module FF( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  output [31:0] io_rPort_0_output_0, // @[:@6.4]
  input  [31:0] io_wPort_0_data_0, // @[:@6.4]
  input         io_wPort_0_reset, // @[:@6.4]
  input         io_wPort_0_en_0 // @[:@6.4]
);
  reg [31:0] ff; // @[MemPrimitives.scala 173:19:@21.4]
  reg [31:0] _RAND_0;
  wire [31:0] _T_68; // @[MemPrimitives.scala 177:32:@23.4]
  wire [31:0] _T_69; // @[MemPrimitives.scala 177:12:@24.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 177:32:@23.4]
  assign _T_69 = io_wPort_0_reset ? 32'h0 : _T_68; // @[MemPrimitives.scala 177:12:@24.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 178:34:@26.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 32'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 32'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SRFF( // @[:@28.2]
  input   clock, // @[:@29.4]
  input   reset, // @[:@30.4]
  input   io_input_set, // @[:@31.4]
  input   io_input_reset, // @[:@31.4]
  input   io_input_asyn_reset, // @[:@31.4]
  output  io_output // @[:@31.4]
);
  reg  _T_15; // @[SRFF.scala 20:21:@33.4]
  reg [31:0] _RAND_0;
  wire  _T_19; // @[SRFF.scala 21:74:@34.4]
  wire  _T_20; // @[SRFF.scala 21:48:@35.4]
  wire  _T_21; // @[SRFF.scala 21:14:@36.4]
  assign _T_19 = io_input_reset ? 1'h0 : _T_15; // @[SRFF.scala 21:74:@34.4]
  assign _T_20 = io_input_set ? 1'h1 : _T_19; // @[SRFF.scala 21:48:@35.4]
  assign _T_21 = io_input_asyn_reset ? 1'h0 : _T_20; // @[SRFF.scala 21:14:@36.4]
  assign io_output = io_input_asyn_reset ? 1'h0 : _T_15; // @[SRFF.scala 22:15:@39.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_15 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_15 <= 1'h0;
    end else begin
      if (io_input_asyn_reset) begin
        _T_15 <= 1'h0;
      end else begin
        if (io_input_set) begin
          _T_15 <= 1'h1;
        end else begin
          if (io_input_reset) begin
            _T_15 <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module SingleCounter( // @[:@41.2]
  input   clock, // @[:@42.4]
  input   reset, // @[:@43.4]
  input   io_input_reset, // @[:@44.4]
  output  io_output_done // @[:@44.4]
);
  wire  bases_0_clock; // @[Counter.scala 253:53:@57.4]
  wire  bases_0_reset; // @[Counter.scala 253:53:@57.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 253:53:@57.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 253:53:@57.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 253:53:@57.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 253:53:@57.4]
  wire  SRFF_clock; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_reset; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_input_set; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_output; // @[Counter.scala 255:22:@73.4]
  wire [31:0] _T_48; // @[Counter.scala 279:52:@101.4]
  wire [32:0] _T_50; // @[Counter.scala 283:33:@102.4]
  wire [31:0] _T_51; // @[Counter.scala 283:33:@103.4]
  wire [31:0] _T_52; // @[Counter.scala 283:33:@104.4]
  wire  _T_57; // @[Counter.scala 285:18:@106.4]
  wire [31:0] _T_68; // @[Counter.scala 291:115:@114.4]
  wire [31:0] _T_71; // @[Counter.scala 291:152:@117.4]
  wire [31:0] _T_72; // @[Counter.scala 291:74:@118.4]
  FF bases_0 ( // @[Counter.scala 253:53:@57.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 255:22:@73.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 279:52:@101.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@102.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@103.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 283:33:@104.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh1); // @[Counter.scala 285:18:@106.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 291:115:@114.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 291:152:@117.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 291:74:@118.4]
  assign io_output_done = $signed(_T_52) >= $signed(32'sh1); // @[Counter.scala 325:20:@127.4]
  assign bases_0_clock = clock; // @[:@58.4]
  assign bases_0_reset = reset; // @[:@59.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 291:31:@120.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 273:27:@99.4]
  assign bases_0_io_wPort_0_en_0 = 1'h1; // @[Counter.scala 276:29:@100.4]
  assign SRFF_clock = clock; // @[:@74.4]
  assign SRFF_reset = reset; // @[:@75.4]
  assign SRFF_io_input_set = io_input_reset == 1'h0; // @[Counter.scala 256:23:@78.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 257:25:@80.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 258:30:@81.4]
endmodule
module RetimeWrapper( // @[:@144.2]
  input   clock, // @[:@145.4]
  input   reset, // @[:@146.4]
  input   io_flow, // @[:@147.4]
  input   io_in, // @[:@147.4]
  output  io_out // @[:@147.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@149.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@149.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@162.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@161.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@160.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@159.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@158.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@156.4]
endmodule
module RootController_sm( // @[:@351.2]
  input   clock, // @[:@352.4]
  input   reset, // @[:@353.4]
  input   io_enable, // @[:@354.4]
  output  io_done, // @[:@354.4]
  input   io_rst, // @[:@354.4]
  input   io_ctrDone, // @[:@354.4]
  output  io_ctrInc, // @[:@354.4]
  input   io_doneIn_0, // @[:@354.4]
  input   io_doneIn_1, // @[:@354.4]
  output  io_enableOut_0, // @[:@354.4]
  output  io_enableOut_1, // @[:@354.4]
  output  io_childAck_0, // @[:@354.4]
  output  io_childAck_1 // @[:@354.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@357.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@357.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@357.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@357.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@357.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@357.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@360.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@360.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@360.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@360.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@360.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@360.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@363.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@363.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@363.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@363.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@363.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@363.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@366.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@366.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@366.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@366.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@366.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@366.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@395.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@395.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@395.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@395.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@395.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@395.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@398.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@398.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@398.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@398.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@398.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@398.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@427.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@427.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@427.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@427.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@427.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@523.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@523.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@523.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@523.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@523.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@540.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@540.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@540.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@540.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@540.4]
  wire  allDone; // @[Controllers.scala 80:47:@369.4]
  wire  _T_77; // @[Controllers.scala 81:26:@370.4]
  wire  finished; // @[Controllers.scala 81:37:@371.4]
  wire  synchronize; // @[package.scala 96:25:@432.4 package.scala 96:25:@433.4]
  wire  _T_144; // @[Controllers.scala 128:33:@441.4]
  wire  _T_146; // @[Controllers.scala 128:54:@442.4]
  wire  _T_147; // @[Controllers.scala 128:52:@443.4]
  wire  _T_148; // @[Controllers.scala 128:66:@444.4]
  wire  _T_150; // @[Controllers.scala 128:98:@446.4]
  wire  _T_151; // @[Controllers.scala 128:96:@447.4]
  wire  _T_153; // @[Controllers.scala 128:123:@448.4]
  wire  _T_155; // @[Controllers.scala 129:48:@451.4]
  wire  _T_160; // @[Controllers.scala 130:52:@456.4]
  wire  _T_161; // @[Controllers.scala 130:50:@457.4]
  wire  _T_169; // @[Controllers.scala 130:129:@463.4]
  wire  _T_172; // @[Controllers.scala 131:45:@466.4]
  wire  _T_175; // @[Controllers.scala 135:80:@470.4]
  wire  _T_176; // @[Controllers.scala 135:78:@471.4]
  wire  _T_178; // @[Controllers.scala 135:105:@472.4]
  wire  _T_179; // @[Controllers.scala 135:103:@473.4]
  wire  _T_180; // @[Controllers.scala 135:119:@474.4]
  wire  _T_182; // @[Controllers.scala 135:51:@476.4]
  wire  _T_205; // @[Controllers.scala 213:68:@501.4]
  wire  _T_207; // @[Controllers.scala 213:90:@503.4]
  wire  _T_209; // @[Controllers.scala 213:132:@505.4]
  wire  _T_210; // @[Controllers.scala 213:130:@506.4]
  wire  _T_211; // @[Controllers.scala 213:156:@507.4]
  wire  _T_213; // @[Controllers.scala 213:68:@510.4]
  wire  _T_215; // @[Controllers.scala 213:90:@512.4]
  wire  _T_222; // @[package.scala 100:49:@518.4]
  reg  _T_225; // @[package.scala 48:56:@519.4]
  reg [31:0] _RAND_0;
  reg  _T_239; // @[package.scala 48:56:@537.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@357.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@360.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@363.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@366.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@395.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@398.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@427.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@523.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@540.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  assign allDone = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@369.4]
  assign _T_77 = allDone | io_done; // @[Controllers.scala 81:26:@370.4]
  assign finished = _T_77 | done_1_io_input_set; // @[Controllers.scala 81:37:@371.4]
  assign synchronize = RetimeWrapper_io_out; // @[package.scala 96:25:@432.4 package.scala 96:25:@433.4]
  assign _T_144 = done_0_io_output == 1'h0; // @[Controllers.scala 128:33:@441.4]
  assign _T_146 = io_ctrDone == 1'h0; // @[Controllers.scala 128:54:@442.4]
  assign _T_147 = _T_144 & _T_146; // @[Controllers.scala 128:52:@443.4]
  assign _T_148 = _T_147 & io_enable; // @[Controllers.scala 128:66:@444.4]
  assign _T_150 = ~ iterDone_0_io_output; // @[Controllers.scala 128:98:@446.4]
  assign _T_151 = _T_148 & _T_150; // @[Controllers.scala 128:96:@447.4]
  assign _T_153 = io_doneIn_0 == 1'h0; // @[Controllers.scala 128:123:@448.4]
  assign _T_155 = io_doneIn_0 | io_rst; // @[Controllers.scala 129:48:@451.4]
  assign _T_160 = synchronize == 1'h0; // @[Controllers.scala 130:52:@456.4]
  assign _T_161 = io_doneIn_0 & _T_160; // @[Controllers.scala 130:50:@457.4]
  assign _T_169 = finished == 1'h0; // @[Controllers.scala 130:129:@463.4]
  assign _T_172 = io_rst == 1'h0; // @[Controllers.scala 131:45:@466.4]
  assign _T_175 = ~ iterDone_1_io_output; // @[Controllers.scala 135:80:@470.4]
  assign _T_176 = iterDone_0_io_output & _T_175; // @[Controllers.scala 135:78:@471.4]
  assign _T_178 = io_doneIn_1 == 1'h0; // @[Controllers.scala 135:105:@472.4]
  assign _T_179 = _T_176 & _T_178; // @[Controllers.scala 135:103:@473.4]
  assign _T_180 = _T_179 & io_enable; // @[Controllers.scala 135:119:@474.4]
  assign _T_182 = io_doneIn_0 | _T_180; // @[Controllers.scala 135:51:@476.4]
  assign _T_205 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@501.4]
  assign _T_207 = _T_205 & _T_150; // @[Controllers.scala 213:90:@503.4]
  assign _T_209 = ~ allDone; // @[Controllers.scala 213:132:@505.4]
  assign _T_210 = _T_207 & _T_209; // @[Controllers.scala 213:130:@506.4]
  assign _T_211 = ~ io_ctrDone; // @[Controllers.scala 213:156:@507.4]
  assign _T_213 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@510.4]
  assign _T_215 = _T_213 & _T_175; // @[Controllers.scala 213:90:@512.4]
  assign _T_222 = allDone == 1'h0; // @[package.scala 100:49:@518.4]
  assign io_done = RetimeWrapper_2_io_out; // @[Controllers.scala 245:13:@547.4]
  assign io_ctrInc = io_doneIn_1; // @[Controllers.scala 122:17:@426.4]
  assign io_enableOut_0 = _T_210 & _T_211; // @[Controllers.scala 213:55:@509.4]
  assign io_enableOut_1 = _T_215 & _T_209; // @[Controllers.scala 213:55:@517.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@498.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@500.4]
  assign active_0_clock = clock; // @[:@358.4]
  assign active_0_reset = reset; // @[:@359.4]
  assign active_0_io_input_set = _T_151 & _T_153; // @[Controllers.scala 128:30:@450.4]
  assign active_0_io_input_reset = _T_155 | allDone; // @[Controllers.scala 129:32:@455.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@372.4]
  assign active_1_clock = clock; // @[:@361.4]
  assign active_1_reset = reset; // @[:@362.4]
  assign active_1_io_input_set = _T_182 & _T_160; // @[Controllers.scala 135:32:@479.4]
  assign active_1_io_input_reset = io_doneIn_1 | io_rst; // @[Controllers.scala 136:34:@483.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@373.4]
  assign done_0_clock = clock; // @[:@364.4]
  assign done_0_reset = reset; // @[:@365.4]
  assign done_0_io_input_set = io_ctrDone & _T_172; // @[Controllers.scala 131:28:@469.4]
  assign done_0_io_input_reset = io_rst | allDone; // @[Controllers.scala 86:33:@384.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@374.4]
  assign done_1_clock = clock; // @[:@367.4]
  assign done_1_reset = reset; // @[:@368.4]
  assign done_1_io_input_set = io_ctrDone & _T_172; // @[Controllers.scala 138:30:@496.4]
  assign done_1_io_input_reset = io_rst | allDone; // @[Controllers.scala 86:33:@393.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@375.4]
  assign iterDone_0_clock = clock; // @[:@396.4]
  assign iterDone_0_reset = reset; // @[:@397.4]
  assign iterDone_0_io_input_set = _T_161 & _T_169; // @[Controllers.scala 130:32:@465.4]
  assign iterDone_0_io_input_reset = synchronize | io_rst; // @[Controllers.scala 92:37:@411.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@401.4]
  assign iterDone_1_clock = clock; // @[:@399.4]
  assign iterDone_1_reset = reset; // @[:@400.4]
  assign iterDone_1_io_input_set = io_doneIn_1 & _T_160; // @[Controllers.scala 137:34:@492.4]
  assign iterDone_1_io_input_reset = synchronize | io_rst; // @[Controllers.scala 92:37:@420.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@402.4]
  assign RetimeWrapper_clock = clock; // @[:@428.4]
  assign RetimeWrapper_reset = reset; // @[:@429.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@431.4]
  assign RetimeWrapper_io_in = io_doneIn_1; // @[package.scala 94:16:@430.4]
  assign RetimeWrapper_1_clock = clock; // @[:@524.4]
  assign RetimeWrapper_1_reset = reset; // @[:@525.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@527.4]
  assign RetimeWrapper_1_io_in = allDone & _T_225; // @[package.scala 94:16:@526.4]
  assign RetimeWrapper_2_clock = clock; // @[:@541.4]
  assign RetimeWrapper_2_reset = reset; // @[:@542.4]
  assign RetimeWrapper_2_io_flow = io_enable; // @[package.scala 95:18:@544.4]
  assign RetimeWrapper_2_io_in = allDone & _T_239; // @[package.scala 94:16:@543.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_225 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_239 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_225 <= 1'h0;
    end else begin
      _T_225 <= _T_222;
    end
    if (reset) begin
      _T_239 <= 1'h0;
    end else begin
      _T_239 <= _T_222;
    end
  end
endmodule
module RetimeWrapper_6( // @[:@641.2]
  input         clock, // @[:@642.4]
  input         reset, // @[:@643.4]
  input         io_flow, // @[:@644.4]
  input  [31:0] io_in, // @[:@644.4]
  output [31:0] io_out // @[:@644.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@646.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@646.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@646.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@646.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@646.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@646.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@646.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@659.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@658.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@657.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@656.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@655.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@653.4]
endmodule
module Mem1D( // @[:@661.2]
  input         clock, // @[:@662.4]
  input         reset, // @[:@663.4]
  input         io_r_ofs_0, // @[:@664.4]
  input         io_r_backpressure, // @[:@664.4]
  input         io_w_ofs_0, // @[:@664.4]
  input  [31:0] io_w_data_0, // @[:@664.4]
  input         io_w_en_0, // @[:@664.4]
  output [31:0] io_output // @[:@664.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@674.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@674.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@674.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@674.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@674.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@683.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@683.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@683.4]
  wire [31:0] RetimeWrapper_1_io_in; // @[package.scala 93:22:@683.4]
  wire [31:0] RetimeWrapper_1_io_out; // @[package.scala 93:22:@683.4]
  reg [31:0] _T_127; // @[MemPrimitives.scala 560:26:@668.4]
  reg [31:0] _RAND_0;
  wire  _T_130; // @[MemPrimitives.scala 561:61:@670.4]
  wire  _T_131; // @[MemPrimitives.scala 561:44:@671.4]
  wire [31:0] _T_132; // @[MemPrimitives.scala 561:19:@672.4]
  wire  _T_135; // @[package.scala 96:25:@679.4 package.scala 96:25:@680.4]
  wire  _T_137; // @[Mux.scala 46:19:@681.4]
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@674.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@683.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign _T_130 = io_w_ofs_0 == 1'h0; // @[MemPrimitives.scala 561:61:@670.4]
  assign _T_131 = io_w_en_0 & _T_130; // @[MemPrimitives.scala 561:44:@671.4]
  assign _T_132 = _T_131 ? io_w_data_0 : _T_127; // @[MemPrimitives.scala 561:19:@672.4]
  assign _T_135 = RetimeWrapper_io_out; // @[package.scala 96:25:@679.4 package.scala 96:25:@680.4]
  assign _T_137 = 1'h0 == _T_135; // @[Mux.scala 46:19:@681.4]
  assign io_output = RetimeWrapper_1_io_out; // @[MemPrimitives.scala 565:17:@690.4]
  assign RetimeWrapper_clock = clock; // @[:@675.4]
  assign RetimeWrapper_reset = reset; // @[:@676.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@678.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@677.4]
  assign RetimeWrapper_1_clock = clock; // @[:@684.4]
  assign RetimeWrapper_1_reset = reset; // @[:@685.4]
  assign RetimeWrapper_1_io_flow = io_r_backpressure; // @[package.scala 95:18:@687.4]
  assign RetimeWrapper_1_io_in = _T_137 ? _T_127 : 32'h0; // @[package.scala 94:16:@686.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_127 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_127 <= 32'h0;
    end else begin
      if (_T_131) begin
        _T_127 <= io_w_data_0;
      end
    end
  end
endmodule
module StickySelects( // @[:@2117.2]
  input   io_ins_0, // @[:@2120.4]
  output  io_outs_0 // @[:@2120.4]
);
  assign io_outs_0 = io_ins_0; // @[StickySelects.scala 12:26:@2122.4]
endmodule
module RetimeWrapper_37( // @[:@2241.2]
  input   clock, // @[:@2242.4]
  input   reset, // @[:@2243.4]
  input   io_in, // @[:@2244.4]
  output  io_out // @[:@2244.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@2246.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@2246.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@2246.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@2246.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@2246.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@2246.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@2246.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@2259.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@2258.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@2257.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@2256.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@2255.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@2253.4]
endmodule
module x273_a_0( // @[:@2741.2]
  input         clock, // @[:@2742.4]
  input         reset, // @[:@2743.4]
  input         io_rPort_15_en_0, // @[:@2744.4]
  output [31:0] io_rPort_15_output_0, // @[:@2744.4]
  input         io_rPort_14_en_0, // @[:@2744.4]
  output [31:0] io_rPort_14_output_0, // @[:@2744.4]
  input         io_rPort_13_en_0, // @[:@2744.4]
  output [31:0] io_rPort_13_output_0, // @[:@2744.4]
  input         io_rPort_12_en_0, // @[:@2744.4]
  output [31:0] io_rPort_12_output_0, // @[:@2744.4]
  input         io_rPort_11_en_0, // @[:@2744.4]
  output [31:0] io_rPort_11_output_0, // @[:@2744.4]
  input         io_rPort_10_en_0, // @[:@2744.4]
  output [31:0] io_rPort_10_output_0, // @[:@2744.4]
  input         io_rPort_9_en_0, // @[:@2744.4]
  output [31:0] io_rPort_9_output_0, // @[:@2744.4]
  input         io_rPort_8_en_0, // @[:@2744.4]
  output [31:0] io_rPort_8_output_0, // @[:@2744.4]
  input         io_rPort_7_en_0, // @[:@2744.4]
  output [31:0] io_rPort_7_output_0, // @[:@2744.4]
  input         io_rPort_6_en_0, // @[:@2744.4]
  output [31:0] io_rPort_6_output_0, // @[:@2744.4]
  input         io_rPort_5_en_0, // @[:@2744.4]
  output [31:0] io_rPort_5_output_0, // @[:@2744.4]
  input         io_rPort_4_en_0, // @[:@2744.4]
  output [31:0] io_rPort_4_output_0, // @[:@2744.4]
  input         io_rPort_3_en_0, // @[:@2744.4]
  output [31:0] io_rPort_3_output_0, // @[:@2744.4]
  input         io_rPort_2_en_0, // @[:@2744.4]
  output [31:0] io_rPort_2_output_0, // @[:@2744.4]
  input         io_rPort_1_en_0, // @[:@2744.4]
  output [31:0] io_rPort_1_output_0, // @[:@2744.4]
  input         io_rPort_0_en_0, // @[:@2744.4]
  output [31:0] io_rPort_0_output_0, // @[:@2744.4]
  input  [4:0]  io_wPort_0_banks_0, // @[:@2744.4]
  input         io_wPort_0_ofs_0, // @[:@2744.4]
  input  [31:0] io_wPort_0_data_0, // @[:@2744.4]
  input         io_wPort_0_en_0 // @[:@2744.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@2834.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@2834.4]
  wire  Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@2834.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@2834.4]
  wire  Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@2834.4]
  wire [31:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@2834.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@2834.4]
  wire [31:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@2834.4]
  wire  Mem1D_1_clock; // @[MemPrimitives.scala 64:21:@2850.4]
  wire  Mem1D_1_reset; // @[MemPrimitives.scala 64:21:@2850.4]
  wire  Mem1D_1_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@2850.4]
  wire  Mem1D_1_io_r_backpressure; // @[MemPrimitives.scala 64:21:@2850.4]
  wire  Mem1D_1_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@2850.4]
  wire [31:0] Mem1D_1_io_w_data_0; // @[MemPrimitives.scala 64:21:@2850.4]
  wire  Mem1D_1_io_w_en_0; // @[MemPrimitives.scala 64:21:@2850.4]
  wire [31:0] Mem1D_1_io_output; // @[MemPrimitives.scala 64:21:@2850.4]
  wire  Mem1D_2_clock; // @[MemPrimitives.scala 64:21:@2866.4]
  wire  Mem1D_2_reset; // @[MemPrimitives.scala 64:21:@2866.4]
  wire  Mem1D_2_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@2866.4]
  wire  Mem1D_2_io_r_backpressure; // @[MemPrimitives.scala 64:21:@2866.4]
  wire  Mem1D_2_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@2866.4]
  wire [31:0] Mem1D_2_io_w_data_0; // @[MemPrimitives.scala 64:21:@2866.4]
  wire  Mem1D_2_io_w_en_0; // @[MemPrimitives.scala 64:21:@2866.4]
  wire [31:0] Mem1D_2_io_output; // @[MemPrimitives.scala 64:21:@2866.4]
  wire  Mem1D_3_clock; // @[MemPrimitives.scala 64:21:@2882.4]
  wire  Mem1D_3_reset; // @[MemPrimitives.scala 64:21:@2882.4]
  wire  Mem1D_3_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@2882.4]
  wire  Mem1D_3_io_r_backpressure; // @[MemPrimitives.scala 64:21:@2882.4]
  wire  Mem1D_3_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@2882.4]
  wire [31:0] Mem1D_3_io_w_data_0; // @[MemPrimitives.scala 64:21:@2882.4]
  wire  Mem1D_3_io_w_en_0; // @[MemPrimitives.scala 64:21:@2882.4]
  wire [31:0] Mem1D_3_io_output; // @[MemPrimitives.scala 64:21:@2882.4]
  wire  Mem1D_4_clock; // @[MemPrimitives.scala 64:21:@2898.4]
  wire  Mem1D_4_reset; // @[MemPrimitives.scala 64:21:@2898.4]
  wire  Mem1D_4_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@2898.4]
  wire  Mem1D_4_io_r_backpressure; // @[MemPrimitives.scala 64:21:@2898.4]
  wire  Mem1D_4_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@2898.4]
  wire [31:0] Mem1D_4_io_w_data_0; // @[MemPrimitives.scala 64:21:@2898.4]
  wire  Mem1D_4_io_w_en_0; // @[MemPrimitives.scala 64:21:@2898.4]
  wire [31:0] Mem1D_4_io_output; // @[MemPrimitives.scala 64:21:@2898.4]
  wire  Mem1D_5_clock; // @[MemPrimitives.scala 64:21:@2914.4]
  wire  Mem1D_5_reset; // @[MemPrimitives.scala 64:21:@2914.4]
  wire  Mem1D_5_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@2914.4]
  wire  Mem1D_5_io_r_backpressure; // @[MemPrimitives.scala 64:21:@2914.4]
  wire  Mem1D_5_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@2914.4]
  wire [31:0] Mem1D_5_io_w_data_0; // @[MemPrimitives.scala 64:21:@2914.4]
  wire  Mem1D_5_io_w_en_0; // @[MemPrimitives.scala 64:21:@2914.4]
  wire [31:0] Mem1D_5_io_output; // @[MemPrimitives.scala 64:21:@2914.4]
  wire  Mem1D_6_clock; // @[MemPrimitives.scala 64:21:@2930.4]
  wire  Mem1D_6_reset; // @[MemPrimitives.scala 64:21:@2930.4]
  wire  Mem1D_6_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@2930.4]
  wire  Mem1D_6_io_r_backpressure; // @[MemPrimitives.scala 64:21:@2930.4]
  wire  Mem1D_6_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@2930.4]
  wire [31:0] Mem1D_6_io_w_data_0; // @[MemPrimitives.scala 64:21:@2930.4]
  wire  Mem1D_6_io_w_en_0; // @[MemPrimitives.scala 64:21:@2930.4]
  wire [31:0] Mem1D_6_io_output; // @[MemPrimitives.scala 64:21:@2930.4]
  wire  Mem1D_7_clock; // @[MemPrimitives.scala 64:21:@2946.4]
  wire  Mem1D_7_reset; // @[MemPrimitives.scala 64:21:@2946.4]
  wire  Mem1D_7_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@2946.4]
  wire  Mem1D_7_io_r_backpressure; // @[MemPrimitives.scala 64:21:@2946.4]
  wire  Mem1D_7_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@2946.4]
  wire [31:0] Mem1D_7_io_w_data_0; // @[MemPrimitives.scala 64:21:@2946.4]
  wire  Mem1D_7_io_w_en_0; // @[MemPrimitives.scala 64:21:@2946.4]
  wire [31:0] Mem1D_7_io_output; // @[MemPrimitives.scala 64:21:@2946.4]
  wire  Mem1D_8_clock; // @[MemPrimitives.scala 64:21:@2962.4]
  wire  Mem1D_8_reset; // @[MemPrimitives.scala 64:21:@2962.4]
  wire  Mem1D_8_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@2962.4]
  wire  Mem1D_8_io_r_backpressure; // @[MemPrimitives.scala 64:21:@2962.4]
  wire  Mem1D_8_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@2962.4]
  wire [31:0] Mem1D_8_io_w_data_0; // @[MemPrimitives.scala 64:21:@2962.4]
  wire  Mem1D_8_io_w_en_0; // @[MemPrimitives.scala 64:21:@2962.4]
  wire [31:0] Mem1D_8_io_output; // @[MemPrimitives.scala 64:21:@2962.4]
  wire  Mem1D_9_clock; // @[MemPrimitives.scala 64:21:@2978.4]
  wire  Mem1D_9_reset; // @[MemPrimitives.scala 64:21:@2978.4]
  wire  Mem1D_9_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@2978.4]
  wire  Mem1D_9_io_r_backpressure; // @[MemPrimitives.scala 64:21:@2978.4]
  wire  Mem1D_9_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@2978.4]
  wire [31:0] Mem1D_9_io_w_data_0; // @[MemPrimitives.scala 64:21:@2978.4]
  wire  Mem1D_9_io_w_en_0; // @[MemPrimitives.scala 64:21:@2978.4]
  wire [31:0] Mem1D_9_io_output; // @[MemPrimitives.scala 64:21:@2978.4]
  wire  Mem1D_10_clock; // @[MemPrimitives.scala 64:21:@2994.4]
  wire  Mem1D_10_reset; // @[MemPrimitives.scala 64:21:@2994.4]
  wire  Mem1D_10_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@2994.4]
  wire  Mem1D_10_io_r_backpressure; // @[MemPrimitives.scala 64:21:@2994.4]
  wire  Mem1D_10_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@2994.4]
  wire [31:0] Mem1D_10_io_w_data_0; // @[MemPrimitives.scala 64:21:@2994.4]
  wire  Mem1D_10_io_w_en_0; // @[MemPrimitives.scala 64:21:@2994.4]
  wire [31:0] Mem1D_10_io_output; // @[MemPrimitives.scala 64:21:@2994.4]
  wire  Mem1D_11_clock; // @[MemPrimitives.scala 64:21:@3010.4]
  wire  Mem1D_11_reset; // @[MemPrimitives.scala 64:21:@3010.4]
  wire  Mem1D_11_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@3010.4]
  wire  Mem1D_11_io_r_backpressure; // @[MemPrimitives.scala 64:21:@3010.4]
  wire  Mem1D_11_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@3010.4]
  wire [31:0] Mem1D_11_io_w_data_0; // @[MemPrimitives.scala 64:21:@3010.4]
  wire  Mem1D_11_io_w_en_0; // @[MemPrimitives.scala 64:21:@3010.4]
  wire [31:0] Mem1D_11_io_output; // @[MemPrimitives.scala 64:21:@3010.4]
  wire  Mem1D_12_clock; // @[MemPrimitives.scala 64:21:@3026.4]
  wire  Mem1D_12_reset; // @[MemPrimitives.scala 64:21:@3026.4]
  wire  Mem1D_12_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@3026.4]
  wire  Mem1D_12_io_r_backpressure; // @[MemPrimitives.scala 64:21:@3026.4]
  wire  Mem1D_12_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@3026.4]
  wire [31:0] Mem1D_12_io_w_data_0; // @[MemPrimitives.scala 64:21:@3026.4]
  wire  Mem1D_12_io_w_en_0; // @[MemPrimitives.scala 64:21:@3026.4]
  wire [31:0] Mem1D_12_io_output; // @[MemPrimitives.scala 64:21:@3026.4]
  wire  Mem1D_13_clock; // @[MemPrimitives.scala 64:21:@3042.4]
  wire  Mem1D_13_reset; // @[MemPrimitives.scala 64:21:@3042.4]
  wire  Mem1D_13_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@3042.4]
  wire  Mem1D_13_io_r_backpressure; // @[MemPrimitives.scala 64:21:@3042.4]
  wire  Mem1D_13_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@3042.4]
  wire [31:0] Mem1D_13_io_w_data_0; // @[MemPrimitives.scala 64:21:@3042.4]
  wire  Mem1D_13_io_w_en_0; // @[MemPrimitives.scala 64:21:@3042.4]
  wire [31:0] Mem1D_13_io_output; // @[MemPrimitives.scala 64:21:@3042.4]
  wire  Mem1D_14_clock; // @[MemPrimitives.scala 64:21:@3058.4]
  wire  Mem1D_14_reset; // @[MemPrimitives.scala 64:21:@3058.4]
  wire  Mem1D_14_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@3058.4]
  wire  Mem1D_14_io_r_backpressure; // @[MemPrimitives.scala 64:21:@3058.4]
  wire  Mem1D_14_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@3058.4]
  wire [31:0] Mem1D_14_io_w_data_0; // @[MemPrimitives.scala 64:21:@3058.4]
  wire  Mem1D_14_io_w_en_0; // @[MemPrimitives.scala 64:21:@3058.4]
  wire [31:0] Mem1D_14_io_output; // @[MemPrimitives.scala 64:21:@3058.4]
  wire  Mem1D_15_clock; // @[MemPrimitives.scala 64:21:@3074.4]
  wire  Mem1D_15_reset; // @[MemPrimitives.scala 64:21:@3074.4]
  wire  Mem1D_15_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@3074.4]
  wire  Mem1D_15_io_r_backpressure; // @[MemPrimitives.scala 64:21:@3074.4]
  wire  Mem1D_15_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@3074.4]
  wire [31:0] Mem1D_15_io_w_data_0; // @[MemPrimitives.scala 64:21:@3074.4]
  wire  Mem1D_15_io_w_en_0; // @[MemPrimitives.scala 64:21:@3074.4]
  wire [31:0] Mem1D_15_io_output; // @[MemPrimitives.scala 64:21:@3074.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 121:29:@3251.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 121:29:@3251.4]
  wire  StickySelects_1_io_ins_0; // @[MemPrimitives.scala 121:29:@3265.4]
  wire  StickySelects_1_io_outs_0; // @[MemPrimitives.scala 121:29:@3265.4]
  wire  StickySelects_2_io_ins_0; // @[MemPrimitives.scala 121:29:@3279.4]
  wire  StickySelects_2_io_outs_0; // @[MemPrimitives.scala 121:29:@3279.4]
  wire  StickySelects_3_io_ins_0; // @[MemPrimitives.scala 121:29:@3293.4]
  wire  StickySelects_3_io_outs_0; // @[MemPrimitives.scala 121:29:@3293.4]
  wire  StickySelects_4_io_ins_0; // @[MemPrimitives.scala 121:29:@3307.4]
  wire  StickySelects_4_io_outs_0; // @[MemPrimitives.scala 121:29:@3307.4]
  wire  StickySelects_5_io_ins_0; // @[MemPrimitives.scala 121:29:@3321.4]
  wire  StickySelects_5_io_outs_0; // @[MemPrimitives.scala 121:29:@3321.4]
  wire  StickySelects_6_io_ins_0; // @[MemPrimitives.scala 121:29:@3335.4]
  wire  StickySelects_6_io_outs_0; // @[MemPrimitives.scala 121:29:@3335.4]
  wire  StickySelects_7_io_ins_0; // @[MemPrimitives.scala 121:29:@3349.4]
  wire  StickySelects_7_io_outs_0; // @[MemPrimitives.scala 121:29:@3349.4]
  wire  StickySelects_8_io_ins_0; // @[MemPrimitives.scala 121:29:@3363.4]
  wire  StickySelects_8_io_outs_0; // @[MemPrimitives.scala 121:29:@3363.4]
  wire  StickySelects_9_io_ins_0; // @[MemPrimitives.scala 121:29:@3377.4]
  wire  StickySelects_9_io_outs_0; // @[MemPrimitives.scala 121:29:@3377.4]
  wire  StickySelects_10_io_ins_0; // @[MemPrimitives.scala 121:29:@3391.4]
  wire  StickySelects_10_io_outs_0; // @[MemPrimitives.scala 121:29:@3391.4]
  wire  StickySelects_11_io_ins_0; // @[MemPrimitives.scala 121:29:@3405.4]
  wire  StickySelects_11_io_outs_0; // @[MemPrimitives.scala 121:29:@3405.4]
  wire  StickySelects_12_io_ins_0; // @[MemPrimitives.scala 121:29:@3419.4]
  wire  StickySelects_12_io_outs_0; // @[MemPrimitives.scala 121:29:@3419.4]
  wire  StickySelects_13_io_ins_0; // @[MemPrimitives.scala 121:29:@3433.4]
  wire  StickySelects_13_io_outs_0; // @[MemPrimitives.scala 121:29:@3433.4]
  wire  StickySelects_14_io_ins_0; // @[MemPrimitives.scala 121:29:@3447.4]
  wire  StickySelects_14_io_outs_0; // @[MemPrimitives.scala 121:29:@3447.4]
  wire  StickySelects_15_io_ins_0; // @[MemPrimitives.scala 121:29:@3461.4]
  wire  StickySelects_15_io_outs_0; // @[MemPrimitives.scala 121:29:@3461.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3475.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3475.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@3475.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@3475.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@3484.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@3484.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@3484.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@3484.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@3493.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@3493.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@3493.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@3493.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@3502.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@3502.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@3502.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@3502.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@3511.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@3511.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@3511.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@3511.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@3520.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@3520.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@3520.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@3520.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@3529.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@3529.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@3529.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@3529.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@3538.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@3538.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@3538.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@3538.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@3547.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@3547.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@3547.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@3547.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@3556.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@3556.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@3556.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@3556.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@3565.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@3565.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@3565.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@3565.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@3574.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@3574.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@3574.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@3574.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@3583.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@3583.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@3583.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@3583.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@3592.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@3592.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@3592.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@3592.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@3601.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@3601.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@3601.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@3601.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@3610.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@3610.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@3610.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@3610.4]
  wire  _T_458; // @[MemPrimitives.scala 82:210:@3090.4]
  wire  _T_459; // @[MemPrimitives.scala 83:102:@3091.4]
  wire [33:0] _T_461; // @[Cat.scala 30:58:@3093.4]
  wire  _T_466; // @[MemPrimitives.scala 82:210:@3100.4]
  wire  _T_467; // @[MemPrimitives.scala 83:102:@3101.4]
  wire [33:0] _T_469; // @[Cat.scala 30:58:@3103.4]
  wire  _T_474; // @[MemPrimitives.scala 82:210:@3110.4]
  wire  _T_475; // @[MemPrimitives.scala 83:102:@3111.4]
  wire [33:0] _T_477; // @[Cat.scala 30:58:@3113.4]
  wire  _T_482; // @[MemPrimitives.scala 82:210:@3120.4]
  wire  _T_483; // @[MemPrimitives.scala 83:102:@3121.4]
  wire [33:0] _T_485; // @[Cat.scala 30:58:@3123.4]
  wire  _T_490; // @[MemPrimitives.scala 82:210:@3130.4]
  wire  _T_491; // @[MemPrimitives.scala 83:102:@3131.4]
  wire [33:0] _T_493; // @[Cat.scala 30:58:@3133.4]
  wire  _T_498; // @[MemPrimitives.scala 82:210:@3140.4]
  wire  _T_499; // @[MemPrimitives.scala 83:102:@3141.4]
  wire [33:0] _T_501; // @[Cat.scala 30:58:@3143.4]
  wire  _T_506; // @[MemPrimitives.scala 82:210:@3150.4]
  wire  _T_507; // @[MemPrimitives.scala 83:102:@3151.4]
  wire [33:0] _T_509; // @[Cat.scala 30:58:@3153.4]
  wire  _T_514; // @[MemPrimitives.scala 82:210:@3160.4]
  wire  _T_515; // @[MemPrimitives.scala 83:102:@3161.4]
  wire [33:0] _T_517; // @[Cat.scala 30:58:@3163.4]
  wire  _T_522; // @[MemPrimitives.scala 82:210:@3170.4]
  wire  _T_523; // @[MemPrimitives.scala 83:102:@3171.4]
  wire [33:0] _T_525; // @[Cat.scala 30:58:@3173.4]
  wire  _T_530; // @[MemPrimitives.scala 82:210:@3180.4]
  wire  _T_531; // @[MemPrimitives.scala 83:102:@3181.4]
  wire [33:0] _T_533; // @[Cat.scala 30:58:@3183.4]
  wire  _T_538; // @[MemPrimitives.scala 82:210:@3190.4]
  wire  _T_539; // @[MemPrimitives.scala 83:102:@3191.4]
  wire [33:0] _T_541; // @[Cat.scala 30:58:@3193.4]
  wire  _T_546; // @[MemPrimitives.scala 82:210:@3200.4]
  wire  _T_547; // @[MemPrimitives.scala 83:102:@3201.4]
  wire [33:0] _T_549; // @[Cat.scala 30:58:@3203.4]
  wire  _T_554; // @[MemPrimitives.scala 82:210:@3210.4]
  wire  _T_555; // @[MemPrimitives.scala 83:102:@3211.4]
  wire [33:0] _T_557; // @[Cat.scala 30:58:@3213.4]
  wire  _T_562; // @[MemPrimitives.scala 82:210:@3220.4]
  wire  _T_563; // @[MemPrimitives.scala 83:102:@3221.4]
  wire [33:0] _T_565; // @[Cat.scala 30:58:@3223.4]
  wire  _T_570; // @[MemPrimitives.scala 82:210:@3230.4]
  wire  _T_571; // @[MemPrimitives.scala 83:102:@3231.4]
  wire [33:0] _T_573; // @[Cat.scala 30:58:@3233.4]
  wire  _T_578; // @[MemPrimitives.scala 82:210:@3240.4]
  wire  _T_579; // @[MemPrimitives.scala 83:102:@3241.4]
  wire [33:0] _T_581; // @[Cat.scala 30:58:@3243.4]
  wire  _T_587; // @[MemPrimitives.scala 123:41:@3255.4]
  wire [2:0] _T_589; // @[Cat.scala 30:58:@3257.4]
  wire  _T_595; // @[MemPrimitives.scala 123:41:@3269.4]
  wire [2:0] _T_597; // @[Cat.scala 30:58:@3271.4]
  wire  _T_603; // @[MemPrimitives.scala 123:41:@3283.4]
  wire [2:0] _T_605; // @[Cat.scala 30:58:@3285.4]
  wire  _T_611; // @[MemPrimitives.scala 123:41:@3297.4]
  wire [2:0] _T_613; // @[Cat.scala 30:58:@3299.4]
  wire  _T_619; // @[MemPrimitives.scala 123:41:@3311.4]
  wire [2:0] _T_621; // @[Cat.scala 30:58:@3313.4]
  wire  _T_627; // @[MemPrimitives.scala 123:41:@3325.4]
  wire [2:0] _T_629; // @[Cat.scala 30:58:@3327.4]
  wire  _T_635; // @[MemPrimitives.scala 123:41:@3339.4]
  wire [2:0] _T_637; // @[Cat.scala 30:58:@3341.4]
  wire  _T_643; // @[MemPrimitives.scala 123:41:@3353.4]
  wire [2:0] _T_645; // @[Cat.scala 30:58:@3355.4]
  wire  _T_651; // @[MemPrimitives.scala 123:41:@3367.4]
  wire [2:0] _T_653; // @[Cat.scala 30:58:@3369.4]
  wire  _T_659; // @[MemPrimitives.scala 123:41:@3381.4]
  wire [2:0] _T_661; // @[Cat.scala 30:58:@3383.4]
  wire  _T_667; // @[MemPrimitives.scala 123:41:@3395.4]
  wire [2:0] _T_669; // @[Cat.scala 30:58:@3397.4]
  wire  _T_675; // @[MemPrimitives.scala 123:41:@3409.4]
  wire [2:0] _T_677; // @[Cat.scala 30:58:@3411.4]
  wire  _T_683; // @[MemPrimitives.scala 123:41:@3423.4]
  wire [2:0] _T_685; // @[Cat.scala 30:58:@3425.4]
  wire  _T_691; // @[MemPrimitives.scala 123:41:@3437.4]
  wire [2:0] _T_693; // @[Cat.scala 30:58:@3439.4]
  wire  _T_699; // @[MemPrimitives.scala 123:41:@3451.4]
  wire [2:0] _T_701; // @[Cat.scala 30:58:@3453.4]
  wire  _T_707; // @[MemPrimitives.scala 123:41:@3465.4]
  wire [2:0] _T_709; // @[Cat.scala 30:58:@3467.4]
  Mem1D Mem1D ( // @[MemPrimitives.scala 64:21:@2834.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  Mem1D Mem1D_1 ( // @[MemPrimitives.scala 64:21:@2850.4]
    .clock(Mem1D_1_clock),
    .reset(Mem1D_1_reset),
    .io_r_ofs_0(Mem1D_1_io_r_ofs_0),
    .io_r_backpressure(Mem1D_1_io_r_backpressure),
    .io_w_ofs_0(Mem1D_1_io_w_ofs_0),
    .io_w_data_0(Mem1D_1_io_w_data_0),
    .io_w_en_0(Mem1D_1_io_w_en_0),
    .io_output(Mem1D_1_io_output)
  );
  Mem1D Mem1D_2 ( // @[MemPrimitives.scala 64:21:@2866.4]
    .clock(Mem1D_2_clock),
    .reset(Mem1D_2_reset),
    .io_r_ofs_0(Mem1D_2_io_r_ofs_0),
    .io_r_backpressure(Mem1D_2_io_r_backpressure),
    .io_w_ofs_0(Mem1D_2_io_w_ofs_0),
    .io_w_data_0(Mem1D_2_io_w_data_0),
    .io_w_en_0(Mem1D_2_io_w_en_0),
    .io_output(Mem1D_2_io_output)
  );
  Mem1D Mem1D_3 ( // @[MemPrimitives.scala 64:21:@2882.4]
    .clock(Mem1D_3_clock),
    .reset(Mem1D_3_reset),
    .io_r_ofs_0(Mem1D_3_io_r_ofs_0),
    .io_r_backpressure(Mem1D_3_io_r_backpressure),
    .io_w_ofs_0(Mem1D_3_io_w_ofs_0),
    .io_w_data_0(Mem1D_3_io_w_data_0),
    .io_w_en_0(Mem1D_3_io_w_en_0),
    .io_output(Mem1D_3_io_output)
  );
  Mem1D Mem1D_4 ( // @[MemPrimitives.scala 64:21:@2898.4]
    .clock(Mem1D_4_clock),
    .reset(Mem1D_4_reset),
    .io_r_ofs_0(Mem1D_4_io_r_ofs_0),
    .io_r_backpressure(Mem1D_4_io_r_backpressure),
    .io_w_ofs_0(Mem1D_4_io_w_ofs_0),
    .io_w_data_0(Mem1D_4_io_w_data_0),
    .io_w_en_0(Mem1D_4_io_w_en_0),
    .io_output(Mem1D_4_io_output)
  );
  Mem1D Mem1D_5 ( // @[MemPrimitives.scala 64:21:@2914.4]
    .clock(Mem1D_5_clock),
    .reset(Mem1D_5_reset),
    .io_r_ofs_0(Mem1D_5_io_r_ofs_0),
    .io_r_backpressure(Mem1D_5_io_r_backpressure),
    .io_w_ofs_0(Mem1D_5_io_w_ofs_0),
    .io_w_data_0(Mem1D_5_io_w_data_0),
    .io_w_en_0(Mem1D_5_io_w_en_0),
    .io_output(Mem1D_5_io_output)
  );
  Mem1D Mem1D_6 ( // @[MemPrimitives.scala 64:21:@2930.4]
    .clock(Mem1D_6_clock),
    .reset(Mem1D_6_reset),
    .io_r_ofs_0(Mem1D_6_io_r_ofs_0),
    .io_r_backpressure(Mem1D_6_io_r_backpressure),
    .io_w_ofs_0(Mem1D_6_io_w_ofs_0),
    .io_w_data_0(Mem1D_6_io_w_data_0),
    .io_w_en_0(Mem1D_6_io_w_en_0),
    .io_output(Mem1D_6_io_output)
  );
  Mem1D Mem1D_7 ( // @[MemPrimitives.scala 64:21:@2946.4]
    .clock(Mem1D_7_clock),
    .reset(Mem1D_7_reset),
    .io_r_ofs_0(Mem1D_7_io_r_ofs_0),
    .io_r_backpressure(Mem1D_7_io_r_backpressure),
    .io_w_ofs_0(Mem1D_7_io_w_ofs_0),
    .io_w_data_0(Mem1D_7_io_w_data_0),
    .io_w_en_0(Mem1D_7_io_w_en_0),
    .io_output(Mem1D_7_io_output)
  );
  Mem1D Mem1D_8 ( // @[MemPrimitives.scala 64:21:@2962.4]
    .clock(Mem1D_8_clock),
    .reset(Mem1D_8_reset),
    .io_r_ofs_0(Mem1D_8_io_r_ofs_0),
    .io_r_backpressure(Mem1D_8_io_r_backpressure),
    .io_w_ofs_0(Mem1D_8_io_w_ofs_0),
    .io_w_data_0(Mem1D_8_io_w_data_0),
    .io_w_en_0(Mem1D_8_io_w_en_0),
    .io_output(Mem1D_8_io_output)
  );
  Mem1D Mem1D_9 ( // @[MemPrimitives.scala 64:21:@2978.4]
    .clock(Mem1D_9_clock),
    .reset(Mem1D_9_reset),
    .io_r_ofs_0(Mem1D_9_io_r_ofs_0),
    .io_r_backpressure(Mem1D_9_io_r_backpressure),
    .io_w_ofs_0(Mem1D_9_io_w_ofs_0),
    .io_w_data_0(Mem1D_9_io_w_data_0),
    .io_w_en_0(Mem1D_9_io_w_en_0),
    .io_output(Mem1D_9_io_output)
  );
  Mem1D Mem1D_10 ( // @[MemPrimitives.scala 64:21:@2994.4]
    .clock(Mem1D_10_clock),
    .reset(Mem1D_10_reset),
    .io_r_ofs_0(Mem1D_10_io_r_ofs_0),
    .io_r_backpressure(Mem1D_10_io_r_backpressure),
    .io_w_ofs_0(Mem1D_10_io_w_ofs_0),
    .io_w_data_0(Mem1D_10_io_w_data_0),
    .io_w_en_0(Mem1D_10_io_w_en_0),
    .io_output(Mem1D_10_io_output)
  );
  Mem1D Mem1D_11 ( // @[MemPrimitives.scala 64:21:@3010.4]
    .clock(Mem1D_11_clock),
    .reset(Mem1D_11_reset),
    .io_r_ofs_0(Mem1D_11_io_r_ofs_0),
    .io_r_backpressure(Mem1D_11_io_r_backpressure),
    .io_w_ofs_0(Mem1D_11_io_w_ofs_0),
    .io_w_data_0(Mem1D_11_io_w_data_0),
    .io_w_en_0(Mem1D_11_io_w_en_0),
    .io_output(Mem1D_11_io_output)
  );
  Mem1D Mem1D_12 ( // @[MemPrimitives.scala 64:21:@3026.4]
    .clock(Mem1D_12_clock),
    .reset(Mem1D_12_reset),
    .io_r_ofs_0(Mem1D_12_io_r_ofs_0),
    .io_r_backpressure(Mem1D_12_io_r_backpressure),
    .io_w_ofs_0(Mem1D_12_io_w_ofs_0),
    .io_w_data_0(Mem1D_12_io_w_data_0),
    .io_w_en_0(Mem1D_12_io_w_en_0),
    .io_output(Mem1D_12_io_output)
  );
  Mem1D Mem1D_13 ( // @[MemPrimitives.scala 64:21:@3042.4]
    .clock(Mem1D_13_clock),
    .reset(Mem1D_13_reset),
    .io_r_ofs_0(Mem1D_13_io_r_ofs_0),
    .io_r_backpressure(Mem1D_13_io_r_backpressure),
    .io_w_ofs_0(Mem1D_13_io_w_ofs_0),
    .io_w_data_0(Mem1D_13_io_w_data_0),
    .io_w_en_0(Mem1D_13_io_w_en_0),
    .io_output(Mem1D_13_io_output)
  );
  Mem1D Mem1D_14 ( // @[MemPrimitives.scala 64:21:@3058.4]
    .clock(Mem1D_14_clock),
    .reset(Mem1D_14_reset),
    .io_r_ofs_0(Mem1D_14_io_r_ofs_0),
    .io_r_backpressure(Mem1D_14_io_r_backpressure),
    .io_w_ofs_0(Mem1D_14_io_w_ofs_0),
    .io_w_data_0(Mem1D_14_io_w_data_0),
    .io_w_en_0(Mem1D_14_io_w_en_0),
    .io_output(Mem1D_14_io_output)
  );
  Mem1D Mem1D_15 ( // @[MemPrimitives.scala 64:21:@3074.4]
    .clock(Mem1D_15_clock),
    .reset(Mem1D_15_reset),
    .io_r_ofs_0(Mem1D_15_io_r_ofs_0),
    .io_r_backpressure(Mem1D_15_io_r_backpressure),
    .io_w_ofs_0(Mem1D_15_io_w_ofs_0),
    .io_w_data_0(Mem1D_15_io_w_data_0),
    .io_w_en_0(Mem1D_15_io_w_en_0),
    .io_output(Mem1D_15_io_output)
  );
  StickySelects StickySelects ( // @[MemPrimitives.scala 121:29:@3251.4]
    .io_ins_0(StickySelects_io_ins_0),
    .io_outs_0(StickySelects_io_outs_0)
  );
  StickySelects StickySelects_1 ( // @[MemPrimitives.scala 121:29:@3265.4]
    .io_ins_0(StickySelects_1_io_ins_0),
    .io_outs_0(StickySelects_1_io_outs_0)
  );
  StickySelects StickySelects_2 ( // @[MemPrimitives.scala 121:29:@3279.4]
    .io_ins_0(StickySelects_2_io_ins_0),
    .io_outs_0(StickySelects_2_io_outs_0)
  );
  StickySelects StickySelects_3 ( // @[MemPrimitives.scala 121:29:@3293.4]
    .io_ins_0(StickySelects_3_io_ins_0),
    .io_outs_0(StickySelects_3_io_outs_0)
  );
  StickySelects StickySelects_4 ( // @[MemPrimitives.scala 121:29:@3307.4]
    .io_ins_0(StickySelects_4_io_ins_0),
    .io_outs_0(StickySelects_4_io_outs_0)
  );
  StickySelects StickySelects_5 ( // @[MemPrimitives.scala 121:29:@3321.4]
    .io_ins_0(StickySelects_5_io_ins_0),
    .io_outs_0(StickySelects_5_io_outs_0)
  );
  StickySelects StickySelects_6 ( // @[MemPrimitives.scala 121:29:@3335.4]
    .io_ins_0(StickySelects_6_io_ins_0),
    .io_outs_0(StickySelects_6_io_outs_0)
  );
  StickySelects StickySelects_7 ( // @[MemPrimitives.scala 121:29:@3349.4]
    .io_ins_0(StickySelects_7_io_ins_0),
    .io_outs_0(StickySelects_7_io_outs_0)
  );
  StickySelects StickySelects_8 ( // @[MemPrimitives.scala 121:29:@3363.4]
    .io_ins_0(StickySelects_8_io_ins_0),
    .io_outs_0(StickySelects_8_io_outs_0)
  );
  StickySelects StickySelects_9 ( // @[MemPrimitives.scala 121:29:@3377.4]
    .io_ins_0(StickySelects_9_io_ins_0),
    .io_outs_0(StickySelects_9_io_outs_0)
  );
  StickySelects StickySelects_10 ( // @[MemPrimitives.scala 121:29:@3391.4]
    .io_ins_0(StickySelects_10_io_ins_0),
    .io_outs_0(StickySelects_10_io_outs_0)
  );
  StickySelects StickySelects_11 ( // @[MemPrimitives.scala 121:29:@3405.4]
    .io_ins_0(StickySelects_11_io_ins_0),
    .io_outs_0(StickySelects_11_io_outs_0)
  );
  StickySelects StickySelects_12 ( // @[MemPrimitives.scala 121:29:@3419.4]
    .io_ins_0(StickySelects_12_io_ins_0),
    .io_outs_0(StickySelects_12_io_outs_0)
  );
  StickySelects StickySelects_13 ( // @[MemPrimitives.scala 121:29:@3433.4]
    .io_ins_0(StickySelects_13_io_ins_0),
    .io_outs_0(StickySelects_13_io_outs_0)
  );
  StickySelects StickySelects_14 ( // @[MemPrimitives.scala 121:29:@3447.4]
    .io_ins_0(StickySelects_14_io_ins_0),
    .io_outs_0(StickySelects_14_io_outs_0)
  );
  StickySelects StickySelects_15 ( // @[MemPrimitives.scala 121:29:@3461.4]
    .io_ins_0(StickySelects_15_io_ins_0),
    .io_outs_0(StickySelects_15_io_outs_0)
  );
  RetimeWrapper_37 RetimeWrapper ( // @[package.scala 93:22:@3475.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_37 RetimeWrapper_1 ( // @[package.scala 93:22:@3484.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_37 RetimeWrapper_2 ( // @[package.scala 93:22:@3493.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_37 RetimeWrapper_3 ( // @[package.scala 93:22:@3502.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_37 RetimeWrapper_4 ( // @[package.scala 93:22:@3511.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_37 RetimeWrapper_5 ( // @[package.scala 93:22:@3520.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_37 RetimeWrapper_6 ( // @[package.scala 93:22:@3529.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_37 RetimeWrapper_7 ( // @[package.scala 93:22:@3538.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_37 RetimeWrapper_8 ( // @[package.scala 93:22:@3547.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_37 RetimeWrapper_9 ( // @[package.scala 93:22:@3556.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_37 RetimeWrapper_10 ( // @[package.scala 93:22:@3565.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_37 RetimeWrapper_11 ( // @[package.scala 93:22:@3574.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_37 RetimeWrapper_12 ( // @[package.scala 93:22:@3583.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_37 RetimeWrapper_13 ( // @[package.scala 93:22:@3592.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_37 RetimeWrapper_14 ( // @[package.scala 93:22:@3601.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_37 RetimeWrapper_15 ( // @[package.scala 93:22:@3610.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  assign _T_458 = io_wPort_0_banks_0 == 5'h0; // @[MemPrimitives.scala 82:210:@3090.4]
  assign _T_459 = io_wPort_0_en_0 & _T_458; // @[MemPrimitives.scala 83:102:@3091.4]
  assign _T_461 = {_T_459,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@3093.4]
  assign _T_466 = io_wPort_0_banks_0 == 5'h1; // @[MemPrimitives.scala 82:210:@3100.4]
  assign _T_467 = io_wPort_0_en_0 & _T_466; // @[MemPrimitives.scala 83:102:@3101.4]
  assign _T_469 = {_T_467,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@3103.4]
  assign _T_474 = io_wPort_0_banks_0 == 5'h2; // @[MemPrimitives.scala 82:210:@3110.4]
  assign _T_475 = io_wPort_0_en_0 & _T_474; // @[MemPrimitives.scala 83:102:@3111.4]
  assign _T_477 = {_T_475,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@3113.4]
  assign _T_482 = io_wPort_0_banks_0 == 5'h3; // @[MemPrimitives.scala 82:210:@3120.4]
  assign _T_483 = io_wPort_0_en_0 & _T_482; // @[MemPrimitives.scala 83:102:@3121.4]
  assign _T_485 = {_T_483,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@3123.4]
  assign _T_490 = io_wPort_0_banks_0 == 5'h4; // @[MemPrimitives.scala 82:210:@3130.4]
  assign _T_491 = io_wPort_0_en_0 & _T_490; // @[MemPrimitives.scala 83:102:@3131.4]
  assign _T_493 = {_T_491,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@3133.4]
  assign _T_498 = io_wPort_0_banks_0 == 5'h5; // @[MemPrimitives.scala 82:210:@3140.4]
  assign _T_499 = io_wPort_0_en_0 & _T_498; // @[MemPrimitives.scala 83:102:@3141.4]
  assign _T_501 = {_T_499,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@3143.4]
  assign _T_506 = io_wPort_0_banks_0 == 5'h6; // @[MemPrimitives.scala 82:210:@3150.4]
  assign _T_507 = io_wPort_0_en_0 & _T_506; // @[MemPrimitives.scala 83:102:@3151.4]
  assign _T_509 = {_T_507,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@3153.4]
  assign _T_514 = io_wPort_0_banks_0 == 5'h7; // @[MemPrimitives.scala 82:210:@3160.4]
  assign _T_515 = io_wPort_0_en_0 & _T_514; // @[MemPrimitives.scala 83:102:@3161.4]
  assign _T_517 = {_T_515,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@3163.4]
  assign _T_522 = io_wPort_0_banks_0 == 5'h8; // @[MemPrimitives.scala 82:210:@3170.4]
  assign _T_523 = io_wPort_0_en_0 & _T_522; // @[MemPrimitives.scala 83:102:@3171.4]
  assign _T_525 = {_T_523,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@3173.4]
  assign _T_530 = io_wPort_0_banks_0 == 5'h9; // @[MemPrimitives.scala 82:210:@3180.4]
  assign _T_531 = io_wPort_0_en_0 & _T_530; // @[MemPrimitives.scala 83:102:@3181.4]
  assign _T_533 = {_T_531,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@3183.4]
  assign _T_538 = io_wPort_0_banks_0 == 5'ha; // @[MemPrimitives.scala 82:210:@3190.4]
  assign _T_539 = io_wPort_0_en_0 & _T_538; // @[MemPrimitives.scala 83:102:@3191.4]
  assign _T_541 = {_T_539,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@3193.4]
  assign _T_546 = io_wPort_0_banks_0 == 5'hb; // @[MemPrimitives.scala 82:210:@3200.4]
  assign _T_547 = io_wPort_0_en_0 & _T_546; // @[MemPrimitives.scala 83:102:@3201.4]
  assign _T_549 = {_T_547,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@3203.4]
  assign _T_554 = io_wPort_0_banks_0 == 5'hc; // @[MemPrimitives.scala 82:210:@3210.4]
  assign _T_555 = io_wPort_0_en_0 & _T_554; // @[MemPrimitives.scala 83:102:@3211.4]
  assign _T_557 = {_T_555,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@3213.4]
  assign _T_562 = io_wPort_0_banks_0 == 5'hd; // @[MemPrimitives.scala 82:210:@3220.4]
  assign _T_563 = io_wPort_0_en_0 & _T_562; // @[MemPrimitives.scala 83:102:@3221.4]
  assign _T_565 = {_T_563,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@3223.4]
  assign _T_570 = io_wPort_0_banks_0 == 5'he; // @[MemPrimitives.scala 82:210:@3230.4]
  assign _T_571 = io_wPort_0_en_0 & _T_570; // @[MemPrimitives.scala 83:102:@3231.4]
  assign _T_573 = {_T_571,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@3233.4]
  assign _T_578 = io_wPort_0_banks_0 == 5'hf; // @[MemPrimitives.scala 82:210:@3240.4]
  assign _T_579 = io_wPort_0_en_0 & _T_578; // @[MemPrimitives.scala 83:102:@3241.4]
  assign _T_581 = {_T_579,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@3243.4]
  assign _T_587 = StickySelects_io_outs_0; // @[MemPrimitives.scala 123:41:@3255.4]
  assign _T_589 = {_T_587,1'h1,1'h0}; // @[Cat.scala 30:58:@3257.4]
  assign _T_595 = StickySelects_1_io_outs_0; // @[MemPrimitives.scala 123:41:@3269.4]
  assign _T_597 = {_T_595,1'h1,1'h0}; // @[Cat.scala 30:58:@3271.4]
  assign _T_603 = StickySelects_2_io_outs_0; // @[MemPrimitives.scala 123:41:@3283.4]
  assign _T_605 = {_T_603,1'h1,1'h0}; // @[Cat.scala 30:58:@3285.4]
  assign _T_611 = StickySelects_3_io_outs_0; // @[MemPrimitives.scala 123:41:@3297.4]
  assign _T_613 = {_T_611,1'h1,1'h0}; // @[Cat.scala 30:58:@3299.4]
  assign _T_619 = StickySelects_4_io_outs_0; // @[MemPrimitives.scala 123:41:@3311.4]
  assign _T_621 = {_T_619,1'h1,1'h0}; // @[Cat.scala 30:58:@3313.4]
  assign _T_627 = StickySelects_5_io_outs_0; // @[MemPrimitives.scala 123:41:@3325.4]
  assign _T_629 = {_T_627,1'h1,1'h0}; // @[Cat.scala 30:58:@3327.4]
  assign _T_635 = StickySelects_6_io_outs_0; // @[MemPrimitives.scala 123:41:@3339.4]
  assign _T_637 = {_T_635,1'h1,1'h0}; // @[Cat.scala 30:58:@3341.4]
  assign _T_643 = StickySelects_7_io_outs_0; // @[MemPrimitives.scala 123:41:@3353.4]
  assign _T_645 = {_T_643,1'h1,1'h0}; // @[Cat.scala 30:58:@3355.4]
  assign _T_651 = StickySelects_8_io_outs_0; // @[MemPrimitives.scala 123:41:@3367.4]
  assign _T_653 = {_T_651,1'h1,1'h0}; // @[Cat.scala 30:58:@3369.4]
  assign _T_659 = StickySelects_9_io_outs_0; // @[MemPrimitives.scala 123:41:@3381.4]
  assign _T_661 = {_T_659,1'h1,1'h0}; // @[Cat.scala 30:58:@3383.4]
  assign _T_667 = StickySelects_10_io_outs_0; // @[MemPrimitives.scala 123:41:@3395.4]
  assign _T_669 = {_T_667,1'h1,1'h0}; // @[Cat.scala 30:58:@3397.4]
  assign _T_675 = StickySelects_11_io_outs_0; // @[MemPrimitives.scala 123:41:@3409.4]
  assign _T_677 = {_T_675,1'h1,1'h0}; // @[Cat.scala 30:58:@3411.4]
  assign _T_683 = StickySelects_12_io_outs_0; // @[MemPrimitives.scala 123:41:@3423.4]
  assign _T_685 = {_T_683,1'h1,1'h0}; // @[Cat.scala 30:58:@3425.4]
  assign _T_691 = StickySelects_13_io_outs_0; // @[MemPrimitives.scala 123:41:@3437.4]
  assign _T_693 = {_T_691,1'h1,1'h0}; // @[Cat.scala 30:58:@3439.4]
  assign _T_699 = StickySelects_14_io_outs_0; // @[MemPrimitives.scala 123:41:@3451.4]
  assign _T_701 = {_T_699,1'h1,1'h0}; // @[Cat.scala 30:58:@3453.4]
  assign _T_707 = StickySelects_15_io_outs_0; // @[MemPrimitives.scala 123:41:@3465.4]
  assign _T_709 = {_T_707,1'h1,1'h0}; // @[Cat.scala 30:58:@3467.4]
  assign io_rPort_15_output_0 = Mem1D_14_io_output; // @[MemPrimitives.scala 148:13:@3617.4]
  assign io_rPort_14_output_0 = Mem1D_9_io_output; // @[MemPrimitives.scala 148:13:@3608.4]
  assign io_rPort_13_output_0 = Mem1D_3_io_output; // @[MemPrimitives.scala 148:13:@3599.4]
  assign io_rPort_12_output_0 = Mem1D_8_io_output; // @[MemPrimitives.scala 148:13:@3590.4]
  assign io_rPort_11_output_0 = Mem1D_12_io_output; // @[MemPrimitives.scala 148:13:@3581.4]
  assign io_rPort_10_output_0 = Mem1D_5_io_output; // @[MemPrimitives.scala 148:13:@3572.4]
  assign io_rPort_9_output_0 = Mem1D_io_output; // @[MemPrimitives.scala 148:13:@3563.4]
  assign io_rPort_8_output_0 = Mem1D_6_io_output; // @[MemPrimitives.scala 148:13:@3554.4]
  assign io_rPort_7_output_0 = Mem1D_1_io_output; // @[MemPrimitives.scala 148:13:@3545.4]
  assign io_rPort_6_output_0 = Mem1D_11_io_output; // @[MemPrimitives.scala 148:13:@3536.4]
  assign io_rPort_5_output_0 = Mem1D_13_io_output; // @[MemPrimitives.scala 148:13:@3527.4]
  assign io_rPort_4_output_0 = Mem1D_4_io_output; // @[MemPrimitives.scala 148:13:@3518.4]
  assign io_rPort_3_output_0 = Mem1D_7_io_output; // @[MemPrimitives.scala 148:13:@3509.4]
  assign io_rPort_2_output_0 = Mem1D_10_io_output; // @[MemPrimitives.scala 148:13:@3500.4]
  assign io_rPort_1_output_0 = Mem1D_2_io_output; // @[MemPrimitives.scala 148:13:@3491.4]
  assign io_rPort_0_output_0 = Mem1D_15_io_output; // @[MemPrimitives.scala 148:13:@3482.4]
  assign Mem1D_clock = clock; // @[:@2835.4]
  assign Mem1D_reset = reset; // @[:@2836.4]
  assign Mem1D_io_r_ofs_0 = _T_589[0]; // @[MemPrimitives.scala 127:28:@3261.4]
  assign Mem1D_io_r_backpressure = _T_589[1]; // @[MemPrimitives.scala 128:32:@3262.4]
  assign Mem1D_io_w_ofs_0 = _T_461[0]; // @[MemPrimitives.scala 94:28:@3097.4]
  assign Mem1D_io_w_data_0 = _T_461[32:1]; // @[MemPrimitives.scala 95:29:@3098.4]
  assign Mem1D_io_w_en_0 = _T_461[33]; // @[MemPrimitives.scala 96:27:@3099.4]
  assign Mem1D_1_clock = clock; // @[:@2851.4]
  assign Mem1D_1_reset = reset; // @[:@2852.4]
  assign Mem1D_1_io_r_ofs_0 = _T_597[0]; // @[MemPrimitives.scala 127:28:@3275.4]
  assign Mem1D_1_io_r_backpressure = _T_597[1]; // @[MemPrimitives.scala 128:32:@3276.4]
  assign Mem1D_1_io_w_ofs_0 = _T_469[0]; // @[MemPrimitives.scala 94:28:@3107.4]
  assign Mem1D_1_io_w_data_0 = _T_469[32:1]; // @[MemPrimitives.scala 95:29:@3108.4]
  assign Mem1D_1_io_w_en_0 = _T_469[33]; // @[MemPrimitives.scala 96:27:@3109.4]
  assign Mem1D_2_clock = clock; // @[:@2867.4]
  assign Mem1D_2_reset = reset; // @[:@2868.4]
  assign Mem1D_2_io_r_ofs_0 = _T_605[0]; // @[MemPrimitives.scala 127:28:@3289.4]
  assign Mem1D_2_io_r_backpressure = _T_605[1]; // @[MemPrimitives.scala 128:32:@3290.4]
  assign Mem1D_2_io_w_ofs_0 = _T_477[0]; // @[MemPrimitives.scala 94:28:@3117.4]
  assign Mem1D_2_io_w_data_0 = _T_477[32:1]; // @[MemPrimitives.scala 95:29:@3118.4]
  assign Mem1D_2_io_w_en_0 = _T_477[33]; // @[MemPrimitives.scala 96:27:@3119.4]
  assign Mem1D_3_clock = clock; // @[:@2883.4]
  assign Mem1D_3_reset = reset; // @[:@2884.4]
  assign Mem1D_3_io_r_ofs_0 = _T_613[0]; // @[MemPrimitives.scala 127:28:@3303.4]
  assign Mem1D_3_io_r_backpressure = _T_613[1]; // @[MemPrimitives.scala 128:32:@3304.4]
  assign Mem1D_3_io_w_ofs_0 = _T_485[0]; // @[MemPrimitives.scala 94:28:@3127.4]
  assign Mem1D_3_io_w_data_0 = _T_485[32:1]; // @[MemPrimitives.scala 95:29:@3128.4]
  assign Mem1D_3_io_w_en_0 = _T_485[33]; // @[MemPrimitives.scala 96:27:@3129.4]
  assign Mem1D_4_clock = clock; // @[:@2899.4]
  assign Mem1D_4_reset = reset; // @[:@2900.4]
  assign Mem1D_4_io_r_ofs_0 = _T_621[0]; // @[MemPrimitives.scala 127:28:@3317.4]
  assign Mem1D_4_io_r_backpressure = _T_621[1]; // @[MemPrimitives.scala 128:32:@3318.4]
  assign Mem1D_4_io_w_ofs_0 = _T_493[0]; // @[MemPrimitives.scala 94:28:@3137.4]
  assign Mem1D_4_io_w_data_0 = _T_493[32:1]; // @[MemPrimitives.scala 95:29:@3138.4]
  assign Mem1D_4_io_w_en_0 = _T_493[33]; // @[MemPrimitives.scala 96:27:@3139.4]
  assign Mem1D_5_clock = clock; // @[:@2915.4]
  assign Mem1D_5_reset = reset; // @[:@2916.4]
  assign Mem1D_5_io_r_ofs_0 = _T_629[0]; // @[MemPrimitives.scala 127:28:@3331.4]
  assign Mem1D_5_io_r_backpressure = _T_629[1]; // @[MemPrimitives.scala 128:32:@3332.4]
  assign Mem1D_5_io_w_ofs_0 = _T_501[0]; // @[MemPrimitives.scala 94:28:@3147.4]
  assign Mem1D_5_io_w_data_0 = _T_501[32:1]; // @[MemPrimitives.scala 95:29:@3148.4]
  assign Mem1D_5_io_w_en_0 = _T_501[33]; // @[MemPrimitives.scala 96:27:@3149.4]
  assign Mem1D_6_clock = clock; // @[:@2931.4]
  assign Mem1D_6_reset = reset; // @[:@2932.4]
  assign Mem1D_6_io_r_ofs_0 = _T_637[0]; // @[MemPrimitives.scala 127:28:@3345.4]
  assign Mem1D_6_io_r_backpressure = _T_637[1]; // @[MemPrimitives.scala 128:32:@3346.4]
  assign Mem1D_6_io_w_ofs_0 = _T_509[0]; // @[MemPrimitives.scala 94:28:@3157.4]
  assign Mem1D_6_io_w_data_0 = _T_509[32:1]; // @[MemPrimitives.scala 95:29:@3158.4]
  assign Mem1D_6_io_w_en_0 = _T_509[33]; // @[MemPrimitives.scala 96:27:@3159.4]
  assign Mem1D_7_clock = clock; // @[:@2947.4]
  assign Mem1D_7_reset = reset; // @[:@2948.4]
  assign Mem1D_7_io_r_ofs_0 = _T_645[0]; // @[MemPrimitives.scala 127:28:@3359.4]
  assign Mem1D_7_io_r_backpressure = _T_645[1]; // @[MemPrimitives.scala 128:32:@3360.4]
  assign Mem1D_7_io_w_ofs_0 = _T_517[0]; // @[MemPrimitives.scala 94:28:@3167.4]
  assign Mem1D_7_io_w_data_0 = _T_517[32:1]; // @[MemPrimitives.scala 95:29:@3168.4]
  assign Mem1D_7_io_w_en_0 = _T_517[33]; // @[MemPrimitives.scala 96:27:@3169.4]
  assign Mem1D_8_clock = clock; // @[:@2963.4]
  assign Mem1D_8_reset = reset; // @[:@2964.4]
  assign Mem1D_8_io_r_ofs_0 = _T_653[0]; // @[MemPrimitives.scala 127:28:@3373.4]
  assign Mem1D_8_io_r_backpressure = _T_653[1]; // @[MemPrimitives.scala 128:32:@3374.4]
  assign Mem1D_8_io_w_ofs_0 = _T_525[0]; // @[MemPrimitives.scala 94:28:@3177.4]
  assign Mem1D_8_io_w_data_0 = _T_525[32:1]; // @[MemPrimitives.scala 95:29:@3178.4]
  assign Mem1D_8_io_w_en_0 = _T_525[33]; // @[MemPrimitives.scala 96:27:@3179.4]
  assign Mem1D_9_clock = clock; // @[:@2979.4]
  assign Mem1D_9_reset = reset; // @[:@2980.4]
  assign Mem1D_9_io_r_ofs_0 = _T_661[0]; // @[MemPrimitives.scala 127:28:@3387.4]
  assign Mem1D_9_io_r_backpressure = _T_661[1]; // @[MemPrimitives.scala 128:32:@3388.4]
  assign Mem1D_9_io_w_ofs_0 = _T_533[0]; // @[MemPrimitives.scala 94:28:@3187.4]
  assign Mem1D_9_io_w_data_0 = _T_533[32:1]; // @[MemPrimitives.scala 95:29:@3188.4]
  assign Mem1D_9_io_w_en_0 = _T_533[33]; // @[MemPrimitives.scala 96:27:@3189.4]
  assign Mem1D_10_clock = clock; // @[:@2995.4]
  assign Mem1D_10_reset = reset; // @[:@2996.4]
  assign Mem1D_10_io_r_ofs_0 = _T_669[0]; // @[MemPrimitives.scala 127:28:@3401.4]
  assign Mem1D_10_io_r_backpressure = _T_669[1]; // @[MemPrimitives.scala 128:32:@3402.4]
  assign Mem1D_10_io_w_ofs_0 = _T_541[0]; // @[MemPrimitives.scala 94:28:@3197.4]
  assign Mem1D_10_io_w_data_0 = _T_541[32:1]; // @[MemPrimitives.scala 95:29:@3198.4]
  assign Mem1D_10_io_w_en_0 = _T_541[33]; // @[MemPrimitives.scala 96:27:@3199.4]
  assign Mem1D_11_clock = clock; // @[:@3011.4]
  assign Mem1D_11_reset = reset; // @[:@3012.4]
  assign Mem1D_11_io_r_ofs_0 = _T_677[0]; // @[MemPrimitives.scala 127:28:@3415.4]
  assign Mem1D_11_io_r_backpressure = _T_677[1]; // @[MemPrimitives.scala 128:32:@3416.4]
  assign Mem1D_11_io_w_ofs_0 = _T_549[0]; // @[MemPrimitives.scala 94:28:@3207.4]
  assign Mem1D_11_io_w_data_0 = _T_549[32:1]; // @[MemPrimitives.scala 95:29:@3208.4]
  assign Mem1D_11_io_w_en_0 = _T_549[33]; // @[MemPrimitives.scala 96:27:@3209.4]
  assign Mem1D_12_clock = clock; // @[:@3027.4]
  assign Mem1D_12_reset = reset; // @[:@3028.4]
  assign Mem1D_12_io_r_ofs_0 = _T_685[0]; // @[MemPrimitives.scala 127:28:@3429.4]
  assign Mem1D_12_io_r_backpressure = _T_685[1]; // @[MemPrimitives.scala 128:32:@3430.4]
  assign Mem1D_12_io_w_ofs_0 = _T_557[0]; // @[MemPrimitives.scala 94:28:@3217.4]
  assign Mem1D_12_io_w_data_0 = _T_557[32:1]; // @[MemPrimitives.scala 95:29:@3218.4]
  assign Mem1D_12_io_w_en_0 = _T_557[33]; // @[MemPrimitives.scala 96:27:@3219.4]
  assign Mem1D_13_clock = clock; // @[:@3043.4]
  assign Mem1D_13_reset = reset; // @[:@3044.4]
  assign Mem1D_13_io_r_ofs_0 = _T_693[0]; // @[MemPrimitives.scala 127:28:@3443.4]
  assign Mem1D_13_io_r_backpressure = _T_693[1]; // @[MemPrimitives.scala 128:32:@3444.4]
  assign Mem1D_13_io_w_ofs_0 = _T_565[0]; // @[MemPrimitives.scala 94:28:@3227.4]
  assign Mem1D_13_io_w_data_0 = _T_565[32:1]; // @[MemPrimitives.scala 95:29:@3228.4]
  assign Mem1D_13_io_w_en_0 = _T_565[33]; // @[MemPrimitives.scala 96:27:@3229.4]
  assign Mem1D_14_clock = clock; // @[:@3059.4]
  assign Mem1D_14_reset = reset; // @[:@3060.4]
  assign Mem1D_14_io_r_ofs_0 = _T_701[0]; // @[MemPrimitives.scala 127:28:@3457.4]
  assign Mem1D_14_io_r_backpressure = _T_701[1]; // @[MemPrimitives.scala 128:32:@3458.4]
  assign Mem1D_14_io_w_ofs_0 = _T_573[0]; // @[MemPrimitives.scala 94:28:@3237.4]
  assign Mem1D_14_io_w_data_0 = _T_573[32:1]; // @[MemPrimitives.scala 95:29:@3238.4]
  assign Mem1D_14_io_w_en_0 = _T_573[33]; // @[MemPrimitives.scala 96:27:@3239.4]
  assign Mem1D_15_clock = clock; // @[:@3075.4]
  assign Mem1D_15_reset = reset; // @[:@3076.4]
  assign Mem1D_15_io_r_ofs_0 = _T_709[0]; // @[MemPrimitives.scala 127:28:@3471.4]
  assign Mem1D_15_io_r_backpressure = _T_709[1]; // @[MemPrimitives.scala 128:32:@3472.4]
  assign Mem1D_15_io_w_ofs_0 = _T_581[0]; // @[MemPrimitives.scala 94:28:@3247.4]
  assign Mem1D_15_io_w_data_0 = _T_581[32:1]; // @[MemPrimitives.scala 95:29:@3248.4]
  assign Mem1D_15_io_w_en_0 = _T_581[33]; // @[MemPrimitives.scala 96:27:@3249.4]
  assign StickySelects_io_ins_0 = io_rPort_9_en_0; // @[MemPrimitives.scala 122:60:@3254.4]
  assign StickySelects_1_io_ins_0 = io_rPort_7_en_0; // @[MemPrimitives.scala 122:60:@3268.4]
  assign StickySelects_2_io_ins_0 = io_rPort_1_en_0; // @[MemPrimitives.scala 122:60:@3282.4]
  assign StickySelects_3_io_ins_0 = io_rPort_13_en_0; // @[MemPrimitives.scala 122:60:@3296.4]
  assign StickySelects_4_io_ins_0 = io_rPort_4_en_0; // @[MemPrimitives.scala 122:60:@3310.4]
  assign StickySelects_5_io_ins_0 = io_rPort_10_en_0; // @[MemPrimitives.scala 122:60:@3324.4]
  assign StickySelects_6_io_ins_0 = io_rPort_8_en_0; // @[MemPrimitives.scala 122:60:@3338.4]
  assign StickySelects_7_io_ins_0 = io_rPort_3_en_0; // @[MemPrimitives.scala 122:60:@3352.4]
  assign StickySelects_8_io_ins_0 = io_rPort_12_en_0; // @[MemPrimitives.scala 122:60:@3366.4]
  assign StickySelects_9_io_ins_0 = io_rPort_14_en_0; // @[MemPrimitives.scala 122:60:@3380.4]
  assign StickySelects_10_io_ins_0 = io_rPort_2_en_0; // @[MemPrimitives.scala 122:60:@3394.4]
  assign StickySelects_11_io_ins_0 = io_rPort_6_en_0; // @[MemPrimitives.scala 122:60:@3408.4]
  assign StickySelects_12_io_ins_0 = io_rPort_11_en_0; // @[MemPrimitives.scala 122:60:@3422.4]
  assign StickySelects_13_io_ins_0 = io_rPort_5_en_0; // @[MemPrimitives.scala 122:60:@3436.4]
  assign StickySelects_14_io_ins_0 = io_rPort_15_en_0; // @[MemPrimitives.scala 122:60:@3450.4]
  assign StickySelects_15_io_ins_0 = io_rPort_0_en_0; // @[MemPrimitives.scala 122:60:@3464.4]
  assign RetimeWrapper_clock = clock; // @[:@3476.4]
  assign RetimeWrapper_reset = reset; // @[:@3477.4]
  assign RetimeWrapper_io_in = io_rPort_0_en_0; // @[package.scala 94:16:@3478.4]
  assign RetimeWrapper_1_clock = clock; // @[:@3485.4]
  assign RetimeWrapper_1_reset = reset; // @[:@3486.4]
  assign RetimeWrapper_1_io_in = io_rPort_1_en_0; // @[package.scala 94:16:@3487.4]
  assign RetimeWrapper_2_clock = clock; // @[:@3494.4]
  assign RetimeWrapper_2_reset = reset; // @[:@3495.4]
  assign RetimeWrapper_2_io_in = io_rPort_2_en_0; // @[package.scala 94:16:@3496.4]
  assign RetimeWrapper_3_clock = clock; // @[:@3503.4]
  assign RetimeWrapper_3_reset = reset; // @[:@3504.4]
  assign RetimeWrapper_3_io_in = io_rPort_3_en_0; // @[package.scala 94:16:@3505.4]
  assign RetimeWrapper_4_clock = clock; // @[:@3512.4]
  assign RetimeWrapper_4_reset = reset; // @[:@3513.4]
  assign RetimeWrapper_4_io_in = io_rPort_4_en_0; // @[package.scala 94:16:@3514.4]
  assign RetimeWrapper_5_clock = clock; // @[:@3521.4]
  assign RetimeWrapper_5_reset = reset; // @[:@3522.4]
  assign RetimeWrapper_5_io_in = io_rPort_5_en_0; // @[package.scala 94:16:@3523.4]
  assign RetimeWrapper_6_clock = clock; // @[:@3530.4]
  assign RetimeWrapper_6_reset = reset; // @[:@3531.4]
  assign RetimeWrapper_6_io_in = io_rPort_6_en_0; // @[package.scala 94:16:@3532.4]
  assign RetimeWrapper_7_clock = clock; // @[:@3539.4]
  assign RetimeWrapper_7_reset = reset; // @[:@3540.4]
  assign RetimeWrapper_7_io_in = io_rPort_7_en_0; // @[package.scala 94:16:@3541.4]
  assign RetimeWrapper_8_clock = clock; // @[:@3548.4]
  assign RetimeWrapper_8_reset = reset; // @[:@3549.4]
  assign RetimeWrapper_8_io_in = io_rPort_8_en_0; // @[package.scala 94:16:@3550.4]
  assign RetimeWrapper_9_clock = clock; // @[:@3557.4]
  assign RetimeWrapper_9_reset = reset; // @[:@3558.4]
  assign RetimeWrapper_9_io_in = io_rPort_9_en_0; // @[package.scala 94:16:@3559.4]
  assign RetimeWrapper_10_clock = clock; // @[:@3566.4]
  assign RetimeWrapper_10_reset = reset; // @[:@3567.4]
  assign RetimeWrapper_10_io_in = io_rPort_10_en_0; // @[package.scala 94:16:@3568.4]
  assign RetimeWrapper_11_clock = clock; // @[:@3575.4]
  assign RetimeWrapper_11_reset = reset; // @[:@3576.4]
  assign RetimeWrapper_11_io_in = io_rPort_11_en_0; // @[package.scala 94:16:@3577.4]
  assign RetimeWrapper_12_clock = clock; // @[:@3584.4]
  assign RetimeWrapper_12_reset = reset; // @[:@3585.4]
  assign RetimeWrapper_12_io_in = io_rPort_12_en_0; // @[package.scala 94:16:@3586.4]
  assign RetimeWrapper_13_clock = clock; // @[:@3593.4]
  assign RetimeWrapper_13_reset = reset; // @[:@3594.4]
  assign RetimeWrapper_13_io_in = io_rPort_13_en_0; // @[package.scala 94:16:@3595.4]
  assign RetimeWrapper_14_clock = clock; // @[:@3602.4]
  assign RetimeWrapper_14_reset = reset; // @[:@3603.4]
  assign RetimeWrapper_14_io_in = io_rPort_14_en_0; // @[package.scala 94:16:@3604.4]
  assign RetimeWrapper_15_clock = clock; // @[:@3611.4]
  assign RetimeWrapper_15_reset = reset; // @[:@3612.4]
  assign RetimeWrapper_15_io_in = io_rPort_15_en_0; // @[package.scala 94:16:@3613.4]
endmodule
module x294_outr_UnitPipe_sm( // @[:@3953.2]
  input   clock, // @[:@3954.4]
  input   reset, // @[:@3955.4]
  input   io_enable, // @[:@3956.4]
  output  io_done, // @[:@3956.4]
  input   io_parentAck, // @[:@3956.4]
  input   io_doneIn_0, // @[:@3956.4]
  input   io_doneIn_1, // @[:@3956.4]
  output  io_enableOut_0, // @[:@3956.4]
  output  io_enableOut_1, // @[:@3956.4]
  output  io_childAck_0, // @[:@3956.4]
  output  io_childAck_1, // @[:@3956.4]
  input   io_ctrCopyDone_0, // @[:@3956.4]
  input   io_ctrCopyDone_1 // @[:@3956.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@3959.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@3959.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@3959.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@3959.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@3959.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@3959.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@3962.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@3962.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@3962.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@3962.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@3962.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@3962.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@3965.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@3965.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@3965.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@3965.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@3965.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@3965.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@3968.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@3968.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@3968.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@3968.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@3968.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@3968.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@3997.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@3997.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@3997.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@3997.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@3997.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@3997.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@4000.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@4000.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@4000.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@4000.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@4000.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@4000.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@4041.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@4041.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@4041.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@4041.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@4041.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@4055.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@4055.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@4055.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@4055.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@4055.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@4073.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@4073.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@4073.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@4073.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@4073.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@4110.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@4110.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@4110.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@4110.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@4110.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@4124.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@4124.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@4124.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@4124.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@4124.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@4142.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@4142.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@4142.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@4142.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@4142.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@4189.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@4189.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@4189.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@4189.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@4189.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@4206.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@4206.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@4206.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@4206.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@4206.4]
  wire  allDone; // @[Controllers.scala 80:47:@3971.4]
  wire  _T_127; // @[Controllers.scala 165:35:@4025.4]
  wire  _T_129; // @[Controllers.scala 165:60:@4026.4]
  wire  _T_130; // @[Controllers.scala 165:58:@4027.4]
  wire  _T_132; // @[Controllers.scala 165:76:@4028.4]
  wire  _T_133; // @[Controllers.scala 165:74:@4029.4]
  wire  _T_137; // @[Controllers.scala 165:109:@4032.4]
  wire  _T_140; // @[Controllers.scala 165:141:@4034.4]
  wire  _T_148; // @[package.scala 96:25:@4046.4 package.scala 96:25:@4047.4]
  wire  _T_152; // @[Controllers.scala 167:54:@4049.4]
  wire  _T_153; // @[Controllers.scala 167:52:@4050.4]
  wire  _T_160; // @[package.scala 96:25:@4060.4 package.scala 96:25:@4061.4]
  wire  _T_178; // @[package.scala 96:25:@4078.4 package.scala 96:25:@4079.4]
  wire  _T_182; // @[Controllers.scala 169:67:@4081.4]
  wire  _T_183; // @[Controllers.scala 169:86:@4082.4]
  wire  _T_195; // @[Controllers.scala 165:35:@4094.4]
  wire  _T_197; // @[Controllers.scala 165:60:@4095.4]
  wire  _T_198; // @[Controllers.scala 165:58:@4096.4]
  wire  _T_200; // @[Controllers.scala 165:76:@4097.4]
  wire  _T_201; // @[Controllers.scala 165:74:@4098.4]
  wire  _T_205; // @[Controllers.scala 165:109:@4101.4]
  wire  _T_208; // @[Controllers.scala 165:141:@4103.4]
  wire  _T_216; // @[package.scala 96:25:@4115.4 package.scala 96:25:@4116.4]
  wire  _T_220; // @[Controllers.scala 167:54:@4118.4]
  wire  _T_221; // @[Controllers.scala 167:52:@4119.4]
  wire  _T_228; // @[package.scala 96:25:@4129.4 package.scala 96:25:@4130.4]
  wire  _T_246; // @[package.scala 96:25:@4147.4 package.scala 96:25:@4148.4]
  wire  _T_250; // @[Controllers.scala 169:67:@4150.4]
  wire  _T_251; // @[Controllers.scala 169:86:@4151.4]
  wire  _T_265; // @[Controllers.scala 213:68:@4167.4]
  wire  _T_267; // @[Controllers.scala 213:90:@4169.4]
  wire  _T_269; // @[Controllers.scala 213:132:@4171.4]
  wire  _T_273; // @[Controllers.scala 213:68:@4176.4]
  wire  _T_275; // @[Controllers.scala 213:90:@4178.4]
  wire  _T_282; // @[package.scala 100:49:@4184.4]
  reg  _T_285; // @[package.scala 48:56:@4185.4]
  reg [31:0] _RAND_0;
  wire  _T_286; // @[package.scala 100:41:@4187.4]
  reg  _T_299; // @[package.scala 48:56:@4203.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@3959.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@3962.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@3965.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@3968.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@3997.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@4000.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@4041.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@4055.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@4073.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@4110.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@4124.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@4142.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@4189.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@4206.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  assign allDone = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@3971.4]
  assign _T_127 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@4025.4]
  assign _T_129 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@4026.4]
  assign _T_130 = _T_127 & _T_129; // @[Controllers.scala 165:58:@4027.4]
  assign _T_132 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@4028.4]
  assign _T_133 = _T_130 & _T_132; // @[Controllers.scala 165:74:@4029.4]
  assign _T_137 = _T_133 & io_enable; // @[Controllers.scala 165:109:@4032.4]
  assign _T_140 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@4034.4]
  assign _T_148 = RetimeWrapper_io_out; // @[package.scala 96:25:@4046.4 package.scala 96:25:@4047.4]
  assign _T_152 = _T_148 == 1'h0; // @[Controllers.scala 167:54:@4049.4]
  assign _T_153 = io_doneIn_0 | _T_152; // @[Controllers.scala 167:52:@4050.4]
  assign _T_160 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@4060.4 package.scala 96:25:@4061.4]
  assign _T_178 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@4078.4 package.scala 96:25:@4079.4]
  assign _T_182 = _T_178 == 1'h0; // @[Controllers.scala 169:67:@4081.4]
  assign _T_183 = _T_182 & io_enable; // @[Controllers.scala 169:86:@4082.4]
  assign _T_195 = ~ iterDone_1_io_output; // @[Controllers.scala 165:35:@4094.4]
  assign _T_197 = io_doneIn_1 == 1'h0; // @[Controllers.scala 165:60:@4095.4]
  assign _T_198 = _T_195 & _T_197; // @[Controllers.scala 165:58:@4096.4]
  assign _T_200 = done_1_io_output == 1'h0; // @[Controllers.scala 165:76:@4097.4]
  assign _T_201 = _T_198 & _T_200; // @[Controllers.scala 165:74:@4098.4]
  assign _T_205 = _T_201 & io_enable; // @[Controllers.scala 165:109:@4101.4]
  assign _T_208 = io_ctrCopyDone_1 == 1'h0; // @[Controllers.scala 165:141:@4103.4]
  assign _T_216 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@4115.4 package.scala 96:25:@4116.4]
  assign _T_220 = _T_216 == 1'h0; // @[Controllers.scala 167:54:@4118.4]
  assign _T_221 = io_doneIn_1 | _T_220; // @[Controllers.scala 167:52:@4119.4]
  assign _T_228 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@4129.4 package.scala 96:25:@4130.4]
  assign _T_246 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@4147.4 package.scala 96:25:@4148.4]
  assign _T_250 = _T_246 == 1'h0; // @[Controllers.scala 169:67:@4150.4]
  assign _T_251 = _T_250 & io_enable; // @[Controllers.scala 169:86:@4151.4]
  assign _T_265 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@4167.4]
  assign _T_267 = _T_265 & _T_127; // @[Controllers.scala 213:90:@4169.4]
  assign _T_269 = ~ allDone; // @[Controllers.scala 213:132:@4171.4]
  assign _T_273 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@4176.4]
  assign _T_275 = _T_273 & _T_195; // @[Controllers.scala 213:90:@4178.4]
  assign _T_282 = allDone == 1'h0; // @[package.scala 100:49:@4184.4]
  assign _T_286 = allDone & _T_285; // @[package.scala 100:41:@4187.4]
  assign io_done = RetimeWrapper_7_io_out; // @[Controllers.scala 245:13:@4213.4]
  assign io_enableOut_0 = _T_267 & _T_269; // @[Controllers.scala 213:55:@4175.4]
  assign io_enableOut_1 = _T_275 & _T_269; // @[Controllers.scala 213:55:@4183.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@4164.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@4166.4]
  assign active_0_clock = clock; // @[:@3960.4]
  assign active_0_reset = reset; // @[:@3961.4]
  assign active_0_io_input_set = _T_137 & _T_140; // @[Controllers.scala 165:32:@4036.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@4040.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@3974.4]
  assign active_1_clock = clock; // @[:@3963.4]
  assign active_1_reset = reset; // @[:@3964.4]
  assign active_1_io_input_set = _T_205 & _T_208; // @[Controllers.scala 165:32:@4105.4]
  assign active_1_io_input_reset = io_ctrCopyDone_1 | io_parentAck; // @[Controllers.scala 166:34:@4109.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@3975.4]
  assign done_0_clock = clock; // @[:@3966.4]
  assign done_0_reset = reset; // @[:@3967.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_183; // @[Controllers.scala 169:30:@4086.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@3986.4 Controllers.scala 170:32:@4093.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@3976.4]
  assign done_1_clock = clock; // @[:@3969.4]
  assign done_1_reset = reset; // @[:@3970.4]
  assign done_1_io_input_set = io_ctrCopyDone_1 | _T_251; // @[Controllers.scala 169:30:@4155.4]
  assign done_1_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@3995.4 Controllers.scala 170:32:@4162.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@3977.4]
  assign iterDone_0_clock = clock; // @[:@3998.4]
  assign iterDone_0_reset = reset; // @[:@3999.4]
  assign iterDone_0_io_input_set = _T_153 & io_enable; // @[Controllers.scala 167:34:@4054.4]
  assign iterDone_0_io_input_reset = _T_160 | io_parentAck; // @[Controllers.scala 92:37:@4013.4 Controllers.scala 168:36:@4070.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@4003.4]
  assign iterDone_1_clock = clock; // @[:@4001.4]
  assign iterDone_1_reset = reset; // @[:@4002.4]
  assign iterDone_1_io_input_set = _T_221 & io_enable; // @[Controllers.scala 167:34:@4123.4]
  assign iterDone_1_io_input_reset = _T_228 | io_parentAck; // @[Controllers.scala 92:37:@4022.4 Controllers.scala 168:36:@4139.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@4004.4]
  assign RetimeWrapper_clock = clock; // @[:@4042.4]
  assign RetimeWrapper_reset = reset; // @[:@4043.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@4045.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@4044.4]
  assign RetimeWrapper_1_clock = clock; // @[:@4056.4]
  assign RetimeWrapper_1_reset = reset; // @[:@4057.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@4059.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@4058.4]
  assign RetimeWrapper_2_clock = clock; // @[:@4074.4]
  assign RetimeWrapper_2_reset = reset; // @[:@4075.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@4077.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@4076.4]
  assign RetimeWrapper_3_clock = clock; // @[:@4111.4]
  assign RetimeWrapper_3_reset = reset; // @[:@4112.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@4114.4]
  assign RetimeWrapper_3_io_in = 1'h1; // @[package.scala 94:16:@4113.4]
  assign RetimeWrapper_4_clock = clock; // @[:@4125.4]
  assign RetimeWrapper_4_reset = reset; // @[:@4126.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@4128.4]
  assign RetimeWrapper_4_io_in = io_doneIn_1; // @[package.scala 94:16:@4127.4]
  assign RetimeWrapper_5_clock = clock; // @[:@4143.4]
  assign RetimeWrapper_5_reset = reset; // @[:@4144.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@4146.4]
  assign RetimeWrapper_5_io_in = 1'h1; // @[package.scala 94:16:@4145.4]
  assign RetimeWrapper_6_clock = clock; // @[:@4190.4]
  assign RetimeWrapper_6_reset = reset; // @[:@4191.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@4193.4]
  assign RetimeWrapper_6_io_in = _T_286 | io_parentAck; // @[package.scala 94:16:@4192.4]
  assign RetimeWrapper_7_clock = clock; // @[:@4207.4]
  assign RetimeWrapper_7_reset = reset; // @[:@4208.4]
  assign RetimeWrapper_7_io_flow = io_enable; // @[package.scala 95:18:@4210.4]
  assign RetimeWrapper_7_io_in = allDone & _T_299; // @[package.scala 94:16:@4209.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_285 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_299 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_285 <= 1'h0;
    end else begin
      _T_285 <= _T_282;
    end
    if (reset) begin
      _T_299 <= 1'h0;
    end else begin
      _T_299 <= _T_282;
    end
  end
endmodule
module x280_inr_UnitPipe_sm( // @[:@4385.2]
  input   clock, // @[:@4386.4]
  input   reset, // @[:@4387.4]
  input   io_enable, // @[:@4388.4]
  output  io_done, // @[:@4388.4]
  output  io_doneLatch, // @[:@4388.4]
  input   io_ctrDone, // @[:@4388.4]
  output  io_datapathEn, // @[:@4388.4]
  output  io_ctrInc, // @[:@4388.4]
  input   io_parentAck, // @[:@4388.4]
  input   io_backpressure // @[:@4388.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@4390.4]
  wire  active_reset; // @[Controllers.scala 261:22:@4390.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@4390.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@4390.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@4390.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@4390.4]
  wire  done_clock; // @[Controllers.scala 262:20:@4393.4]
  wire  done_reset; // @[Controllers.scala 262:20:@4393.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@4393.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@4393.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@4393.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@4393.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@4447.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@4447.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@4447.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@4447.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@4447.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@4455.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@4455.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@4455.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@4455.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@4455.4]
  wire  _T_80; // @[Controllers.scala 264:48:@4398.4]
  wire  _T_81; // @[Controllers.scala 264:46:@4399.4]
  wire  _T_82; // @[Controllers.scala 264:62:@4400.4]
  wire  _T_83; // @[Controllers.scala 264:60:@4401.4]
  wire  _T_100; // @[package.scala 100:49:@4418.4]
  reg  _T_103; // @[package.scala 48:56:@4419.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 100:49:@4427.4]
  wire  _T_116; // @[Controllers.scala 283:41:@4435.4]
  wire  _T_117; // @[Controllers.scala 283:59:@4436.4]
  wire  _T_119; // @[Controllers.scala 284:37:@4439.4]
  reg  _T_125; // @[package.scala 48:56:@4443.4]
  reg [31:0] _RAND_1;
  reg  _T_142; // @[Controllers.scala 291:31:@4465.4]
  reg [31:0] _RAND_2;
  reg  _T_149; // @[package.scala 48:56:@4468.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:41:@4470.4]
  wire  _T_152; // @[Controllers.scala 292:61:@4471.4]
  wire  _T_153; // @[Controllers.scala 292:24:@4472.4]
  SRFF active ( // @[Controllers.scala 261:22:@4390.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@4393.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@4447.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@4455.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@4398.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@4399.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@4400.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@4401.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@4418.4]
  assign _T_108 = done_io_output == 1'h0; // @[package.scala 100:49:@4427.4]
  assign _T_116 = active_io_output & _T_82; // @[Controllers.scala 283:41:@4435.4]
  assign _T_117 = _T_116 & io_enable; // @[Controllers.scala 283:59:@4436.4]
  assign _T_119 = active_io_output & io_enable; // @[Controllers.scala 284:37:@4439.4]
  assign _T_150 = done_io_output & _T_149; // @[package.scala 100:41:@4470.4]
  assign _T_152 = _T_150 ? 1'h1 : _T_142; // @[Controllers.scala 292:61:@4471.4]
  assign _T_153 = io_parentAck ? 1'h0 : _T_152; // @[Controllers.scala 292:24:@4472.4]
  assign io_done = done_io_output & _T_125; // @[Controllers.scala 287:13:@4446.4]
  assign io_doneLatch = _T_142; // @[Controllers.scala 293:18:@4474.4]
  assign io_datapathEn = _T_117 & io_backpressure; // @[Controllers.scala 283:21:@4438.4]
  assign io_ctrInc = _T_119 & io_backpressure; // @[Controllers.scala 284:17:@4441.4]
  assign active_clock = clock; // @[:@4391.4]
  assign active_reset = reset; // @[:@4392.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@4403.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@4407.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@4408.4]
  assign done_clock = clock; // @[:@4394.4]
  assign done_reset = reset; // @[:@4395.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@4423.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@4416.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@4417.4]
  assign RetimeWrapper_clock = clock; // @[:@4448.4]
  assign RetimeWrapper_reset = reset; // @[:@4449.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@4451.4]
  assign RetimeWrapper_io_in = 1'h0; // @[package.scala 94:16:@4450.4]
  assign RetimeWrapper_1_clock = clock; // @[:@4456.4]
  assign RetimeWrapper_1_reset = reset; // @[:@4457.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@4459.4]
  assign RetimeWrapper_1_io_in = io_ctrDone; // @[package.scala 94:16:@4458.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_125 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_142 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_149 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_125 <= 1'h0;
    end else begin
      _T_125 <= _T_108;
    end
    if (reset) begin
      _T_142 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_142 <= 1'h0;
      end else begin
        if (_T_150) begin
          _T_142 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_149 <= 1'h0;
    end else begin
      _T_149 <= _T_108;
    end
  end
endmodule
module x280_inr_UnitPipe_kernelx280_inr_UnitPipe_concrete1( // @[:@4548.2]
  output        io_in_x274_valid, // @[:@4551.4]
  output [63:0] io_in_x274_bits_addr, // @[:@4551.4]
  output [31:0] io_in_x274_bits_size, // @[:@4551.4]
  input  [63:0] io_in_x254_in_number, // @[:@4551.4]
  input         io_sigsIn_backpressure, // @[:@4551.4]
  input         io_sigsIn_datapathEn, // @[:@4551.4]
  input         io_rr // @[:@4551.4]
);
  wire [96:0] x277_tuple; // @[Cat.scala 30:58:@4565.4]
  wire  _T_135; // @[implicits.scala 55:10:@4568.4]
  assign x277_tuple = {33'h100000040,io_in_x254_in_number}; // @[Cat.scala 30:58:@4565.4]
  assign _T_135 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 55:10:@4568.4]
  assign io_in_x274_valid = _T_135 & io_sigsIn_backpressure; // @[sm_x280_inr_UnitPipe.scala 64:18:@4571.4]
  assign io_in_x274_bits_addr = x277_tuple[63:0]; // @[sm_x280_inr_UnitPipe.scala 65:22:@4573.4]
  assign io_in_x274_bits_size = x277_tuple[95:64]; // @[sm_x280_inr_UnitPipe.scala 66:22:@4575.4]
endmodule
module SingleCounter_1( // @[:@4615.2]
  input         clock, // @[:@4616.4]
  input         reset, // @[:@4617.4]
  input         io_input_reset, // @[:@4618.4]
  input         io_input_enable, // @[:@4618.4]
  output [31:0] io_output_count_0, // @[:@4618.4]
  output        io_output_oobs_0, // @[:@4618.4]
  output        io_output_done // @[:@4618.4]
);
  wire  bases_0_clock; // @[Counter.scala 253:53:@4631.4]
  wire  bases_0_reset; // @[Counter.scala 253:53:@4631.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 253:53:@4631.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 253:53:@4631.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 253:53:@4631.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 253:53:@4631.4]
  wire  SRFF_clock; // @[Counter.scala 255:22:@4647.4]
  wire  SRFF_reset; // @[Counter.scala 255:22:@4647.4]
  wire  SRFF_io_input_set; // @[Counter.scala 255:22:@4647.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 255:22:@4647.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 255:22:@4647.4]
  wire  SRFF_io_output; // @[Counter.scala 255:22:@4647.4]
  wire  _T_36; // @[Counter.scala 256:45:@4650.4]
  wire [31:0] _T_48; // @[Counter.scala 279:52:@4675.4]
  wire [32:0] _T_50; // @[Counter.scala 283:33:@4676.4]
  wire [31:0] _T_51; // @[Counter.scala 283:33:@4677.4]
  wire [31:0] _T_52; // @[Counter.scala 283:33:@4678.4]
  wire  _T_57; // @[Counter.scala 285:18:@4680.4]
  wire [31:0] _T_68; // @[Counter.scala 291:115:@4688.4]
  wire [31:0] _T_71; // @[Counter.scala 291:152:@4691.4]
  wire [31:0] _T_72; // @[Counter.scala 291:74:@4692.4]
  wire  _T_75; // @[Counter.scala 314:102:@4696.4]
  wire  _T_77; // @[Counter.scala 314:130:@4697.4]
  FF bases_0 ( // @[Counter.scala 253:53:@4631.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 255:22:@4647.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 256:45:@4650.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 279:52:@4675.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@4676.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@4677.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 283:33:@4678.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh10); // @[Counter.scala 285:18:@4680.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 291:115:@4688.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 291:152:@4691.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 291:74:@4692.4]
  assign _T_75 = $signed(_T_48) < $signed(32'sh0); // @[Counter.scala 314:102:@4696.4]
  assign _T_77 = $signed(_T_48) >= $signed(32'sh10); // @[Counter.scala 314:130:@4697.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 296:28:@4695.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 314:60:@4699.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 325:20:@4701.4]
  assign bases_0_clock = clock; // @[:@4632.4]
  assign bases_0_reset = reset; // @[:@4633.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 291:31:@4694.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 273:27:@4673.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 276:29:@4674.4]
  assign SRFF_clock = clock; // @[:@4648.4]
  assign SRFF_reset = reset; // @[:@4649.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 256:23:@4652.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 257:25:@4654.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 258:30:@4655.4]
endmodule
module x283_ctrchain( // @[:@4706.2]
  input         clock, // @[:@4707.4]
  input         reset, // @[:@4708.4]
  input         io_input_reset, // @[:@4709.4]
  input         io_input_enable, // @[:@4709.4]
  output [31:0] io_output_counts_0, // @[:@4709.4]
  output        io_output_oobs_0, // @[:@4709.4]
  output        io_output_done // @[:@4709.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 505:46:@4711.4]
  wire  ctrs_0_reset; // @[Counter.scala 505:46:@4711.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 505:46:@4711.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 505:46:@4711.4]
  wire [31:0] ctrs_0_io_output_count_0; // @[Counter.scala 505:46:@4711.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 505:46:@4711.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 505:46:@4711.4]
  reg  wasDone; // @[Counter.scala 534:24:@4720.4]
  reg [31:0] _RAND_0;
  wire  _T_45; // @[Counter.scala 538:69:@4726.4]
  wire  _T_47; // @[Counter.scala 538:80:@4727.4]
  reg  doneLatch; // @[Counter.scala 542:26:@4732.4]
  reg [31:0] _RAND_1;
  wire  _T_54; // @[Counter.scala 543:48:@4733.4]
  wire  _T_55; // @[Counter.scala 543:19:@4734.4]
  SingleCounter_1 ctrs_0 ( // @[Counter.scala 505:46:@4711.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done)
  );
  assign _T_45 = io_input_enable & ctrs_0_io_output_done; // @[Counter.scala 538:69:@4726.4]
  assign _T_47 = wasDone == 1'h0; // @[Counter.scala 538:80:@4727.4]
  assign _T_54 = ctrs_0_io_output_done ? 1'h1 : doneLatch; // @[Counter.scala 543:48:@4733.4]
  assign _T_55 = io_input_reset ? 1'h0 : _T_54; // @[Counter.scala 543:19:@4734.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 549:32:@4736.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 550:30:@4738.4]
  assign io_output_done = _T_45 & _T_47; // @[Counter.scala 538:18:@4729.4]
  assign ctrs_0_clock = clock; // @[:@4712.4]
  assign ctrs_0_reset = reset; // @[:@4713.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 512:24:@4717.4]
  assign ctrs_0_io_input_enable = io_input_enable; // @[Counter.scala 516:33:@4718.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= ctrs_0_io_output_done;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (ctrs_0_io_output_done) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module x293_inr_Foreach_sm( // @[:@4926.2]
  input   clock, // @[:@4927.4]
  input   reset, // @[:@4928.4]
  input   io_enable, // @[:@4929.4]
  output  io_done, // @[:@4929.4]
  output  io_doneLatch, // @[:@4929.4]
  input   io_ctrDone, // @[:@4929.4]
  output  io_datapathEn, // @[:@4929.4]
  output  io_ctrInc, // @[:@4929.4]
  output  io_ctrRst, // @[:@4929.4]
  input   io_parentAck, // @[:@4929.4]
  input   io_break // @[:@4929.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@4931.4]
  wire  active_reset; // @[Controllers.scala 261:22:@4931.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@4931.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@4931.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@4931.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@4931.4]
  wire  done_clock; // @[Controllers.scala 262:20:@4934.4]
  wire  done_reset; // @[Controllers.scala 262:20:@4934.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@4934.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@4934.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@4934.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@4934.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@4968.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@4968.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@4968.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@4968.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@4990.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@4990.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@4990.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@4990.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@5002.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@5002.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@5002.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@5002.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@5002.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@5010.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@5010.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@5010.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@5010.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@5010.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@5026.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@5026.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@5026.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@5026.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@5026.4]
  wire  _T_80; // @[Controllers.scala 264:48:@4939.4]
  wire  _T_81; // @[Controllers.scala 264:46:@4940.4]
  wire  _T_82; // @[Controllers.scala 264:62:@4941.4]
  wire  _T_100; // @[package.scala 100:49:@4959.4]
  reg  _T_103; // @[package.scala 48:56:@4960.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@4973.4 package.scala 96:25:@4974.4]
  wire  _T_110; // @[package.scala 100:49:@4975.4]
  reg  _T_113; // @[package.scala 48:56:@4976.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@4978.4]
  wire  _T_118; // @[Controllers.scala 283:41:@4983.4]
  wire  _T_124; // @[package.scala 96:25:@4995.4 package.scala 96:25:@4996.4]
  wire  _T_126; // @[package.scala 100:49:@4997.4]
  reg  _T_129; // @[package.scala 48:56:@4998.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@5020.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@5022.4]
  reg  _T_153; // @[package.scala 48:56:@5023.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@5031.4 package.scala 96:25:@5032.4]
  wire  _T_158; // @[Controllers.scala 292:61:@5033.4]
  wire  _T_159; // @[Controllers.scala 292:24:@5034.4]
  SRFF active ( // @[Controllers.scala 261:22:@4931.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@4934.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_37 RetimeWrapper ( // @[package.scala 93:22:@4968.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_37 RetimeWrapper_1 ( // @[package.scala 93:22:@4990.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@5002.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@5010.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@5026.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@4939.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@4940.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@4941.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@4959.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@4973.4 package.scala 96:25:@4974.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@4975.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@4978.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@4983.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@4995.4 package.scala 96:25:@4996.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@4997.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@5022.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@5031.4 package.scala 96:25:@5032.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@5033.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@5034.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@5001.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@5036.4]
  assign io_datapathEn = _T_118 & io_enable; // @[Controllers.scala 283:21:@4986.4]
  assign io_ctrInc = active_io_output & io_enable; // @[Controllers.scala 284:17:@4989.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@4981.4]
  assign active_clock = clock; // @[:@4932.4]
  assign active_reset = reset; // @[:@4933.4]
  assign active_io_input_set = _T_81 & _T_82; // @[Controllers.scala 264:23:@4944.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@4948.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@4949.4]
  assign done_clock = clock; // @[:@4935.4]
  assign done_reset = reset; // @[:@4936.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@4964.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@4957.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@4958.4]
  assign RetimeWrapper_clock = clock; // @[:@4969.4]
  assign RetimeWrapper_reset = reset; // @[:@4970.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@4971.4]
  assign RetimeWrapper_1_clock = clock; // @[:@4991.4]
  assign RetimeWrapper_1_reset = reset; // @[:@4992.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@4993.4]
  assign RetimeWrapper_2_clock = clock; // @[:@5003.4]
  assign RetimeWrapper_2_reset = reset; // @[:@5004.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@5006.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@5005.4]
  assign RetimeWrapper_3_clock = clock; // @[:@5011.4]
  assign RetimeWrapper_3_reset = reset; // @[:@5012.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@5014.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@5013.4]
  assign RetimeWrapper_4_clock = clock; // @[:@5027.4]
  assign RetimeWrapper_4_reset = reset; // @[:@5028.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@5030.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@5029.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module fix2fixBox( // @[:@5142.2]
  input  [31:0] io_a, // @[:@5145.4]
  output [31:0] io_b // @[:@5145.4]
);
  assign io_b = io_a; // @[Converter.scala 95:38:@5155.4]
endmodule
module _( // @[:@5157.2]
  input  [31:0] io_b, // @[:@5160.4]
  output [31:0] io_result // @[:@5160.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@5165.4]
  wire [31:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@5165.4]
  fix2fixBox fix2fixBox ( // @[BigIPZynq.scala 219:30:@5165.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 706:17:@5173.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@5168.4]
endmodule
module x293_inr_Foreach_kernelx293_inr_Foreach_concrete1( // @[:@5335.2]
  input         clock, // @[:@5336.4]
  input         reset, // @[:@5337.4]
  output        io_in_x275_ready, // @[:@5338.4]
  input  [31:0] io_in_x275_bits_rdata_0, // @[:@5338.4]
  output [4:0]  io_in_x273_a_0_wPort_0_banks_0, // @[:@5338.4]
  output        io_in_x273_a_0_wPort_0_ofs_0, // @[:@5338.4]
  output [31:0] io_in_x273_a_0_wPort_0_data_0, // @[:@5338.4]
  output        io_in_x273_a_0_wPort_0_en_0, // @[:@5338.4]
  input         io_sigsIn_datapathEn, // @[:@5338.4]
  input         io_sigsIn_break, // @[:@5338.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@5338.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@5338.4]
  input         io_rr // @[:@5338.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@5440.4]
  wire [31:0] __io_result; // @[Math.scala 709:24:@5440.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@5454.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@5454.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@5454.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@5454.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@5454.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@5485.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@5485.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@5485.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@5485.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@5485.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@5494.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@5494.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@5494.4]
  wire [31:0] RetimeWrapper_2_io_in; // @[package.scala 93:22:@5494.4]
  wire [31:0] RetimeWrapper_2_io_out; // @[package.scala 93:22:@5494.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@5503.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@5503.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@5503.4]
  wire [31:0] RetimeWrapper_3_io_in; // @[package.scala 93:22:@5503.4]
  wire [31:0] RetimeWrapper_3_io_out; // @[package.scala 93:22:@5503.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@5514.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@5514.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@5514.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@5514.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@5514.4]
  wire  b285; // @[sm_x293_inr_Foreach.scala 61:18:@5448.4]
  wire [31:0] b284_number; // @[Math.scala 712:22:@5445.4 Math.scala 713:14:@5446.4]
  wire [31:0] _T_1078; // @[Math.scala 406:49:@5468.4]
  wire [31:0] _T_1080; // @[Math.scala 406:56:@5470.4]
  wire [31:0] _T_1081; // @[Math.scala 406:56:@5471.4]
  wire  _T_1087; // @[FixedPoint.scala 50:25:@5477.4]
  wire [3:0] _T_1091; // @[Bitwise.scala 72:12:@5479.4]
  wire [27:0] _T_1092; // @[FixedPoint.scala 18:52:@5480.4]
  wire  _T_1103; // @[sm_x293_inr_Foreach.scala 83:96:@5511.4]
  wire  _T_1107; // @[package.scala 96:25:@5519.4 package.scala 96:25:@5520.4]
  wire  _T_1109; // @[implicits.scala 55:10:@5521.4]
  wire  _T_1110; // @[sm_x293_inr_Foreach.scala 83:113:@5522.4]
  wire  _T_1112; // @[sm_x293_inr_Foreach.scala 83:200:@5524.4]
  wire  x458_b285_D1; // @[package.scala 96:25:@5490.4 package.scala 96:25:@5491.4]
  wire [31:0] x459_x456_D1_number; // @[package.scala 96:25:@5499.4 package.scala 96:25:@5500.4]
  wire [31:0] x460_x289_D1_number; // @[package.scala 96:25:@5508.4 package.scala 96:25:@5509.4]
  _ _ ( // @[Math.scala 709:24:@5440.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@5454.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@5485.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_2 ( // @[package.scala 93:22:@5494.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_3 ( // @[package.scala 93:22:@5503.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@5514.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign b285 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x293_inr_Foreach.scala 61:18:@5448.4]
  assign b284_number = __io_result; // @[Math.scala 712:22:@5445.4 Math.scala 713:14:@5446.4]
  assign _T_1078 = $signed(b284_number); // @[Math.scala 406:49:@5468.4]
  assign _T_1080 = $signed(_T_1078) & $signed(32'shf); // @[Math.scala 406:56:@5470.4]
  assign _T_1081 = $signed(_T_1080); // @[Math.scala 406:56:@5471.4]
  assign _T_1087 = b284_number[31]; // @[FixedPoint.scala 50:25:@5477.4]
  assign _T_1091 = _T_1087 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12:@5479.4]
  assign _T_1092 = b284_number[31:4]; // @[FixedPoint.scala 18:52:@5480.4]
  assign _T_1103 = ~ io_sigsIn_break; // @[sm_x293_inr_Foreach.scala 83:96:@5511.4]
  assign _T_1107 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@5519.4 package.scala 96:25:@5520.4]
  assign _T_1109 = io_rr ? _T_1107 : 1'h0; // @[implicits.scala 55:10:@5521.4]
  assign _T_1110 = _T_1103 & _T_1109; // @[sm_x293_inr_Foreach.scala 83:113:@5522.4]
  assign _T_1112 = _T_1110 & _T_1103; // @[sm_x293_inr_Foreach.scala 83:200:@5524.4]
  assign x458_b285_D1 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@5490.4 package.scala 96:25:@5491.4]
  assign x459_x456_D1_number = RetimeWrapper_2_io_out; // @[package.scala 96:25:@5499.4 package.scala 96:25:@5500.4]
  assign x460_x289_D1_number = RetimeWrapper_3_io_out; // @[package.scala 96:25:@5508.4 package.scala 96:25:@5509.4]
  assign io_in_x275_ready = b285 & io_sigsIn_datapathEn; // @[sm_x293_inr_Foreach.scala 63:18:@5451.4]
  assign io_in_x273_a_0_wPort_0_banks_0 = x459_x456_D1_number[4:0]; // @[MemInterfaceType.scala 88:58:@5527.4]
  assign io_in_x273_a_0_wPort_0_ofs_0 = x460_x289_D1_number[0]; // @[MemInterfaceType.scala 89:54:@5528.4]
  assign io_in_x273_a_0_wPort_0_data_0 = RetimeWrapper_io_out; // @[MemInterfaceType.scala 90:56:@5529.4]
  assign io_in_x273_a_0_wPort_0_en_0 = _T_1112 & x458_b285_D1; // @[MemInterfaceType.scala 93:57:@5531.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 710:17:@5443.4]
  assign RetimeWrapper_clock = clock; // @[:@5455.4]
  assign RetimeWrapper_reset = reset; // @[:@5456.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@5458.4]
  assign RetimeWrapper_io_in = io_in_x275_bits_rdata_0; // @[package.scala 94:16:@5457.4]
  assign RetimeWrapper_1_clock = clock; // @[:@5486.4]
  assign RetimeWrapper_1_reset = reset; // @[:@5487.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@5489.4]
  assign RetimeWrapper_1_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@5488.4]
  assign RetimeWrapper_2_clock = clock; // @[:@5495.4]
  assign RetimeWrapper_2_reset = reset; // @[:@5496.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@5498.4]
  assign RetimeWrapper_2_io_in = $unsigned(_T_1081); // @[package.scala 94:16:@5497.4]
  assign RetimeWrapper_3_clock = clock; // @[:@5504.4]
  assign RetimeWrapper_3_reset = reset; // @[:@5505.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@5507.4]
  assign RetimeWrapper_3_io_in = {_T_1091,_T_1092}; // @[package.scala 94:16:@5506.4]
  assign RetimeWrapper_4_clock = clock; // @[:@5515.4]
  assign RetimeWrapper_4_reset = reset; // @[:@5516.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@5518.4]
  assign RetimeWrapper_4_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@5517.4]
endmodule
module x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1( // @[:@5533.2]
  input         clock, // @[:@5534.4]
  input         reset, // @[:@5535.4]
  output [4:0]  io_in_x273_a_0_wPort_0_banks_0, // @[:@5536.4]
  output        io_in_x273_a_0_wPort_0_ofs_0, // @[:@5536.4]
  output [31:0] io_in_x273_a_0_wPort_0_data_0, // @[:@5536.4]
  output        io_in_x273_a_0_wPort_0_en_0, // @[:@5536.4]
  input  [63:0] io_in_x254_in_number, // @[:@5536.4]
  input         io_in_x274_ready, // @[:@5536.4]
  output        io_in_x274_valid, // @[:@5536.4]
  output [63:0] io_in_x274_bits_addr, // @[:@5536.4]
  output [31:0] io_in_x274_bits_size, // @[:@5536.4]
  output        io_in_x275_ready, // @[:@5536.4]
  input         io_in_x275_valid, // @[:@5536.4]
  input  [31:0] io_in_x275_bits_rdata_0, // @[:@5536.4]
  input         io_sigsIn_smEnableOuts_0, // @[:@5536.4]
  input         io_sigsIn_smEnableOuts_1, // @[:@5536.4]
  input         io_sigsIn_smChildAcks_0, // @[:@5536.4]
  input         io_sigsIn_smChildAcks_1, // @[:@5536.4]
  output        io_sigsOut_smDoneIn_0, // @[:@5536.4]
  output        io_sigsOut_smDoneIn_1, // @[:@5536.4]
  output        io_sigsOut_smCtrCopyDone_0, // @[:@5536.4]
  output        io_sigsOut_smCtrCopyDone_1, // @[:@5536.4]
  input         io_rr // @[:@5536.4]
);
  wire  x280_inr_UnitPipe_sm_clock; // @[sm_x280_inr_UnitPipe.scala 32:18:@5673.4]
  wire  x280_inr_UnitPipe_sm_reset; // @[sm_x280_inr_UnitPipe.scala 32:18:@5673.4]
  wire  x280_inr_UnitPipe_sm_io_enable; // @[sm_x280_inr_UnitPipe.scala 32:18:@5673.4]
  wire  x280_inr_UnitPipe_sm_io_done; // @[sm_x280_inr_UnitPipe.scala 32:18:@5673.4]
  wire  x280_inr_UnitPipe_sm_io_doneLatch; // @[sm_x280_inr_UnitPipe.scala 32:18:@5673.4]
  wire  x280_inr_UnitPipe_sm_io_ctrDone; // @[sm_x280_inr_UnitPipe.scala 32:18:@5673.4]
  wire  x280_inr_UnitPipe_sm_io_datapathEn; // @[sm_x280_inr_UnitPipe.scala 32:18:@5673.4]
  wire  x280_inr_UnitPipe_sm_io_ctrInc; // @[sm_x280_inr_UnitPipe.scala 32:18:@5673.4]
  wire  x280_inr_UnitPipe_sm_io_parentAck; // @[sm_x280_inr_UnitPipe.scala 32:18:@5673.4]
  wire  x280_inr_UnitPipe_sm_io_backpressure; // @[sm_x280_inr_UnitPipe.scala 32:18:@5673.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@5730.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@5730.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@5730.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@5730.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@5730.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@5738.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@5738.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@5738.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@5738.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@5738.4]
  wire  x280_inr_UnitPipe_kernelx280_inr_UnitPipe_concrete1_io_in_x274_valid; // @[sm_x280_inr_UnitPipe.scala 68:24:@5765.4]
  wire [63:0] x280_inr_UnitPipe_kernelx280_inr_UnitPipe_concrete1_io_in_x274_bits_addr; // @[sm_x280_inr_UnitPipe.scala 68:24:@5765.4]
  wire [31:0] x280_inr_UnitPipe_kernelx280_inr_UnitPipe_concrete1_io_in_x274_bits_size; // @[sm_x280_inr_UnitPipe.scala 68:24:@5765.4]
  wire [63:0] x280_inr_UnitPipe_kernelx280_inr_UnitPipe_concrete1_io_in_x254_in_number; // @[sm_x280_inr_UnitPipe.scala 68:24:@5765.4]
  wire  x280_inr_UnitPipe_kernelx280_inr_UnitPipe_concrete1_io_sigsIn_backpressure; // @[sm_x280_inr_UnitPipe.scala 68:24:@5765.4]
  wire  x280_inr_UnitPipe_kernelx280_inr_UnitPipe_concrete1_io_sigsIn_datapathEn; // @[sm_x280_inr_UnitPipe.scala 68:24:@5765.4]
  wire  x280_inr_UnitPipe_kernelx280_inr_UnitPipe_concrete1_io_rr; // @[sm_x280_inr_UnitPipe.scala 68:24:@5765.4]
  wire  x283_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@5831.4]
  wire  x283_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@5831.4]
  wire  x283_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@5831.4]
  wire  x283_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@5831.4]
  wire [31:0] x283_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@5831.4]
  wire  x283_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@5831.4]
  wire  x283_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@5831.4]
  wire  x293_inr_Foreach_sm_clock; // @[sm_x293_inr_Foreach.scala 32:18:@5883.4]
  wire  x293_inr_Foreach_sm_reset; // @[sm_x293_inr_Foreach.scala 32:18:@5883.4]
  wire  x293_inr_Foreach_sm_io_enable; // @[sm_x293_inr_Foreach.scala 32:18:@5883.4]
  wire  x293_inr_Foreach_sm_io_done; // @[sm_x293_inr_Foreach.scala 32:18:@5883.4]
  wire  x293_inr_Foreach_sm_io_doneLatch; // @[sm_x293_inr_Foreach.scala 32:18:@5883.4]
  wire  x293_inr_Foreach_sm_io_ctrDone; // @[sm_x293_inr_Foreach.scala 32:18:@5883.4]
  wire  x293_inr_Foreach_sm_io_datapathEn; // @[sm_x293_inr_Foreach.scala 32:18:@5883.4]
  wire  x293_inr_Foreach_sm_io_ctrInc; // @[sm_x293_inr_Foreach.scala 32:18:@5883.4]
  wire  x293_inr_Foreach_sm_io_ctrRst; // @[sm_x293_inr_Foreach.scala 32:18:@5883.4]
  wire  x293_inr_Foreach_sm_io_parentAck; // @[sm_x293_inr_Foreach.scala 32:18:@5883.4]
  wire  x293_inr_Foreach_sm_io_break; // @[sm_x293_inr_Foreach.scala 32:18:@5883.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@5911.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@5911.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@5911.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@5911.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@5911.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@5951.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@5951.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@5951.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@5951.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@5951.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@5959.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@5959.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@5959.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@5959.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@5959.4]
  wire  x293_inr_Foreach_kernelx293_inr_Foreach_concrete1_clock; // @[sm_x293_inr_Foreach.scala 85:24:@5991.4]
  wire  x293_inr_Foreach_kernelx293_inr_Foreach_concrete1_reset; // @[sm_x293_inr_Foreach.scala 85:24:@5991.4]
  wire  x293_inr_Foreach_kernelx293_inr_Foreach_concrete1_io_in_x275_ready; // @[sm_x293_inr_Foreach.scala 85:24:@5991.4]
  wire [31:0] x293_inr_Foreach_kernelx293_inr_Foreach_concrete1_io_in_x275_bits_rdata_0; // @[sm_x293_inr_Foreach.scala 85:24:@5991.4]
  wire [4:0] x293_inr_Foreach_kernelx293_inr_Foreach_concrete1_io_in_x273_a_0_wPort_0_banks_0; // @[sm_x293_inr_Foreach.scala 85:24:@5991.4]
  wire  x293_inr_Foreach_kernelx293_inr_Foreach_concrete1_io_in_x273_a_0_wPort_0_ofs_0; // @[sm_x293_inr_Foreach.scala 85:24:@5991.4]
  wire [31:0] x293_inr_Foreach_kernelx293_inr_Foreach_concrete1_io_in_x273_a_0_wPort_0_data_0; // @[sm_x293_inr_Foreach.scala 85:24:@5991.4]
  wire  x293_inr_Foreach_kernelx293_inr_Foreach_concrete1_io_in_x273_a_0_wPort_0_en_0; // @[sm_x293_inr_Foreach.scala 85:24:@5991.4]
  wire  x293_inr_Foreach_kernelx293_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x293_inr_Foreach.scala 85:24:@5991.4]
  wire  x293_inr_Foreach_kernelx293_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x293_inr_Foreach.scala 85:24:@5991.4]
  wire [31:0] x293_inr_Foreach_kernelx293_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x293_inr_Foreach.scala 85:24:@5991.4]
  wire  x293_inr_Foreach_kernelx293_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x293_inr_Foreach.scala 85:24:@5991.4]
  wire  x293_inr_Foreach_kernelx293_inr_Foreach_concrete1_io_rr; // @[sm_x293_inr_Foreach.scala 85:24:@5991.4]
  wire  _T_1125; // @[package.scala 100:49:@5701.4]
  reg  _T_1128; // @[package.scala 48:56:@5702.4]
  reg [31:0] _RAND_0;
  wire  _T_1141; // @[package.scala 96:25:@5735.4 package.scala 96:25:@5736.4]
  wire  _T_1147; // @[package.scala 96:25:@5743.4 package.scala 96:25:@5744.4]
  wire  _T_1150; // @[SpatialBlocks.scala 110:93:@5746.4]
  wire  _T_1218; // @[package.scala 96:25:@5916.4 package.scala 96:25:@5917.4]
  wire  x293_inr_Foreach_sigsIn_forwardpressure; // @[sm_x294_outr_UnitPipe.scala 86:54:@5922.4]
  wire  _T_1232; // @[package.scala 96:25:@5956.4 package.scala 96:25:@5957.4]
  wire  _T_1238; // @[package.scala 96:25:@5964.4 package.scala 96:25:@5965.4]
  wire  _T_1241; // @[SpatialBlocks.scala 110:93:@5967.4]
  wire  x293_inr_Foreach_sigsIn_baseEn; // @[SpatialBlocks.scala 110:90:@5968.4]
  wire  _T_1243; // @[SpatialBlocks.scala 128:36:@5976.4]
  wire  _T_1244; // @[SpatialBlocks.scala 128:78:@5977.4]
  wire  _T_1249; // @[SpatialBlocks.scala 130:61:@5986.4]
  x280_inr_UnitPipe_sm x280_inr_UnitPipe_sm ( // @[sm_x280_inr_UnitPipe.scala 32:18:@5673.4]
    .clock(x280_inr_UnitPipe_sm_clock),
    .reset(x280_inr_UnitPipe_sm_reset),
    .io_enable(x280_inr_UnitPipe_sm_io_enable),
    .io_done(x280_inr_UnitPipe_sm_io_done),
    .io_doneLatch(x280_inr_UnitPipe_sm_io_doneLatch),
    .io_ctrDone(x280_inr_UnitPipe_sm_io_ctrDone),
    .io_datapathEn(x280_inr_UnitPipe_sm_io_datapathEn),
    .io_ctrInc(x280_inr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x280_inr_UnitPipe_sm_io_parentAck),
    .io_backpressure(x280_inr_UnitPipe_sm_io_backpressure)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@5730.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@5738.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x280_inr_UnitPipe_kernelx280_inr_UnitPipe_concrete1 x280_inr_UnitPipe_kernelx280_inr_UnitPipe_concrete1 ( // @[sm_x280_inr_UnitPipe.scala 68:24:@5765.4]
    .io_in_x274_valid(x280_inr_UnitPipe_kernelx280_inr_UnitPipe_concrete1_io_in_x274_valid),
    .io_in_x274_bits_addr(x280_inr_UnitPipe_kernelx280_inr_UnitPipe_concrete1_io_in_x274_bits_addr),
    .io_in_x274_bits_size(x280_inr_UnitPipe_kernelx280_inr_UnitPipe_concrete1_io_in_x274_bits_size),
    .io_in_x254_in_number(x280_inr_UnitPipe_kernelx280_inr_UnitPipe_concrete1_io_in_x254_in_number),
    .io_sigsIn_backpressure(x280_inr_UnitPipe_kernelx280_inr_UnitPipe_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x280_inr_UnitPipe_kernelx280_inr_UnitPipe_concrete1_io_sigsIn_datapathEn),
    .io_rr(x280_inr_UnitPipe_kernelx280_inr_UnitPipe_concrete1_io_rr)
  );
  x283_ctrchain x283_ctrchain ( // @[SpatialBlocks.scala 37:22:@5831.4]
    .clock(x283_ctrchain_clock),
    .reset(x283_ctrchain_reset),
    .io_input_reset(x283_ctrchain_io_input_reset),
    .io_input_enable(x283_ctrchain_io_input_enable),
    .io_output_counts_0(x283_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x283_ctrchain_io_output_oobs_0),
    .io_output_done(x283_ctrchain_io_output_done)
  );
  x293_inr_Foreach_sm x293_inr_Foreach_sm ( // @[sm_x293_inr_Foreach.scala 32:18:@5883.4]
    .clock(x293_inr_Foreach_sm_clock),
    .reset(x293_inr_Foreach_sm_reset),
    .io_enable(x293_inr_Foreach_sm_io_enable),
    .io_done(x293_inr_Foreach_sm_io_done),
    .io_doneLatch(x293_inr_Foreach_sm_io_doneLatch),
    .io_ctrDone(x293_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x293_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x293_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x293_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x293_inr_Foreach_sm_io_parentAck),
    .io_break(x293_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@5911.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@5951.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@5959.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  x293_inr_Foreach_kernelx293_inr_Foreach_concrete1 x293_inr_Foreach_kernelx293_inr_Foreach_concrete1 ( // @[sm_x293_inr_Foreach.scala 85:24:@5991.4]
    .clock(x293_inr_Foreach_kernelx293_inr_Foreach_concrete1_clock),
    .reset(x293_inr_Foreach_kernelx293_inr_Foreach_concrete1_reset),
    .io_in_x275_ready(x293_inr_Foreach_kernelx293_inr_Foreach_concrete1_io_in_x275_ready),
    .io_in_x275_bits_rdata_0(x293_inr_Foreach_kernelx293_inr_Foreach_concrete1_io_in_x275_bits_rdata_0),
    .io_in_x273_a_0_wPort_0_banks_0(x293_inr_Foreach_kernelx293_inr_Foreach_concrete1_io_in_x273_a_0_wPort_0_banks_0),
    .io_in_x273_a_0_wPort_0_ofs_0(x293_inr_Foreach_kernelx293_inr_Foreach_concrete1_io_in_x273_a_0_wPort_0_ofs_0),
    .io_in_x273_a_0_wPort_0_data_0(x293_inr_Foreach_kernelx293_inr_Foreach_concrete1_io_in_x273_a_0_wPort_0_data_0),
    .io_in_x273_a_0_wPort_0_en_0(x293_inr_Foreach_kernelx293_inr_Foreach_concrete1_io_in_x273_a_0_wPort_0_en_0),
    .io_sigsIn_datapathEn(x293_inr_Foreach_kernelx293_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x293_inr_Foreach_kernelx293_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_0(x293_inr_Foreach_kernelx293_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x293_inr_Foreach_kernelx293_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_rr(x293_inr_Foreach_kernelx293_inr_Foreach_concrete1_io_rr)
  );
  assign _T_1125 = x280_inr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@5701.4]
  assign _T_1141 = RetimeWrapper_io_out; // @[package.scala 96:25:@5735.4 package.scala 96:25:@5736.4]
  assign _T_1147 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@5743.4 package.scala 96:25:@5744.4]
  assign _T_1150 = ~ _T_1147; // @[SpatialBlocks.scala 110:93:@5746.4]
  assign _T_1218 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@5916.4 package.scala 96:25:@5917.4]
  assign x293_inr_Foreach_sigsIn_forwardpressure = io_in_x275_valid | x293_inr_Foreach_sm_io_doneLatch; // @[sm_x294_outr_UnitPipe.scala 86:54:@5922.4]
  assign _T_1232 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@5956.4 package.scala 96:25:@5957.4]
  assign _T_1238 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@5964.4 package.scala 96:25:@5965.4]
  assign _T_1241 = ~ _T_1238; // @[SpatialBlocks.scala 110:93:@5967.4]
  assign x293_inr_Foreach_sigsIn_baseEn = _T_1232 & _T_1241; // @[SpatialBlocks.scala 110:90:@5968.4]
  assign _T_1243 = x293_inr_Foreach_sm_io_datapathEn; // @[SpatialBlocks.scala 128:36:@5976.4]
  assign _T_1244 = ~ x293_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 128:78:@5977.4]
  assign _T_1249 = x293_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 130:61:@5986.4]
  assign io_in_x273_a_0_wPort_0_banks_0 = x293_inr_Foreach_kernelx293_inr_Foreach_concrete1_io_in_x273_a_0_wPort_0_banks_0; // @[MemInterfaceType.scala 67:44:@6121.4]
  assign io_in_x273_a_0_wPort_0_ofs_0 = x293_inr_Foreach_kernelx293_inr_Foreach_concrete1_io_in_x273_a_0_wPort_0_ofs_0; // @[MemInterfaceType.scala 67:44:@6120.4]
  assign io_in_x273_a_0_wPort_0_data_0 = x293_inr_Foreach_kernelx293_inr_Foreach_concrete1_io_in_x273_a_0_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@6119.4]
  assign io_in_x273_a_0_wPort_0_en_0 = x293_inr_Foreach_kernelx293_inr_Foreach_concrete1_io_in_x273_a_0_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@6115.4]
  assign io_in_x274_valid = x280_inr_UnitPipe_kernelx280_inr_UnitPipe_concrete1_io_in_x274_valid; // @[sm_x280_inr_UnitPipe.scala 48:23:@5802.4]
  assign io_in_x274_bits_addr = x280_inr_UnitPipe_kernelx280_inr_UnitPipe_concrete1_io_in_x274_bits_addr; // @[sm_x280_inr_UnitPipe.scala 48:23:@5801.4]
  assign io_in_x274_bits_size = x280_inr_UnitPipe_kernelx280_inr_UnitPipe_concrete1_io_in_x274_bits_size; // @[sm_x280_inr_UnitPipe.scala 48:23:@5800.4]
  assign io_in_x275_ready = x293_inr_Foreach_kernelx293_inr_Foreach_concrete1_io_in_x275_ready; // @[sm_x293_inr_Foreach.scala 48:23:@6114.4]
  assign io_sigsOut_smDoneIn_0 = x280_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 127:53:@5753.4]
  assign io_sigsOut_smDoneIn_1 = x293_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 127:53:@5974.4]
  assign io_sigsOut_smCtrCopyDone_0 = x280_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 139:125:@5764.4]
  assign io_sigsOut_smCtrCopyDone_1 = x293_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 139:125:@5990.4]
  assign x280_inr_UnitPipe_sm_clock = clock; // @[:@5674.4]
  assign x280_inr_UnitPipe_sm_reset = reset; // @[:@5675.4]
  assign x280_inr_UnitPipe_sm_io_enable = _T_1141 & _T_1150; // @[SpatialBlocks.scala 112:18:@5750.4]
  assign x280_inr_UnitPipe_sm_io_ctrDone = x280_inr_UnitPipe_sm_io_ctrInc & _T_1128; // @[sm_x294_outr_UnitPipe.scala 71:39:@5705.4]
  assign x280_inr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 114:21:@5752.4]
  assign x280_inr_UnitPipe_sm_io_backpressure = io_in_x274_ready | x280_inr_UnitPipe_sm_io_doneLatch; // @[SpatialBlocks.scala 105:24:@5724.4]
  assign RetimeWrapper_clock = clock; // @[:@5731.4]
  assign RetimeWrapper_reset = reset; // @[:@5732.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@5734.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@5733.4]
  assign RetimeWrapper_1_clock = clock; // @[:@5739.4]
  assign RetimeWrapper_1_reset = reset; // @[:@5740.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@5742.4]
  assign RetimeWrapper_1_io_in = x280_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@5741.4]
  assign x280_inr_UnitPipe_kernelx280_inr_UnitPipe_concrete1_io_in_x254_in_number = io_in_x254_in_number; // @[sm_x280_inr_UnitPipe.scala 49:26:@5804.4]
  assign x280_inr_UnitPipe_kernelx280_inr_UnitPipe_concrete1_io_sigsIn_backpressure = io_in_x274_ready | x280_inr_UnitPipe_sm_io_doneLatch; // @[sm_x280_inr_UnitPipe.scala 72:22:@5819.4]
  assign x280_inr_UnitPipe_kernelx280_inr_UnitPipe_concrete1_io_sigsIn_datapathEn = x280_inr_UnitPipe_sm_io_datapathEn; // @[sm_x280_inr_UnitPipe.scala 72:22:@5817.4]
  assign x280_inr_UnitPipe_kernelx280_inr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x280_inr_UnitPipe.scala 71:18:@5805.4]
  assign x283_ctrchain_clock = clock; // @[:@5832.4]
  assign x283_ctrchain_reset = reset; // @[:@5833.4]
  assign x283_ctrchain_io_input_reset = x293_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 130:103:@5989.4]
  assign x283_ctrchain_io_input_enable = _T_1249 & x293_inr_Foreach_sigsIn_forwardpressure; // @[SpatialBlocks.scala 104:75:@5944.4 SpatialBlocks.scala 130:45:@5988.4]
  assign x293_inr_Foreach_sm_clock = clock; // @[:@5884.4]
  assign x293_inr_Foreach_sm_reset = reset; // @[:@5885.4]
  assign x293_inr_Foreach_sm_io_enable = x293_inr_Foreach_sigsIn_baseEn & x293_inr_Foreach_sigsIn_forwardpressure; // @[SpatialBlocks.scala 112:18:@5971.4]
  assign x293_inr_Foreach_sm_io_ctrDone = io_rr ? _T_1218 : 1'h0; // @[sm_x294_outr_UnitPipe.scala 84:38:@5919.4]
  assign x293_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 114:21:@5973.4]
  assign x293_inr_Foreach_sm_io_break = 1'h0; // @[sm_x294_outr_UnitPipe.scala 88:36:@5925.4]
  assign RetimeWrapper_2_clock = clock; // @[:@5912.4]
  assign RetimeWrapper_2_reset = reset; // @[:@5913.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@5915.4]
  assign RetimeWrapper_2_io_in = x283_ctrchain_io_output_done; // @[package.scala 94:16:@5914.4]
  assign RetimeWrapper_3_clock = clock; // @[:@5952.4]
  assign RetimeWrapper_3_reset = reset; // @[:@5953.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@5955.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@5954.4]
  assign RetimeWrapper_4_clock = clock; // @[:@5960.4]
  assign RetimeWrapper_4_reset = reset; // @[:@5961.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@5963.4]
  assign RetimeWrapper_4_io_in = x293_inr_Foreach_sm_io_done; // @[package.scala 94:16:@5962.4]
  assign x293_inr_Foreach_kernelx293_inr_Foreach_concrete1_clock = clock; // @[:@5992.4]
  assign x293_inr_Foreach_kernelx293_inr_Foreach_concrete1_reset = reset; // @[:@5993.4]
  assign x293_inr_Foreach_kernelx293_inr_Foreach_concrete1_io_in_x275_bits_rdata_0 = io_in_x275_bits_rdata_0; // @[sm_x293_inr_Foreach.scala 48:23:@6112.4]
  assign x293_inr_Foreach_kernelx293_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_1243 & _T_1244; // @[sm_x293_inr_Foreach.scala 89:22:@6134.4]
  assign x293_inr_Foreach_kernelx293_inr_Foreach_concrete1_io_sigsIn_break = x293_inr_Foreach_sm_io_break; // @[sm_x293_inr_Foreach.scala 89:22:@6132.4]
  assign x293_inr_Foreach_kernelx293_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = x283_ctrchain_io_output_counts_0; // @[sm_x293_inr_Foreach.scala 89:22:@6127.4]
  assign x293_inr_Foreach_kernelx293_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x283_ctrchain_io_output_oobs_0; // @[sm_x293_inr_Foreach.scala 89:22:@6126.4]
  assign x293_inr_Foreach_kernelx293_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x293_inr_Foreach.scala 88:18:@6122.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1128 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_1128 <= 1'h0;
    end else begin
      _T_1128 <= _T_1125;
    end
  end
endmodule
module RetimeWrapper_80( // @[:@6187.2]
  input   clock, // @[:@6188.4]
  input   reset, // @[:@6189.4]
  input   io_in, // @[:@6190.4]
  output  io_out // @[:@6190.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@6192.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@6192.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@6192.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@6192.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@6192.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@6192.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@6192.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@6205.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@6204.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@6203.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@6202.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@6201.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@6199.4]
endmodule
module x343_inr_UnitPipe_sm( // @[:@6335.2]
  input   clock, // @[:@6336.4]
  input   reset, // @[:@6337.4]
  input   io_enable, // @[:@6338.4]
  output  io_done, // @[:@6338.4]
  input   io_ctrDone, // @[:@6338.4]
  output  io_datapathEn, // @[:@6338.4]
  output  io_ctrInc, // @[:@6338.4]
  input   io_parentAck, // @[:@6338.4]
  input   io_break // @[:@6338.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@6340.4]
  wire  active_reset; // @[Controllers.scala 261:22:@6340.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@6340.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@6340.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@6340.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@6340.4]
  wire  done_clock; // @[Controllers.scala 262:20:@6343.4]
  wire  done_reset; // @[Controllers.scala 262:20:@6343.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@6343.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@6343.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@6343.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@6343.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@6377.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@6377.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@6377.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@6377.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@6399.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@6399.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@6399.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@6399.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@6411.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@6411.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@6411.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@6411.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@6411.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@6419.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@6419.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@6419.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@6419.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@6419.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@6435.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@6435.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@6435.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@6435.4]
  wire  _T_80; // @[Controllers.scala 264:48:@6348.4]
  wire  _T_81; // @[Controllers.scala 264:46:@6349.4]
  wire  _T_82; // @[Controllers.scala 264:62:@6350.4]
  wire  _T_100; // @[package.scala 100:49:@6368.4]
  reg  _T_103; // @[package.scala 48:56:@6369.4]
  reg [31:0] _RAND_0;
  wire  _T_118; // @[Controllers.scala 283:41:@6392.4]
  wire  _T_124; // @[package.scala 96:25:@6404.4 package.scala 96:25:@6405.4]
  wire  _T_126; // @[package.scala 100:49:@6406.4]
  reg  _T_129; // @[package.scala 48:56:@6407.4]
  reg [31:0] _RAND_1;
  wire  _T_150; // @[package.scala 100:49:@6431.4]
  reg  _T_153; // @[package.scala 48:56:@6432.4]
  reg [31:0] _RAND_2;
  SRFF active ( // @[Controllers.scala 261:22:@6340.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@6343.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_80 RetimeWrapper ( // @[package.scala 93:22:@6377.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_80 RetimeWrapper_1 ( // @[package.scala 93:22:@6399.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@6411.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@6419.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_37 RetimeWrapper_4 ( // @[package.scala 93:22:@6435.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@6348.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@6349.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@6350.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@6368.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@6392.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@6404.4 package.scala 96:25:@6405.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@6406.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@6431.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@6410.4]
  assign io_datapathEn = _T_118 & io_enable; // @[Controllers.scala 283:21:@6395.4]
  assign io_ctrInc = active_io_output & io_enable; // @[Controllers.scala 284:17:@6398.4]
  assign active_clock = clock; // @[:@6341.4]
  assign active_reset = reset; // @[:@6342.4]
  assign active_io_input_set = _T_81 & _T_82; // @[Controllers.scala 264:23:@6353.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@6357.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@6358.4]
  assign done_clock = clock; // @[:@6344.4]
  assign done_reset = reset; // @[:@6345.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@6373.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@6366.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@6367.4]
  assign RetimeWrapper_clock = clock; // @[:@6378.4]
  assign RetimeWrapper_reset = reset; // @[:@6379.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@6380.4]
  assign RetimeWrapper_1_clock = clock; // @[:@6400.4]
  assign RetimeWrapper_1_reset = reset; // @[:@6401.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@6402.4]
  assign RetimeWrapper_2_clock = clock; // @[:@6412.4]
  assign RetimeWrapper_2_reset = reset; // @[:@6413.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@6415.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@6414.4]
  assign RetimeWrapper_3_clock = clock; // @[:@6420.4]
  assign RetimeWrapper_3_reset = reset; // @[:@6421.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@6423.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@6422.4]
  assign RetimeWrapper_4_clock = clock; // @[:@6436.4]
  assign RetimeWrapper_4_reset = reset; // @[:@6437.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@6438.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_129 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_153 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1( // @[:@7031.2]
  input         clock, // @[:@7032.4]
  input         reset, // @[:@7033.4]
  output        io_in_x269_argOut_port_0_valid, // @[:@7034.4]
  output [63:0] io_in_x269_argOut_port_0_bits, // @[:@7034.4]
  output        io_in_x257_argOut_port_0_valid, // @[:@7034.4]
  output [63:0] io_in_x257_argOut_port_0_bits, // @[:@7034.4]
  output        io_in_x261_argOut_port_0_valid, // @[:@7034.4]
  output [63:0] io_in_x261_argOut_port_0_bits, // @[:@7034.4]
  output        io_in_x265_argOut_port_0_valid, // @[:@7034.4]
  output [63:0] io_in_x265_argOut_port_0_bits, // @[:@7034.4]
  output        io_in_x270_argOut_port_0_valid, // @[:@7034.4]
  output [63:0] io_in_x270_argOut_port_0_bits, // @[:@7034.4]
  output        io_in_x260_argOut_port_0_valid, // @[:@7034.4]
  output [63:0] io_in_x260_argOut_port_0_bits, // @[:@7034.4]
  output        io_in_x256_argOut_port_0_valid, // @[:@7034.4]
  output [63:0] io_in_x256_argOut_port_0_bits, // @[:@7034.4]
  output        io_in_x266_argOut_port_0_valid, // @[:@7034.4]
  output [63:0] io_in_x266_argOut_port_0_bits, // @[:@7034.4]
  output        io_in_x264_argOut_port_0_valid, // @[:@7034.4]
  output [63:0] io_in_x264_argOut_port_0_bits, // @[:@7034.4]
  output        io_in_x259_argOut_port_0_valid, // @[:@7034.4]
  output [63:0] io_in_x259_argOut_port_0_bits, // @[:@7034.4]
  output        io_in_x267_argOut_port_0_valid, // @[:@7034.4]
  output [63:0] io_in_x267_argOut_port_0_bits, // @[:@7034.4]
  output        io_in_x255_argOut_port_0_valid, // @[:@7034.4]
  output [63:0] io_in_x255_argOut_port_0_bits, // @[:@7034.4]
  output        io_in_x263_argOut_port_0_valid, // @[:@7034.4]
  output [63:0] io_in_x263_argOut_port_0_bits, // @[:@7034.4]
  output        io_in_x258_argOut_port_0_valid, // @[:@7034.4]
  output [63:0] io_in_x258_argOut_port_0_bits, // @[:@7034.4]
  output        io_in_x262_argOut_port_0_valid, // @[:@7034.4]
  output [63:0] io_in_x262_argOut_port_0_bits, // @[:@7034.4]
  output        io_in_x273_a_0_rPort_15_en_0, // @[:@7034.4]
  input  [31:0] io_in_x273_a_0_rPort_15_output_0, // @[:@7034.4]
  output        io_in_x273_a_0_rPort_14_en_0, // @[:@7034.4]
  input  [31:0] io_in_x273_a_0_rPort_14_output_0, // @[:@7034.4]
  output        io_in_x273_a_0_rPort_13_en_0, // @[:@7034.4]
  input  [31:0] io_in_x273_a_0_rPort_13_output_0, // @[:@7034.4]
  output        io_in_x273_a_0_rPort_12_en_0, // @[:@7034.4]
  input  [31:0] io_in_x273_a_0_rPort_12_output_0, // @[:@7034.4]
  output        io_in_x273_a_0_rPort_11_en_0, // @[:@7034.4]
  input  [31:0] io_in_x273_a_0_rPort_11_output_0, // @[:@7034.4]
  output        io_in_x273_a_0_rPort_10_en_0, // @[:@7034.4]
  input  [31:0] io_in_x273_a_0_rPort_10_output_0, // @[:@7034.4]
  output        io_in_x273_a_0_rPort_9_en_0, // @[:@7034.4]
  input  [31:0] io_in_x273_a_0_rPort_9_output_0, // @[:@7034.4]
  output        io_in_x273_a_0_rPort_8_en_0, // @[:@7034.4]
  input  [31:0] io_in_x273_a_0_rPort_8_output_0, // @[:@7034.4]
  output        io_in_x273_a_0_rPort_7_en_0, // @[:@7034.4]
  input  [31:0] io_in_x273_a_0_rPort_7_output_0, // @[:@7034.4]
  output        io_in_x273_a_0_rPort_6_en_0, // @[:@7034.4]
  input  [31:0] io_in_x273_a_0_rPort_6_output_0, // @[:@7034.4]
  output        io_in_x273_a_0_rPort_5_en_0, // @[:@7034.4]
  input  [31:0] io_in_x273_a_0_rPort_5_output_0, // @[:@7034.4]
  output        io_in_x273_a_0_rPort_4_en_0, // @[:@7034.4]
  input  [31:0] io_in_x273_a_0_rPort_4_output_0, // @[:@7034.4]
  output        io_in_x273_a_0_rPort_3_en_0, // @[:@7034.4]
  input  [31:0] io_in_x273_a_0_rPort_3_output_0, // @[:@7034.4]
  output        io_in_x273_a_0_rPort_2_en_0, // @[:@7034.4]
  input  [31:0] io_in_x273_a_0_rPort_2_output_0, // @[:@7034.4]
  output        io_in_x273_a_0_rPort_1_en_0, // @[:@7034.4]
  input  [31:0] io_in_x273_a_0_rPort_1_output_0, // @[:@7034.4]
  output        io_in_x273_a_0_rPort_0_en_0, // @[:@7034.4]
  input  [31:0] io_in_x273_a_0_rPort_0_output_0, // @[:@7034.4]
  output        io_in_x268_argOut_port_0_valid, // @[:@7034.4]
  output [63:0] io_in_x268_argOut_port_0_bits, // @[:@7034.4]
  input         io_sigsIn_datapathEn, // @[:@7034.4]
  input         io_sigsIn_break, // @[:@7034.4]
  input         io_rr // @[:@7034.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@7219.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@7219.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@7219.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@7219.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@7252.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@7252.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@7252.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@7252.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@7285.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@7285.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@7285.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@7285.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@7318.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@7318.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@7318.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@7318.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@7351.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@7351.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@7351.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@7351.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@7384.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@7384.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@7384.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@7384.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@7417.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@7417.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@7417.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@7417.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@7450.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@7450.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@7450.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@7450.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@7483.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@7483.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@7483.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@7483.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@7516.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@7516.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@7516.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@7516.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@7549.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@7549.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@7549.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@7549.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@7582.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@7582.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@7582.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@7582.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@7615.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@7615.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@7615.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@7615.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@7648.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@7648.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@7648.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@7648.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@7681.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@7681.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@7681.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@7681.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@7714.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@7714.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@7714.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@7714.4]
  wire  _T_1357; // @[sm_x343_inr_UnitPipe.scala 140:124:@7201.4]
  wire  _T_1361; // @[implicits.scala 55:10:@7204.4]
  wire  _T_1366; // @[FixedPoint.scala 50:25:@7214.4]
  wire [31:0] _T_1370; // @[Bitwise.scala 72:12:@7216.4]
  wire  _T_1400; // @[FixedPoint.scala 50:25:@7247.4]
  wire [31:0] _T_1404; // @[Bitwise.scala 72:12:@7249.4]
  wire  _T_1434; // @[FixedPoint.scala 50:25:@7280.4]
  wire [31:0] _T_1438; // @[Bitwise.scala 72:12:@7282.4]
  wire  _T_1468; // @[FixedPoint.scala 50:25:@7313.4]
  wire [31:0] _T_1472; // @[Bitwise.scala 72:12:@7315.4]
  wire  _T_1502; // @[FixedPoint.scala 50:25:@7346.4]
  wire [31:0] _T_1506; // @[Bitwise.scala 72:12:@7348.4]
  wire  _T_1536; // @[FixedPoint.scala 50:25:@7379.4]
  wire [31:0] _T_1540; // @[Bitwise.scala 72:12:@7381.4]
  wire  _T_1570; // @[FixedPoint.scala 50:25:@7412.4]
  wire [31:0] _T_1574; // @[Bitwise.scala 72:12:@7414.4]
  wire  _T_1604; // @[FixedPoint.scala 50:25:@7445.4]
  wire [31:0] _T_1608; // @[Bitwise.scala 72:12:@7447.4]
  wire  _T_1638; // @[FixedPoint.scala 50:25:@7478.4]
  wire [31:0] _T_1642; // @[Bitwise.scala 72:12:@7480.4]
  wire  _T_1672; // @[FixedPoint.scala 50:25:@7511.4]
  wire [31:0] _T_1676; // @[Bitwise.scala 72:12:@7513.4]
  wire  _T_1706; // @[FixedPoint.scala 50:25:@7544.4]
  wire [31:0] _T_1710; // @[Bitwise.scala 72:12:@7546.4]
  wire  _T_1740; // @[FixedPoint.scala 50:25:@7577.4]
  wire [31:0] _T_1744; // @[Bitwise.scala 72:12:@7579.4]
  wire  _T_1774; // @[FixedPoint.scala 50:25:@7610.4]
  wire [31:0] _T_1778; // @[Bitwise.scala 72:12:@7612.4]
  wire  _T_1808; // @[FixedPoint.scala 50:25:@7643.4]
  wire [31:0] _T_1812; // @[Bitwise.scala 72:12:@7645.4]
  wire  _T_1842; // @[FixedPoint.scala 50:25:@7676.4]
  wire [31:0] _T_1846; // @[Bitwise.scala 72:12:@7678.4]
  wire  _T_1876; // @[FixedPoint.scala 50:25:@7709.4]
  wire [31:0] _T_1880; // @[Bitwise.scala 72:12:@7711.4]
  RetimeWrapper_37 RetimeWrapper ( // @[package.scala 93:22:@7219.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_37 RetimeWrapper_1 ( // @[package.scala 93:22:@7252.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_37 RetimeWrapper_2 ( // @[package.scala 93:22:@7285.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_37 RetimeWrapper_3 ( // @[package.scala 93:22:@7318.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_37 RetimeWrapper_4 ( // @[package.scala 93:22:@7351.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_37 RetimeWrapper_5 ( // @[package.scala 93:22:@7384.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_37 RetimeWrapper_6 ( // @[package.scala 93:22:@7417.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_37 RetimeWrapper_7 ( // @[package.scala 93:22:@7450.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_37 RetimeWrapper_8 ( // @[package.scala 93:22:@7483.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_37 RetimeWrapper_9 ( // @[package.scala 93:22:@7516.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_37 RetimeWrapper_10 ( // @[package.scala 93:22:@7549.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_37 RetimeWrapper_11 ( // @[package.scala 93:22:@7582.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_37 RetimeWrapper_12 ( // @[package.scala 93:22:@7615.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_37 RetimeWrapper_13 ( // @[package.scala 93:22:@7648.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_37 RetimeWrapper_14 ( // @[package.scala 93:22:@7681.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_37 RetimeWrapper_15 ( // @[package.scala 93:22:@7714.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  assign _T_1357 = ~ io_sigsIn_break; // @[sm_x343_inr_UnitPipe.scala 140:124:@7201.4]
  assign _T_1361 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 55:10:@7204.4]
  assign _T_1366 = io_in_x273_a_0_rPort_9_output_0[31]; // @[FixedPoint.scala 50:25:@7214.4]
  assign _T_1370 = _T_1366 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12:@7216.4]
  assign _T_1400 = io_in_x273_a_0_rPort_7_output_0[31]; // @[FixedPoint.scala 50:25:@7247.4]
  assign _T_1404 = _T_1400 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12:@7249.4]
  assign _T_1434 = io_in_x273_a_0_rPort_1_output_0[31]; // @[FixedPoint.scala 50:25:@7280.4]
  assign _T_1438 = _T_1434 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12:@7282.4]
  assign _T_1468 = io_in_x273_a_0_rPort_13_output_0[31]; // @[FixedPoint.scala 50:25:@7313.4]
  assign _T_1472 = _T_1468 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12:@7315.4]
  assign _T_1502 = io_in_x273_a_0_rPort_4_output_0[31]; // @[FixedPoint.scala 50:25:@7346.4]
  assign _T_1506 = _T_1502 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12:@7348.4]
  assign _T_1536 = io_in_x273_a_0_rPort_10_output_0[31]; // @[FixedPoint.scala 50:25:@7379.4]
  assign _T_1540 = _T_1536 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12:@7381.4]
  assign _T_1570 = io_in_x273_a_0_rPort_8_output_0[31]; // @[FixedPoint.scala 50:25:@7412.4]
  assign _T_1574 = _T_1570 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12:@7414.4]
  assign _T_1604 = io_in_x273_a_0_rPort_3_output_0[31]; // @[FixedPoint.scala 50:25:@7445.4]
  assign _T_1608 = _T_1604 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12:@7447.4]
  assign _T_1638 = io_in_x273_a_0_rPort_12_output_0[31]; // @[FixedPoint.scala 50:25:@7478.4]
  assign _T_1642 = _T_1638 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12:@7480.4]
  assign _T_1672 = io_in_x273_a_0_rPort_14_output_0[31]; // @[FixedPoint.scala 50:25:@7511.4]
  assign _T_1676 = _T_1672 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12:@7513.4]
  assign _T_1706 = io_in_x273_a_0_rPort_2_output_0[31]; // @[FixedPoint.scala 50:25:@7544.4]
  assign _T_1710 = _T_1706 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12:@7546.4]
  assign _T_1740 = io_in_x273_a_0_rPort_6_output_0[31]; // @[FixedPoint.scala 50:25:@7577.4]
  assign _T_1744 = _T_1740 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12:@7579.4]
  assign _T_1774 = io_in_x273_a_0_rPort_11_output_0[31]; // @[FixedPoint.scala 50:25:@7610.4]
  assign _T_1778 = _T_1774 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12:@7612.4]
  assign _T_1808 = io_in_x273_a_0_rPort_5_output_0[31]; // @[FixedPoint.scala 50:25:@7643.4]
  assign _T_1812 = _T_1808 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12:@7645.4]
  assign _T_1842 = io_in_x273_a_0_rPort_15_output_0[31]; // @[FixedPoint.scala 50:25:@7676.4]
  assign _T_1846 = _T_1842 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12:@7678.4]
  assign _T_1876 = io_in_x273_a_0_rPort_0_output_0[31]; // @[FixedPoint.scala 50:25:@7709.4]
  assign _T_1880 = _T_1876 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12:@7711.4]
  assign io_in_x269_argOut_port_0_valid = RetimeWrapper_14_io_out; // @[MemInterfaceType.scala 311:132:@7690.4]
  assign io_in_x269_argOut_port_0_bits = {_T_1846,io_in_x273_a_0_rPort_15_output_0}; // @[MemInterfaceType.scala 311:109:@7689.4]
  assign io_in_x257_argOut_port_0_valid = RetimeWrapper_2_io_out; // @[MemInterfaceType.scala 311:132:@7294.4]
  assign io_in_x257_argOut_port_0_bits = {_T_1438,io_in_x273_a_0_rPort_1_output_0}; // @[MemInterfaceType.scala 311:109:@7293.4]
  assign io_in_x261_argOut_port_0_valid = RetimeWrapper_6_io_out; // @[MemInterfaceType.scala 311:132:@7426.4]
  assign io_in_x261_argOut_port_0_bits = {_T_1574,io_in_x273_a_0_rPort_8_output_0}; // @[MemInterfaceType.scala 311:109:@7425.4]
  assign io_in_x265_argOut_port_0_valid = RetimeWrapper_10_io_out; // @[MemInterfaceType.scala 311:132:@7558.4]
  assign io_in_x265_argOut_port_0_bits = {_T_1710,io_in_x273_a_0_rPort_2_output_0}; // @[MemInterfaceType.scala 311:109:@7557.4]
  assign io_in_x270_argOut_port_0_valid = RetimeWrapper_15_io_out; // @[MemInterfaceType.scala 311:132:@7723.4]
  assign io_in_x270_argOut_port_0_bits = {_T_1880,io_in_x273_a_0_rPort_0_output_0}; // @[MemInterfaceType.scala 311:109:@7722.4]
  assign io_in_x260_argOut_port_0_valid = RetimeWrapper_5_io_out; // @[MemInterfaceType.scala 311:132:@7393.4]
  assign io_in_x260_argOut_port_0_bits = {_T_1540,io_in_x273_a_0_rPort_10_output_0}; // @[MemInterfaceType.scala 311:109:@7392.4]
  assign io_in_x256_argOut_port_0_valid = RetimeWrapper_1_io_out; // @[MemInterfaceType.scala 311:132:@7261.4]
  assign io_in_x256_argOut_port_0_bits = {_T_1404,io_in_x273_a_0_rPort_7_output_0}; // @[MemInterfaceType.scala 311:109:@7260.4]
  assign io_in_x266_argOut_port_0_valid = RetimeWrapper_11_io_out; // @[MemInterfaceType.scala 311:132:@7591.4]
  assign io_in_x266_argOut_port_0_bits = {_T_1744,io_in_x273_a_0_rPort_6_output_0}; // @[MemInterfaceType.scala 311:109:@7590.4]
  assign io_in_x264_argOut_port_0_valid = RetimeWrapper_9_io_out; // @[MemInterfaceType.scala 311:132:@7525.4]
  assign io_in_x264_argOut_port_0_bits = {_T_1676,io_in_x273_a_0_rPort_14_output_0}; // @[MemInterfaceType.scala 311:109:@7524.4]
  assign io_in_x259_argOut_port_0_valid = RetimeWrapper_4_io_out; // @[MemInterfaceType.scala 311:132:@7360.4]
  assign io_in_x259_argOut_port_0_bits = {_T_1506,io_in_x273_a_0_rPort_4_output_0}; // @[MemInterfaceType.scala 311:109:@7359.4]
  assign io_in_x267_argOut_port_0_valid = RetimeWrapper_12_io_out; // @[MemInterfaceType.scala 311:132:@7624.4]
  assign io_in_x267_argOut_port_0_bits = {_T_1778,io_in_x273_a_0_rPort_11_output_0}; // @[MemInterfaceType.scala 311:109:@7623.4]
  assign io_in_x255_argOut_port_0_valid = RetimeWrapper_io_out; // @[MemInterfaceType.scala 311:132:@7228.4]
  assign io_in_x255_argOut_port_0_bits = {_T_1370,io_in_x273_a_0_rPort_9_output_0}; // @[MemInterfaceType.scala 311:109:@7227.4]
  assign io_in_x263_argOut_port_0_valid = RetimeWrapper_8_io_out; // @[MemInterfaceType.scala 311:132:@7492.4]
  assign io_in_x263_argOut_port_0_bits = {_T_1642,io_in_x273_a_0_rPort_12_output_0}; // @[MemInterfaceType.scala 311:109:@7491.4]
  assign io_in_x258_argOut_port_0_valid = RetimeWrapper_3_io_out; // @[MemInterfaceType.scala 311:132:@7327.4]
  assign io_in_x258_argOut_port_0_bits = {_T_1472,io_in_x273_a_0_rPort_13_output_0}; // @[MemInterfaceType.scala 311:109:@7326.4]
  assign io_in_x262_argOut_port_0_valid = RetimeWrapper_7_io_out; // @[MemInterfaceType.scala 311:132:@7459.4]
  assign io_in_x262_argOut_port_0_bits = {_T_1608,io_in_x273_a_0_rPort_3_output_0}; // @[MemInterfaceType.scala 311:109:@7458.4]
  assign io_in_x273_a_0_rPort_15_en_0 = _T_1357 & _T_1361; // @[MemInterfaceType.scala 110:79:@7672.4]
  assign io_in_x273_a_0_rPort_14_en_0 = _T_1357 & _T_1361; // @[MemInterfaceType.scala 110:79:@7507.4]
  assign io_in_x273_a_0_rPort_13_en_0 = _T_1357 & _T_1361; // @[MemInterfaceType.scala 110:79:@7309.4]
  assign io_in_x273_a_0_rPort_12_en_0 = _T_1357 & _T_1361; // @[MemInterfaceType.scala 110:79:@7474.4]
  assign io_in_x273_a_0_rPort_11_en_0 = _T_1357 & _T_1361; // @[MemInterfaceType.scala 110:79:@7606.4]
  assign io_in_x273_a_0_rPort_10_en_0 = _T_1357 & _T_1361; // @[MemInterfaceType.scala 110:79:@7375.4]
  assign io_in_x273_a_0_rPort_9_en_0 = _T_1357 & _T_1361; // @[MemInterfaceType.scala 110:79:@7210.4]
  assign io_in_x273_a_0_rPort_8_en_0 = _T_1357 & _T_1361; // @[MemInterfaceType.scala 110:79:@7408.4]
  assign io_in_x273_a_0_rPort_7_en_0 = _T_1357 & _T_1361; // @[MemInterfaceType.scala 110:79:@7243.4]
  assign io_in_x273_a_0_rPort_6_en_0 = _T_1357 & _T_1361; // @[MemInterfaceType.scala 110:79:@7573.4]
  assign io_in_x273_a_0_rPort_5_en_0 = _T_1357 & _T_1361; // @[MemInterfaceType.scala 110:79:@7639.4]
  assign io_in_x273_a_0_rPort_4_en_0 = _T_1357 & _T_1361; // @[MemInterfaceType.scala 110:79:@7342.4]
  assign io_in_x273_a_0_rPort_3_en_0 = _T_1357 & _T_1361; // @[MemInterfaceType.scala 110:79:@7441.4]
  assign io_in_x273_a_0_rPort_2_en_0 = _T_1357 & _T_1361; // @[MemInterfaceType.scala 110:79:@7540.4]
  assign io_in_x273_a_0_rPort_1_en_0 = _T_1357 & _T_1361; // @[MemInterfaceType.scala 110:79:@7276.4]
  assign io_in_x273_a_0_rPort_0_en_0 = _T_1357 & _T_1361; // @[MemInterfaceType.scala 110:79:@7705.4]
  assign io_in_x268_argOut_port_0_valid = RetimeWrapper_13_io_out; // @[MemInterfaceType.scala 311:132:@7657.4]
  assign io_in_x268_argOut_port_0_bits = {_T_1812,io_in_x273_a_0_rPort_5_output_0}; // @[MemInterfaceType.scala 311:109:@7656.4]
  assign RetimeWrapper_clock = clock; // @[:@7220.4]
  assign RetimeWrapper_reset = reset; // @[:@7221.4]
  assign RetimeWrapper_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@7222.4]
  assign RetimeWrapper_1_clock = clock; // @[:@7253.4]
  assign RetimeWrapper_1_reset = reset; // @[:@7254.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@7255.4]
  assign RetimeWrapper_2_clock = clock; // @[:@7286.4]
  assign RetimeWrapper_2_reset = reset; // @[:@7287.4]
  assign RetimeWrapper_2_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@7288.4]
  assign RetimeWrapper_3_clock = clock; // @[:@7319.4]
  assign RetimeWrapper_3_reset = reset; // @[:@7320.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@7321.4]
  assign RetimeWrapper_4_clock = clock; // @[:@7352.4]
  assign RetimeWrapper_4_reset = reset; // @[:@7353.4]
  assign RetimeWrapper_4_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@7354.4]
  assign RetimeWrapper_5_clock = clock; // @[:@7385.4]
  assign RetimeWrapper_5_reset = reset; // @[:@7386.4]
  assign RetimeWrapper_5_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@7387.4]
  assign RetimeWrapper_6_clock = clock; // @[:@7418.4]
  assign RetimeWrapper_6_reset = reset; // @[:@7419.4]
  assign RetimeWrapper_6_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@7420.4]
  assign RetimeWrapper_7_clock = clock; // @[:@7451.4]
  assign RetimeWrapper_7_reset = reset; // @[:@7452.4]
  assign RetimeWrapper_7_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@7453.4]
  assign RetimeWrapper_8_clock = clock; // @[:@7484.4]
  assign RetimeWrapper_8_reset = reset; // @[:@7485.4]
  assign RetimeWrapper_8_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@7486.4]
  assign RetimeWrapper_9_clock = clock; // @[:@7517.4]
  assign RetimeWrapper_9_reset = reset; // @[:@7518.4]
  assign RetimeWrapper_9_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@7519.4]
  assign RetimeWrapper_10_clock = clock; // @[:@7550.4]
  assign RetimeWrapper_10_reset = reset; // @[:@7551.4]
  assign RetimeWrapper_10_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@7552.4]
  assign RetimeWrapper_11_clock = clock; // @[:@7583.4]
  assign RetimeWrapper_11_reset = reset; // @[:@7584.4]
  assign RetimeWrapper_11_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@7585.4]
  assign RetimeWrapper_12_clock = clock; // @[:@7616.4]
  assign RetimeWrapper_12_reset = reset; // @[:@7617.4]
  assign RetimeWrapper_12_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@7618.4]
  assign RetimeWrapper_13_clock = clock; // @[:@7649.4]
  assign RetimeWrapper_13_reset = reset; // @[:@7650.4]
  assign RetimeWrapper_13_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@7651.4]
  assign RetimeWrapper_14_clock = clock; // @[:@7682.4]
  assign RetimeWrapper_14_reset = reset; // @[:@7683.4]
  assign RetimeWrapper_14_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@7684.4]
  assign RetimeWrapper_15_clock = clock; // @[:@7715.4]
  assign RetimeWrapper_15_reset = reset; // @[:@7716.4]
  assign RetimeWrapper_15_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@7717.4]
endmodule
module RootController_kernelRootController_concrete1( // @[:@7725.2]
  input         clock, // @[:@7726.4]
  input         reset, // @[:@7727.4]
  output        io_in_x269_argOut_port_0_valid, // @[:@7728.4]
  output [63:0] io_in_x269_argOut_port_0_bits, // @[:@7728.4]
  output        io_in_x257_argOut_port_0_valid, // @[:@7728.4]
  output [63:0] io_in_x257_argOut_port_0_bits, // @[:@7728.4]
  output        io_in_x261_argOut_port_0_valid, // @[:@7728.4]
  output [63:0] io_in_x261_argOut_port_0_bits, // @[:@7728.4]
  output        io_in_x265_argOut_port_0_valid, // @[:@7728.4]
  output [63:0] io_in_x265_argOut_port_0_bits, // @[:@7728.4]
  output        io_in_x270_argOut_port_0_valid, // @[:@7728.4]
  output [63:0] io_in_x270_argOut_port_0_bits, // @[:@7728.4]
  output        io_in_x260_argOut_port_0_valid, // @[:@7728.4]
  output [63:0] io_in_x260_argOut_port_0_bits, // @[:@7728.4]
  output        io_in_x275_ready, // @[:@7728.4]
  input         io_in_x275_valid, // @[:@7728.4]
  input  [31:0] io_in_x275_bits_rdata_0, // @[:@7728.4]
  output        io_in_x256_argOut_port_0_valid, // @[:@7728.4]
  output [63:0] io_in_x256_argOut_port_0_bits, // @[:@7728.4]
  output        io_in_x266_argOut_port_0_valid, // @[:@7728.4]
  output [63:0] io_in_x266_argOut_port_0_bits, // @[:@7728.4]
  output        io_in_x264_argOut_port_0_valid, // @[:@7728.4]
  output [63:0] io_in_x264_argOut_port_0_bits, // @[:@7728.4]
  output        io_in_x259_argOut_port_0_valid, // @[:@7728.4]
  output [63:0] io_in_x259_argOut_port_0_bits, // @[:@7728.4]
  input         io_in_x274_ready, // @[:@7728.4]
  output        io_in_x274_valid, // @[:@7728.4]
  output [63:0] io_in_x274_bits_addr, // @[:@7728.4]
  output [31:0] io_in_x274_bits_size, // @[:@7728.4]
  output        io_in_x267_argOut_port_0_valid, // @[:@7728.4]
  output [63:0] io_in_x267_argOut_port_0_bits, // @[:@7728.4]
  output        io_in_x255_argOut_port_0_valid, // @[:@7728.4]
  output [63:0] io_in_x255_argOut_port_0_bits, // @[:@7728.4]
  output        io_in_x263_argOut_port_0_valid, // @[:@7728.4]
  output [63:0] io_in_x263_argOut_port_0_bits, // @[:@7728.4]
  output        io_in_x258_argOut_port_0_valid, // @[:@7728.4]
  output [63:0] io_in_x258_argOut_port_0_bits, // @[:@7728.4]
  output        io_in_x262_argOut_port_0_valid, // @[:@7728.4]
  output [63:0] io_in_x262_argOut_port_0_bits, // @[:@7728.4]
  output        io_in_x268_argOut_port_0_valid, // @[:@7728.4]
  output [63:0] io_in_x268_argOut_port_0_bits, // @[:@7728.4]
  input  [63:0] io_in_x254_in_number, // @[:@7728.4]
  input         io_sigsIn_smEnableOuts_0, // @[:@7728.4]
  input         io_sigsIn_smEnableOuts_1, // @[:@7728.4]
  input         io_sigsIn_smChildAcks_0, // @[:@7728.4]
  input         io_sigsIn_smChildAcks_1, // @[:@7728.4]
  output        io_sigsOut_smDoneIn_0, // @[:@7728.4]
  output        io_sigsOut_smDoneIn_1, // @[:@7728.4]
  input         io_rr // @[:@7728.4]
);
  wire  x273_a_0_clock; // @[m_x273_a_0.scala 41:17:@7804.4]
  wire  x273_a_0_reset; // @[m_x273_a_0.scala 41:17:@7804.4]
  wire  x273_a_0_io_rPort_15_en_0; // @[m_x273_a_0.scala 41:17:@7804.4]
  wire [31:0] x273_a_0_io_rPort_15_output_0; // @[m_x273_a_0.scala 41:17:@7804.4]
  wire  x273_a_0_io_rPort_14_en_0; // @[m_x273_a_0.scala 41:17:@7804.4]
  wire [31:0] x273_a_0_io_rPort_14_output_0; // @[m_x273_a_0.scala 41:17:@7804.4]
  wire  x273_a_0_io_rPort_13_en_0; // @[m_x273_a_0.scala 41:17:@7804.4]
  wire [31:0] x273_a_0_io_rPort_13_output_0; // @[m_x273_a_0.scala 41:17:@7804.4]
  wire  x273_a_0_io_rPort_12_en_0; // @[m_x273_a_0.scala 41:17:@7804.4]
  wire [31:0] x273_a_0_io_rPort_12_output_0; // @[m_x273_a_0.scala 41:17:@7804.4]
  wire  x273_a_0_io_rPort_11_en_0; // @[m_x273_a_0.scala 41:17:@7804.4]
  wire [31:0] x273_a_0_io_rPort_11_output_0; // @[m_x273_a_0.scala 41:17:@7804.4]
  wire  x273_a_0_io_rPort_10_en_0; // @[m_x273_a_0.scala 41:17:@7804.4]
  wire [31:0] x273_a_0_io_rPort_10_output_0; // @[m_x273_a_0.scala 41:17:@7804.4]
  wire  x273_a_0_io_rPort_9_en_0; // @[m_x273_a_0.scala 41:17:@7804.4]
  wire [31:0] x273_a_0_io_rPort_9_output_0; // @[m_x273_a_0.scala 41:17:@7804.4]
  wire  x273_a_0_io_rPort_8_en_0; // @[m_x273_a_0.scala 41:17:@7804.4]
  wire [31:0] x273_a_0_io_rPort_8_output_0; // @[m_x273_a_0.scala 41:17:@7804.4]
  wire  x273_a_0_io_rPort_7_en_0; // @[m_x273_a_0.scala 41:17:@7804.4]
  wire [31:0] x273_a_0_io_rPort_7_output_0; // @[m_x273_a_0.scala 41:17:@7804.4]
  wire  x273_a_0_io_rPort_6_en_0; // @[m_x273_a_0.scala 41:17:@7804.4]
  wire [31:0] x273_a_0_io_rPort_6_output_0; // @[m_x273_a_0.scala 41:17:@7804.4]
  wire  x273_a_0_io_rPort_5_en_0; // @[m_x273_a_0.scala 41:17:@7804.4]
  wire [31:0] x273_a_0_io_rPort_5_output_0; // @[m_x273_a_0.scala 41:17:@7804.4]
  wire  x273_a_0_io_rPort_4_en_0; // @[m_x273_a_0.scala 41:17:@7804.4]
  wire [31:0] x273_a_0_io_rPort_4_output_0; // @[m_x273_a_0.scala 41:17:@7804.4]
  wire  x273_a_0_io_rPort_3_en_0; // @[m_x273_a_0.scala 41:17:@7804.4]
  wire [31:0] x273_a_0_io_rPort_3_output_0; // @[m_x273_a_0.scala 41:17:@7804.4]
  wire  x273_a_0_io_rPort_2_en_0; // @[m_x273_a_0.scala 41:17:@7804.4]
  wire [31:0] x273_a_0_io_rPort_2_output_0; // @[m_x273_a_0.scala 41:17:@7804.4]
  wire  x273_a_0_io_rPort_1_en_0; // @[m_x273_a_0.scala 41:17:@7804.4]
  wire [31:0] x273_a_0_io_rPort_1_output_0; // @[m_x273_a_0.scala 41:17:@7804.4]
  wire  x273_a_0_io_rPort_0_en_0; // @[m_x273_a_0.scala 41:17:@7804.4]
  wire [31:0] x273_a_0_io_rPort_0_output_0; // @[m_x273_a_0.scala 41:17:@7804.4]
  wire [4:0] x273_a_0_io_wPort_0_banks_0; // @[m_x273_a_0.scala 41:17:@7804.4]
  wire  x273_a_0_io_wPort_0_ofs_0; // @[m_x273_a_0.scala 41:17:@7804.4]
  wire [31:0] x273_a_0_io_wPort_0_data_0; // @[m_x273_a_0.scala 41:17:@7804.4]
  wire  x273_a_0_io_wPort_0_en_0; // @[m_x273_a_0.scala 41:17:@7804.4]
  wire  x294_outr_UnitPipe_sm_clock; // @[sm_x294_outr_UnitPipe.scala 34:18:@7943.4]
  wire  x294_outr_UnitPipe_sm_reset; // @[sm_x294_outr_UnitPipe.scala 34:18:@7943.4]
  wire  x294_outr_UnitPipe_sm_io_enable; // @[sm_x294_outr_UnitPipe.scala 34:18:@7943.4]
  wire  x294_outr_UnitPipe_sm_io_done; // @[sm_x294_outr_UnitPipe.scala 34:18:@7943.4]
  wire  x294_outr_UnitPipe_sm_io_parentAck; // @[sm_x294_outr_UnitPipe.scala 34:18:@7943.4]
  wire  x294_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x294_outr_UnitPipe.scala 34:18:@7943.4]
  wire  x294_outr_UnitPipe_sm_io_doneIn_1; // @[sm_x294_outr_UnitPipe.scala 34:18:@7943.4]
  wire  x294_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x294_outr_UnitPipe.scala 34:18:@7943.4]
  wire  x294_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x294_outr_UnitPipe.scala 34:18:@7943.4]
  wire  x294_outr_UnitPipe_sm_io_childAck_0; // @[sm_x294_outr_UnitPipe.scala 34:18:@7943.4]
  wire  x294_outr_UnitPipe_sm_io_childAck_1; // @[sm_x294_outr_UnitPipe.scala 34:18:@7943.4]
  wire  x294_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x294_outr_UnitPipe.scala 34:18:@7943.4]
  wire  x294_outr_UnitPipe_sm_io_ctrCopyDone_1; // @[sm_x294_outr_UnitPipe.scala 34:18:@7943.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@8005.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@8005.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@8005.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@8005.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@8005.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@8013.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@8013.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@8013.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@8013.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@8013.4]
  wire  x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_clock; // @[sm_x294_outr_UnitPipe.scala 93:24:@8041.4]
  wire  x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_reset; // @[sm_x294_outr_UnitPipe.scala 93:24:@8041.4]
  wire [4:0] x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_in_x273_a_0_wPort_0_banks_0; // @[sm_x294_outr_UnitPipe.scala 93:24:@8041.4]
  wire  x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_in_x273_a_0_wPort_0_ofs_0; // @[sm_x294_outr_UnitPipe.scala 93:24:@8041.4]
  wire [31:0] x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_in_x273_a_0_wPort_0_data_0; // @[sm_x294_outr_UnitPipe.scala 93:24:@8041.4]
  wire  x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_in_x273_a_0_wPort_0_en_0; // @[sm_x294_outr_UnitPipe.scala 93:24:@8041.4]
  wire [63:0] x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_in_x254_in_number; // @[sm_x294_outr_UnitPipe.scala 93:24:@8041.4]
  wire  x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_in_x274_ready; // @[sm_x294_outr_UnitPipe.scala 93:24:@8041.4]
  wire  x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_in_x274_valid; // @[sm_x294_outr_UnitPipe.scala 93:24:@8041.4]
  wire [63:0] x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_in_x274_bits_addr; // @[sm_x294_outr_UnitPipe.scala 93:24:@8041.4]
  wire [31:0] x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_in_x274_bits_size; // @[sm_x294_outr_UnitPipe.scala 93:24:@8041.4]
  wire  x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_in_x275_ready; // @[sm_x294_outr_UnitPipe.scala 93:24:@8041.4]
  wire  x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_in_x275_valid; // @[sm_x294_outr_UnitPipe.scala 93:24:@8041.4]
  wire [31:0] x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_in_x275_bits_rdata_0; // @[sm_x294_outr_UnitPipe.scala 93:24:@8041.4]
  wire  x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x294_outr_UnitPipe.scala 93:24:@8041.4]
  wire  x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x294_outr_UnitPipe.scala 93:24:@8041.4]
  wire  x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x294_outr_UnitPipe.scala 93:24:@8041.4]
  wire  x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x294_outr_UnitPipe.scala 93:24:@8041.4]
  wire  x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x294_outr_UnitPipe.scala 93:24:@8041.4]
  wire  x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x294_outr_UnitPipe.scala 93:24:@8041.4]
  wire  x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x294_outr_UnitPipe.scala 93:24:@8041.4]
  wire  x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[sm_x294_outr_UnitPipe.scala 93:24:@8041.4]
  wire  x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_rr; // @[sm_x294_outr_UnitPipe.scala 93:24:@8041.4]
  wire  x343_inr_UnitPipe_sm_clock; // @[sm_x343_inr_UnitPipe.scala 32:18:@8267.4]
  wire  x343_inr_UnitPipe_sm_reset; // @[sm_x343_inr_UnitPipe.scala 32:18:@8267.4]
  wire  x343_inr_UnitPipe_sm_io_enable; // @[sm_x343_inr_UnitPipe.scala 32:18:@8267.4]
  wire  x343_inr_UnitPipe_sm_io_done; // @[sm_x343_inr_UnitPipe.scala 32:18:@8267.4]
  wire  x343_inr_UnitPipe_sm_io_ctrDone; // @[sm_x343_inr_UnitPipe.scala 32:18:@8267.4]
  wire  x343_inr_UnitPipe_sm_io_datapathEn; // @[sm_x343_inr_UnitPipe.scala 32:18:@8267.4]
  wire  x343_inr_UnitPipe_sm_io_ctrInc; // @[sm_x343_inr_UnitPipe.scala 32:18:@8267.4]
  wire  x343_inr_UnitPipe_sm_io_parentAck; // @[sm_x343_inr_UnitPipe.scala 32:18:@8267.4]
  wire  x343_inr_UnitPipe_sm_io_break; // @[sm_x343_inr_UnitPipe.scala 32:18:@8267.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@8324.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@8324.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@8324.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@8324.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@8324.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@8332.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@8332.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@8332.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@8332.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@8332.4]
  wire  x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_clock; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire  x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_reset; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire  x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x269_argOut_port_0_valid; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire [63:0] x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x269_argOut_port_0_bits; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire  x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x257_argOut_port_0_valid; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire [63:0] x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x257_argOut_port_0_bits; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire  x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x261_argOut_port_0_valid; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire [63:0] x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x261_argOut_port_0_bits; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire  x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x265_argOut_port_0_valid; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire [63:0] x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x265_argOut_port_0_bits; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire  x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x270_argOut_port_0_valid; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire [63:0] x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x270_argOut_port_0_bits; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire  x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x260_argOut_port_0_valid; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire [63:0] x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x260_argOut_port_0_bits; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire  x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x256_argOut_port_0_valid; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire [63:0] x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x256_argOut_port_0_bits; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire  x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x266_argOut_port_0_valid; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire [63:0] x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x266_argOut_port_0_bits; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire  x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x264_argOut_port_0_valid; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire [63:0] x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x264_argOut_port_0_bits; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire  x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x259_argOut_port_0_valid; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire [63:0] x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x259_argOut_port_0_bits; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire  x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x267_argOut_port_0_valid; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire [63:0] x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x267_argOut_port_0_bits; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire  x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x255_argOut_port_0_valid; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire [63:0] x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x255_argOut_port_0_bits; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire  x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x263_argOut_port_0_valid; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire [63:0] x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x263_argOut_port_0_bits; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire  x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x258_argOut_port_0_valid; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire [63:0] x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x258_argOut_port_0_bits; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire  x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x262_argOut_port_0_valid; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire [63:0] x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x262_argOut_port_0_bits; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire  x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_15_en_0; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire [31:0] x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_15_output_0; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire  x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_14_en_0; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire [31:0] x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_14_output_0; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire  x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_13_en_0; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire [31:0] x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_13_output_0; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire  x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_12_en_0; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire [31:0] x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_12_output_0; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire  x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_11_en_0; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire [31:0] x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_11_output_0; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire  x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_10_en_0; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire [31:0] x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_10_output_0; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire  x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_9_en_0; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire [31:0] x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_9_output_0; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire  x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_8_en_0; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire [31:0] x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_8_output_0; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire  x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_7_en_0; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire [31:0] x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_7_output_0; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire  x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_6_en_0; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire [31:0] x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_6_output_0; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire  x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_5_en_0; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire [31:0] x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_5_output_0; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire  x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_4_en_0; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire [31:0] x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_4_output_0; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire  x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_3_en_0; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire [31:0] x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_3_output_0; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire  x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_2_en_0; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire [31:0] x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_2_output_0; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire  x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_1_en_0; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire [31:0] x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_1_output_0; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire  x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_0_en_0; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire [31:0] x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_0_output_0; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire  x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x268_argOut_port_0_valid; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire [63:0] x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x268_argOut_port_0_bits; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire  x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_sigsIn_datapathEn; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire  x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_sigsIn_break; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire  x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_rr; // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
  wire  _T_545; // @[package.scala 96:25:@8010.4 package.scala 96:25:@8011.4]
  wire  _T_551; // @[package.scala 96:25:@8018.4 package.scala 96:25:@8019.4]
  wire  _T_554; // @[SpatialBlocks.scala 110:93:@8021.4]
  wire  _T_620; // @[package.scala 100:49:@8295.4]
  reg  _T_623; // @[package.scala 48:56:@8296.4]
  reg [31:0] _RAND_0;
  wire  _T_637; // @[package.scala 96:25:@8329.4 package.scala 96:25:@8330.4]
  wire  _T_643; // @[package.scala 96:25:@8337.4 package.scala 96:25:@8338.4]
  wire  _T_646; // @[SpatialBlocks.scala 110:93:@8340.4]
  x273_a_0 x273_a_0 ( // @[m_x273_a_0.scala 41:17:@7804.4]
    .clock(x273_a_0_clock),
    .reset(x273_a_0_reset),
    .io_rPort_15_en_0(x273_a_0_io_rPort_15_en_0),
    .io_rPort_15_output_0(x273_a_0_io_rPort_15_output_0),
    .io_rPort_14_en_0(x273_a_0_io_rPort_14_en_0),
    .io_rPort_14_output_0(x273_a_0_io_rPort_14_output_0),
    .io_rPort_13_en_0(x273_a_0_io_rPort_13_en_0),
    .io_rPort_13_output_0(x273_a_0_io_rPort_13_output_0),
    .io_rPort_12_en_0(x273_a_0_io_rPort_12_en_0),
    .io_rPort_12_output_0(x273_a_0_io_rPort_12_output_0),
    .io_rPort_11_en_0(x273_a_0_io_rPort_11_en_0),
    .io_rPort_11_output_0(x273_a_0_io_rPort_11_output_0),
    .io_rPort_10_en_0(x273_a_0_io_rPort_10_en_0),
    .io_rPort_10_output_0(x273_a_0_io_rPort_10_output_0),
    .io_rPort_9_en_0(x273_a_0_io_rPort_9_en_0),
    .io_rPort_9_output_0(x273_a_0_io_rPort_9_output_0),
    .io_rPort_8_en_0(x273_a_0_io_rPort_8_en_0),
    .io_rPort_8_output_0(x273_a_0_io_rPort_8_output_0),
    .io_rPort_7_en_0(x273_a_0_io_rPort_7_en_0),
    .io_rPort_7_output_0(x273_a_0_io_rPort_7_output_0),
    .io_rPort_6_en_0(x273_a_0_io_rPort_6_en_0),
    .io_rPort_6_output_0(x273_a_0_io_rPort_6_output_0),
    .io_rPort_5_en_0(x273_a_0_io_rPort_5_en_0),
    .io_rPort_5_output_0(x273_a_0_io_rPort_5_output_0),
    .io_rPort_4_en_0(x273_a_0_io_rPort_4_en_0),
    .io_rPort_4_output_0(x273_a_0_io_rPort_4_output_0),
    .io_rPort_3_en_0(x273_a_0_io_rPort_3_en_0),
    .io_rPort_3_output_0(x273_a_0_io_rPort_3_output_0),
    .io_rPort_2_en_0(x273_a_0_io_rPort_2_en_0),
    .io_rPort_2_output_0(x273_a_0_io_rPort_2_output_0),
    .io_rPort_1_en_0(x273_a_0_io_rPort_1_en_0),
    .io_rPort_1_output_0(x273_a_0_io_rPort_1_output_0),
    .io_rPort_0_en_0(x273_a_0_io_rPort_0_en_0),
    .io_rPort_0_output_0(x273_a_0_io_rPort_0_output_0),
    .io_wPort_0_banks_0(x273_a_0_io_wPort_0_banks_0),
    .io_wPort_0_ofs_0(x273_a_0_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x273_a_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x273_a_0_io_wPort_0_en_0)
  );
  x294_outr_UnitPipe_sm x294_outr_UnitPipe_sm ( // @[sm_x294_outr_UnitPipe.scala 34:18:@7943.4]
    .clock(x294_outr_UnitPipe_sm_clock),
    .reset(x294_outr_UnitPipe_sm_reset),
    .io_enable(x294_outr_UnitPipe_sm_io_enable),
    .io_done(x294_outr_UnitPipe_sm_io_done),
    .io_parentAck(x294_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x294_outr_UnitPipe_sm_io_doneIn_0),
    .io_doneIn_1(x294_outr_UnitPipe_sm_io_doneIn_1),
    .io_enableOut_0(x294_outr_UnitPipe_sm_io_enableOut_0),
    .io_enableOut_1(x294_outr_UnitPipe_sm_io_enableOut_1),
    .io_childAck_0(x294_outr_UnitPipe_sm_io_childAck_0),
    .io_childAck_1(x294_outr_UnitPipe_sm_io_childAck_1),
    .io_ctrCopyDone_0(x294_outr_UnitPipe_sm_io_ctrCopyDone_0),
    .io_ctrCopyDone_1(x294_outr_UnitPipe_sm_io_ctrCopyDone_1)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@8005.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@8013.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1 x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1 ( // @[sm_x294_outr_UnitPipe.scala 93:24:@8041.4]
    .clock(x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_clock),
    .reset(x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_reset),
    .io_in_x273_a_0_wPort_0_banks_0(x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_in_x273_a_0_wPort_0_banks_0),
    .io_in_x273_a_0_wPort_0_ofs_0(x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_in_x273_a_0_wPort_0_ofs_0),
    .io_in_x273_a_0_wPort_0_data_0(x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_in_x273_a_0_wPort_0_data_0),
    .io_in_x273_a_0_wPort_0_en_0(x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_in_x273_a_0_wPort_0_en_0),
    .io_in_x254_in_number(x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_in_x254_in_number),
    .io_in_x274_ready(x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_in_x274_ready),
    .io_in_x274_valid(x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_in_x274_valid),
    .io_in_x274_bits_addr(x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_in_x274_bits_addr),
    .io_in_x274_bits_size(x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_in_x274_bits_size),
    .io_in_x275_ready(x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_in_x275_ready),
    .io_in_x275_valid(x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_in_x275_valid),
    .io_in_x275_bits_rdata_0(x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_in_x275_bits_rdata_0),
    .io_sigsIn_smEnableOuts_0(x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smChildAcks_0(x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsOut_smDoneIn_0(x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1),
    .io_sigsOut_smCtrCopyDone_0(x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_sigsOut_smCtrCopyDone_1(x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1),
    .io_rr(x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_rr)
  );
  x343_inr_UnitPipe_sm x343_inr_UnitPipe_sm ( // @[sm_x343_inr_UnitPipe.scala 32:18:@8267.4]
    .clock(x343_inr_UnitPipe_sm_clock),
    .reset(x343_inr_UnitPipe_sm_reset),
    .io_enable(x343_inr_UnitPipe_sm_io_enable),
    .io_done(x343_inr_UnitPipe_sm_io_done),
    .io_ctrDone(x343_inr_UnitPipe_sm_io_ctrDone),
    .io_datapathEn(x343_inr_UnitPipe_sm_io_datapathEn),
    .io_ctrInc(x343_inr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x343_inr_UnitPipe_sm_io_parentAck),
    .io_break(x343_inr_UnitPipe_sm_io_break)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@8324.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@8332.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1 x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1 ( // @[sm_x343_inr_UnitPipe.scala 265:24:@8358.4]
    .clock(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_clock),
    .reset(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_reset),
    .io_in_x269_argOut_port_0_valid(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x269_argOut_port_0_valid),
    .io_in_x269_argOut_port_0_bits(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x269_argOut_port_0_bits),
    .io_in_x257_argOut_port_0_valid(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x257_argOut_port_0_valid),
    .io_in_x257_argOut_port_0_bits(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x257_argOut_port_0_bits),
    .io_in_x261_argOut_port_0_valid(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x261_argOut_port_0_valid),
    .io_in_x261_argOut_port_0_bits(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x261_argOut_port_0_bits),
    .io_in_x265_argOut_port_0_valid(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x265_argOut_port_0_valid),
    .io_in_x265_argOut_port_0_bits(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x265_argOut_port_0_bits),
    .io_in_x270_argOut_port_0_valid(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x270_argOut_port_0_valid),
    .io_in_x270_argOut_port_0_bits(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x270_argOut_port_0_bits),
    .io_in_x260_argOut_port_0_valid(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x260_argOut_port_0_valid),
    .io_in_x260_argOut_port_0_bits(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x260_argOut_port_0_bits),
    .io_in_x256_argOut_port_0_valid(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x256_argOut_port_0_valid),
    .io_in_x256_argOut_port_0_bits(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x256_argOut_port_0_bits),
    .io_in_x266_argOut_port_0_valid(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x266_argOut_port_0_valid),
    .io_in_x266_argOut_port_0_bits(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x266_argOut_port_0_bits),
    .io_in_x264_argOut_port_0_valid(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x264_argOut_port_0_valid),
    .io_in_x264_argOut_port_0_bits(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x264_argOut_port_0_bits),
    .io_in_x259_argOut_port_0_valid(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x259_argOut_port_0_valid),
    .io_in_x259_argOut_port_0_bits(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x259_argOut_port_0_bits),
    .io_in_x267_argOut_port_0_valid(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x267_argOut_port_0_valid),
    .io_in_x267_argOut_port_0_bits(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x267_argOut_port_0_bits),
    .io_in_x255_argOut_port_0_valid(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x255_argOut_port_0_valid),
    .io_in_x255_argOut_port_0_bits(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x255_argOut_port_0_bits),
    .io_in_x263_argOut_port_0_valid(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x263_argOut_port_0_valid),
    .io_in_x263_argOut_port_0_bits(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x263_argOut_port_0_bits),
    .io_in_x258_argOut_port_0_valid(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x258_argOut_port_0_valid),
    .io_in_x258_argOut_port_0_bits(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x258_argOut_port_0_bits),
    .io_in_x262_argOut_port_0_valid(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x262_argOut_port_0_valid),
    .io_in_x262_argOut_port_0_bits(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x262_argOut_port_0_bits),
    .io_in_x273_a_0_rPort_15_en_0(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_15_en_0),
    .io_in_x273_a_0_rPort_15_output_0(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_15_output_0),
    .io_in_x273_a_0_rPort_14_en_0(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_14_en_0),
    .io_in_x273_a_0_rPort_14_output_0(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_14_output_0),
    .io_in_x273_a_0_rPort_13_en_0(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_13_en_0),
    .io_in_x273_a_0_rPort_13_output_0(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_13_output_0),
    .io_in_x273_a_0_rPort_12_en_0(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_12_en_0),
    .io_in_x273_a_0_rPort_12_output_0(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_12_output_0),
    .io_in_x273_a_0_rPort_11_en_0(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_11_en_0),
    .io_in_x273_a_0_rPort_11_output_0(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_11_output_0),
    .io_in_x273_a_0_rPort_10_en_0(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_10_en_0),
    .io_in_x273_a_0_rPort_10_output_0(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_10_output_0),
    .io_in_x273_a_0_rPort_9_en_0(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_9_en_0),
    .io_in_x273_a_0_rPort_9_output_0(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_9_output_0),
    .io_in_x273_a_0_rPort_8_en_0(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_8_en_0),
    .io_in_x273_a_0_rPort_8_output_0(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_8_output_0),
    .io_in_x273_a_0_rPort_7_en_0(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_7_en_0),
    .io_in_x273_a_0_rPort_7_output_0(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_7_output_0),
    .io_in_x273_a_0_rPort_6_en_0(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_6_en_0),
    .io_in_x273_a_0_rPort_6_output_0(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_6_output_0),
    .io_in_x273_a_0_rPort_5_en_0(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_5_en_0),
    .io_in_x273_a_0_rPort_5_output_0(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_5_output_0),
    .io_in_x273_a_0_rPort_4_en_0(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_4_en_0),
    .io_in_x273_a_0_rPort_4_output_0(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_4_output_0),
    .io_in_x273_a_0_rPort_3_en_0(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_3_en_0),
    .io_in_x273_a_0_rPort_3_output_0(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_3_output_0),
    .io_in_x273_a_0_rPort_2_en_0(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_2_en_0),
    .io_in_x273_a_0_rPort_2_output_0(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_2_output_0),
    .io_in_x273_a_0_rPort_1_en_0(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_1_en_0),
    .io_in_x273_a_0_rPort_1_output_0(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_1_output_0),
    .io_in_x273_a_0_rPort_0_en_0(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_0_en_0),
    .io_in_x273_a_0_rPort_0_output_0(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_0_output_0),
    .io_in_x268_argOut_port_0_valid(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x268_argOut_port_0_valid),
    .io_in_x268_argOut_port_0_bits(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x268_argOut_port_0_bits),
    .io_sigsIn_datapathEn(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_sigsIn_break),
    .io_rr(x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_rr)
  );
  assign _T_545 = RetimeWrapper_io_out; // @[package.scala 96:25:@8010.4 package.scala 96:25:@8011.4]
  assign _T_551 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@8018.4 package.scala 96:25:@8019.4]
  assign _T_554 = ~ _T_551; // @[SpatialBlocks.scala 110:93:@8021.4]
  assign _T_620 = x343_inr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@8295.4]
  assign _T_637 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@8329.4 package.scala 96:25:@8330.4]
  assign _T_643 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@8337.4 package.scala 96:25:@8338.4]
  assign _T_646 = ~ _T_643; // @[SpatialBlocks.scala 110:93:@8340.4]
  assign io_in_x269_argOut_port_0_valid = x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x269_argOut_port_0_valid; // @[MemInterfaceType.scala 317:38:@8541.4]
  assign io_in_x269_argOut_port_0_bits = x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x269_argOut_port_0_bits; // @[MemInterfaceType.scala 317:38:@8540.4]
  assign io_in_x257_argOut_port_0_valid = x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x257_argOut_port_0_valid; // @[MemInterfaceType.scala 317:38:@8546.4]
  assign io_in_x257_argOut_port_0_bits = x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x257_argOut_port_0_bits; // @[MemInterfaceType.scala 317:38:@8545.4]
  assign io_in_x261_argOut_port_0_valid = x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x261_argOut_port_0_valid; // @[MemInterfaceType.scala 317:38:@8551.4]
  assign io_in_x261_argOut_port_0_bits = x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x261_argOut_port_0_bits; // @[MemInterfaceType.scala 317:38:@8550.4]
  assign io_in_x265_argOut_port_0_valid = x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x265_argOut_port_0_valid; // @[MemInterfaceType.scala 317:38:@8556.4]
  assign io_in_x265_argOut_port_0_bits = x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x265_argOut_port_0_bits; // @[MemInterfaceType.scala 317:38:@8555.4]
  assign io_in_x270_argOut_port_0_valid = x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x270_argOut_port_0_valid; // @[MemInterfaceType.scala 317:38:@8561.4]
  assign io_in_x270_argOut_port_0_bits = x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x270_argOut_port_0_bits; // @[MemInterfaceType.scala 317:38:@8560.4]
  assign io_in_x260_argOut_port_0_valid = x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x260_argOut_port_0_valid; // @[MemInterfaceType.scala 317:38:@8566.4]
  assign io_in_x260_argOut_port_0_bits = x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x260_argOut_port_0_bits; // @[MemInterfaceType.scala 317:38:@8565.4]
  assign io_in_x275_ready = x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_in_x275_ready; // @[sm_x294_outr_UnitPipe.scala 57:23:@8193.4]
  assign io_in_x256_argOut_port_0_valid = x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x256_argOut_port_0_valid; // @[MemInterfaceType.scala 317:38:@8571.4]
  assign io_in_x256_argOut_port_0_bits = x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x256_argOut_port_0_bits; // @[MemInterfaceType.scala 317:38:@8570.4]
  assign io_in_x266_argOut_port_0_valid = x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x266_argOut_port_0_valid; // @[MemInterfaceType.scala 317:38:@8576.4]
  assign io_in_x266_argOut_port_0_bits = x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x266_argOut_port_0_bits; // @[MemInterfaceType.scala 317:38:@8575.4]
  assign io_in_x264_argOut_port_0_valid = x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x264_argOut_port_0_valid; // @[MemInterfaceType.scala 317:38:@8581.4]
  assign io_in_x264_argOut_port_0_bits = x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x264_argOut_port_0_bits; // @[MemInterfaceType.scala 317:38:@8580.4]
  assign io_in_x259_argOut_port_0_valid = x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x259_argOut_port_0_valid; // @[MemInterfaceType.scala 317:38:@8586.4]
  assign io_in_x259_argOut_port_0_bits = x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x259_argOut_port_0_bits; // @[MemInterfaceType.scala 317:38:@8585.4]
  assign io_in_x274_valid = x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_in_x274_valid; // @[sm_x294_outr_UnitPipe.scala 56:23:@8189.4]
  assign io_in_x274_bits_addr = x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_in_x274_bits_addr; // @[sm_x294_outr_UnitPipe.scala 56:23:@8188.4]
  assign io_in_x274_bits_size = x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_in_x274_bits_size; // @[sm_x294_outr_UnitPipe.scala 56:23:@8187.4]
  assign io_in_x267_argOut_port_0_valid = x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x267_argOut_port_0_valid; // @[MemInterfaceType.scala 317:38:@8591.4]
  assign io_in_x267_argOut_port_0_bits = x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x267_argOut_port_0_bits; // @[MemInterfaceType.scala 317:38:@8590.4]
  assign io_in_x255_argOut_port_0_valid = x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x255_argOut_port_0_valid; // @[MemInterfaceType.scala 317:38:@8596.4]
  assign io_in_x255_argOut_port_0_bits = x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x255_argOut_port_0_bits; // @[MemInterfaceType.scala 317:38:@8595.4]
  assign io_in_x263_argOut_port_0_valid = x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x263_argOut_port_0_valid; // @[MemInterfaceType.scala 317:38:@8601.4]
  assign io_in_x263_argOut_port_0_bits = x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x263_argOut_port_0_bits; // @[MemInterfaceType.scala 317:38:@8600.4]
  assign io_in_x258_argOut_port_0_valid = x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x258_argOut_port_0_valid; // @[MemInterfaceType.scala 317:38:@8606.4]
  assign io_in_x258_argOut_port_0_bits = x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x258_argOut_port_0_bits; // @[MemInterfaceType.scala 317:38:@8605.4]
  assign io_in_x262_argOut_port_0_valid = x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x262_argOut_port_0_valid; // @[MemInterfaceType.scala 317:38:@8611.4]
  assign io_in_x262_argOut_port_0_bits = x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x262_argOut_port_0_bits; // @[MemInterfaceType.scala 317:38:@8610.4]
  assign io_in_x268_argOut_port_0_valid = x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x268_argOut_port_0_valid; // @[MemInterfaceType.scala 317:38:@8696.4]
  assign io_in_x268_argOut_port_0_bits = x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x268_argOut_port_0_bits; // @[MemInterfaceType.scala 317:38:@8695.4]
  assign io_sigsOut_smDoneIn_0 = x294_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 127:53:@8028.4]
  assign io_sigsOut_smDoneIn_1 = x343_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 127:53:@8347.4]
  assign x273_a_0_clock = clock; // @[:@7805.4]
  assign x273_a_0_reset = reset; // @[:@7806.4]
  assign x273_a_0_io_rPort_15_en_0 = x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_15_en_0; // @[MemInterfaceType.scala 66:44:@8687.4]
  assign x273_a_0_io_rPort_14_en_0 = x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_14_en_0; // @[MemInterfaceType.scala 66:44:@8662.4]
  assign x273_a_0_io_rPort_13_en_0 = x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_13_en_0; // @[MemInterfaceType.scala 66:44:@8632.4]
  assign x273_a_0_io_rPort_12_en_0 = x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_12_en_0; // @[MemInterfaceType.scala 66:44:@8657.4]
  assign x273_a_0_io_rPort_11_en_0 = x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_11_en_0; // @[MemInterfaceType.scala 66:44:@8677.4]
  assign x273_a_0_io_rPort_10_en_0 = x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_10_en_0; // @[MemInterfaceType.scala 66:44:@8642.4]
  assign x273_a_0_io_rPort_9_en_0 = x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_9_en_0; // @[MemInterfaceType.scala 66:44:@8617.4]
  assign x273_a_0_io_rPort_8_en_0 = x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_8_en_0; // @[MemInterfaceType.scala 66:44:@8647.4]
  assign x273_a_0_io_rPort_7_en_0 = x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_7_en_0; // @[MemInterfaceType.scala 66:44:@8622.4]
  assign x273_a_0_io_rPort_6_en_0 = x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_6_en_0; // @[MemInterfaceType.scala 66:44:@8672.4]
  assign x273_a_0_io_rPort_5_en_0 = x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_5_en_0; // @[MemInterfaceType.scala 66:44:@8682.4]
  assign x273_a_0_io_rPort_4_en_0 = x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_4_en_0; // @[MemInterfaceType.scala 66:44:@8637.4]
  assign x273_a_0_io_rPort_3_en_0 = x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_3_en_0; // @[MemInterfaceType.scala 66:44:@8652.4]
  assign x273_a_0_io_rPort_2_en_0 = x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_2_en_0; // @[MemInterfaceType.scala 66:44:@8667.4]
  assign x273_a_0_io_rPort_1_en_0 = x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_1_en_0; // @[MemInterfaceType.scala 66:44:@8627.4]
  assign x273_a_0_io_rPort_0_en_0 = x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@8692.4]
  assign x273_a_0_io_wPort_0_banks_0 = x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_in_x273_a_0_wPort_0_banks_0; // @[MemInterfaceType.scala 67:44:@8185.4]
  assign x273_a_0_io_wPort_0_ofs_0 = x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_in_x273_a_0_wPort_0_ofs_0; // @[MemInterfaceType.scala 67:44:@8184.4]
  assign x273_a_0_io_wPort_0_data_0 = x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_in_x273_a_0_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@8183.4]
  assign x273_a_0_io_wPort_0_en_0 = x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_in_x273_a_0_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@8179.4]
  assign x294_outr_UnitPipe_sm_clock = clock; // @[:@7944.4]
  assign x294_outr_UnitPipe_sm_reset = reset; // @[:@7945.4]
  assign x294_outr_UnitPipe_sm_io_enable = _T_545 & _T_554; // @[SpatialBlocks.scala 112:18:@8025.4]
  assign x294_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 114:21:@8027.4]
  assign x294_outr_UnitPipe_sm_io_doneIn_0 = x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 102:67:@7995.4]
  assign x294_outr_UnitPipe_sm_io_doneIn_1 = x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 102:67:@7996.4]
  assign x294_outr_UnitPipe_sm_io_ctrCopyDone_0 = x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 132:80:@8039.4]
  assign x294_outr_UnitPipe_sm_io_ctrCopyDone_1 = x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[SpatialBlocks.scala 132:80:@8040.4]
  assign RetimeWrapper_clock = clock; // @[:@8006.4]
  assign RetimeWrapper_reset = reset; // @[:@8007.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@8009.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@8008.4]
  assign RetimeWrapper_1_clock = clock; // @[:@8014.4]
  assign RetimeWrapper_1_reset = reset; // @[:@8015.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@8017.4]
  assign RetimeWrapper_1_io_in = x294_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@8016.4]
  assign x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_clock = clock; // @[:@8042.4]
  assign x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_reset = reset; // @[:@8043.4]
  assign x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_in_x254_in_number = io_in_x254_in_number; // @[sm_x294_outr_UnitPipe.scala 55:26:@8186.4]
  assign x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_in_x274_ready = io_in_x274_ready; // @[sm_x294_outr_UnitPipe.scala 56:23:@8190.4]
  assign x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_in_x275_valid = io_in_x275_valid; // @[sm_x294_outr_UnitPipe.scala 57:23:@8192.4]
  assign x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_in_x275_bits_rdata_0 = io_in_x275_bits_rdata_0; // @[sm_x294_outr_UnitPipe.scala 57:23:@8191.4]
  assign x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x294_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x294_outr_UnitPipe.scala 97:22:@8209.4]
  assign x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1 = x294_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x294_outr_UnitPipe.scala 97:22:@8210.4]
  assign x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x294_outr_UnitPipe_sm_io_childAck_0; // @[sm_x294_outr_UnitPipe.scala 97:22:@8205.4]
  assign x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1 = x294_outr_UnitPipe_sm_io_childAck_1; // @[sm_x294_outr_UnitPipe.scala 97:22:@8206.4]
  assign x294_outr_UnitPipe_kernelx294_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x294_outr_UnitPipe.scala 96:18:@8194.4]
  assign x343_inr_UnitPipe_sm_clock = clock; // @[:@8268.4]
  assign x343_inr_UnitPipe_sm_reset = reset; // @[:@8269.4]
  assign x343_inr_UnitPipe_sm_io_enable = _T_637 & _T_646; // @[SpatialBlocks.scala 112:18:@8344.4]
  assign x343_inr_UnitPipe_sm_io_ctrDone = x343_inr_UnitPipe_sm_io_ctrInc & _T_623; // @[sm_RootController.scala 156:39:@8299.4]
  assign x343_inr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 114:21:@8346.4]
  assign x343_inr_UnitPipe_sm_io_break = 1'h0; // @[sm_RootController.scala 160:37:@8305.4]
  assign RetimeWrapper_2_clock = clock; // @[:@8325.4]
  assign RetimeWrapper_2_reset = reset; // @[:@8326.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@8328.4]
  assign RetimeWrapper_2_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@8327.4]
  assign RetimeWrapper_3_clock = clock; // @[:@8333.4]
  assign RetimeWrapper_3_reset = reset; // @[:@8334.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@8336.4]
  assign RetimeWrapper_3_io_in = x343_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@8335.4]
  assign x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_clock = clock; // @[:@8359.4]
  assign x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_reset = reset; // @[:@8360.4]
  assign x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_15_output_0 = x273_a_0_io_rPort_15_output_0; // @[MemInterfaceType.scala 66:44:@8685.4]
  assign x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_14_output_0 = x273_a_0_io_rPort_14_output_0; // @[MemInterfaceType.scala 66:44:@8660.4]
  assign x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_13_output_0 = x273_a_0_io_rPort_13_output_0; // @[MemInterfaceType.scala 66:44:@8630.4]
  assign x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_12_output_0 = x273_a_0_io_rPort_12_output_0; // @[MemInterfaceType.scala 66:44:@8655.4]
  assign x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_11_output_0 = x273_a_0_io_rPort_11_output_0; // @[MemInterfaceType.scala 66:44:@8675.4]
  assign x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_10_output_0 = x273_a_0_io_rPort_10_output_0; // @[MemInterfaceType.scala 66:44:@8640.4]
  assign x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_9_output_0 = x273_a_0_io_rPort_9_output_0; // @[MemInterfaceType.scala 66:44:@8615.4]
  assign x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_8_output_0 = x273_a_0_io_rPort_8_output_0; // @[MemInterfaceType.scala 66:44:@8645.4]
  assign x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_7_output_0 = x273_a_0_io_rPort_7_output_0; // @[MemInterfaceType.scala 66:44:@8620.4]
  assign x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_6_output_0 = x273_a_0_io_rPort_6_output_0; // @[MemInterfaceType.scala 66:44:@8670.4]
  assign x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_5_output_0 = x273_a_0_io_rPort_5_output_0; // @[MemInterfaceType.scala 66:44:@8680.4]
  assign x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_4_output_0 = x273_a_0_io_rPort_4_output_0; // @[MemInterfaceType.scala 66:44:@8635.4]
  assign x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_3_output_0 = x273_a_0_io_rPort_3_output_0; // @[MemInterfaceType.scala 66:44:@8650.4]
  assign x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_2_output_0 = x273_a_0_io_rPort_2_output_0; // @[MemInterfaceType.scala 66:44:@8665.4]
  assign x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_1_output_0 = x273_a_0_io_rPort_1_output_0; // @[MemInterfaceType.scala 66:44:@8625.4]
  assign x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_in_x273_a_0_rPort_0_output_0 = x273_a_0_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@8690.4]
  assign x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_sigsIn_datapathEn = x343_inr_UnitPipe_sm_io_datapathEn; // @[sm_x343_inr_UnitPipe.scala 269:22:@8712.4]
  assign x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_sigsIn_break = x343_inr_UnitPipe_sm_io_break; // @[sm_x343_inr_UnitPipe.scala 269:22:@8710.4]
  assign x343_inr_UnitPipe_kernelx343_inr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x343_inr_UnitPipe.scala 268:18:@8700.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_623 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_623 <= 1'h0;
    end else begin
      _T_623 <= _T_620;
    end
  end
endmodule
module AccelTop( // @[:@8727.2]
  input         clock, // @[:@8728.4]
  input         reset, // @[:@8729.4]
  input         io_enable, // @[:@8730.4]
  output        io_done, // @[:@8730.4]
  input         io_reset, // @[:@8730.4]
  input         io_memStreams_loads_0_cmd_ready, // @[:@8730.4]
  output        io_memStreams_loads_0_cmd_valid, // @[:@8730.4]
  output [63:0] io_memStreams_loads_0_cmd_bits_addr, // @[:@8730.4]
  output [31:0] io_memStreams_loads_0_cmd_bits_size, // @[:@8730.4]
  output        io_memStreams_loads_0_data_ready, // @[:@8730.4]
  input         io_memStreams_loads_0_data_valid, // @[:@8730.4]
  input  [31:0] io_memStreams_loads_0_data_bits_rdata_0, // @[:@8730.4]
  input         io_memStreams_stores_0_cmd_ready, // @[:@8730.4]
  output        io_memStreams_stores_0_cmd_valid, // @[:@8730.4]
  output [63:0] io_memStreams_stores_0_cmd_bits_addr, // @[:@8730.4]
  output [31:0] io_memStreams_stores_0_cmd_bits_size, // @[:@8730.4]
  input         io_memStreams_stores_0_data_ready, // @[:@8730.4]
  output        io_memStreams_stores_0_data_valid, // @[:@8730.4]
  output [31:0] io_memStreams_stores_0_data_bits_wdata_0, // @[:@8730.4]
  output [31:0] io_memStreams_stores_0_data_bits_wdata_1, // @[:@8730.4]
  output [31:0] io_memStreams_stores_0_data_bits_wdata_2, // @[:@8730.4]
  output [31:0] io_memStreams_stores_0_data_bits_wdata_3, // @[:@8730.4]
  output [31:0] io_memStreams_stores_0_data_bits_wdata_4, // @[:@8730.4]
  output [31:0] io_memStreams_stores_0_data_bits_wdata_5, // @[:@8730.4]
  output [31:0] io_memStreams_stores_0_data_bits_wdata_6, // @[:@8730.4]
  output [31:0] io_memStreams_stores_0_data_bits_wdata_7, // @[:@8730.4]
  output [31:0] io_memStreams_stores_0_data_bits_wdata_8, // @[:@8730.4]
  output [31:0] io_memStreams_stores_0_data_bits_wdata_9, // @[:@8730.4]
  output [31:0] io_memStreams_stores_0_data_bits_wdata_10, // @[:@8730.4]
  output [31:0] io_memStreams_stores_0_data_bits_wdata_11, // @[:@8730.4]
  output [31:0] io_memStreams_stores_0_data_bits_wdata_12, // @[:@8730.4]
  output [31:0] io_memStreams_stores_0_data_bits_wdata_13, // @[:@8730.4]
  output [31:0] io_memStreams_stores_0_data_bits_wdata_14, // @[:@8730.4]
  output [31:0] io_memStreams_stores_0_data_bits_wdata_15, // @[:@8730.4]
  output [15:0] io_memStreams_stores_0_data_bits_wstrb, // @[:@8730.4]
  output        io_memStreams_stores_0_wresp_ready, // @[:@8730.4]
  input         io_memStreams_stores_0_wresp_valid, // @[:@8730.4]
  input         io_memStreams_stores_0_wresp_bits, // @[:@8730.4]
  input         io_memStreams_gathers_0_cmd_ready, // @[:@8730.4]
  output        io_memStreams_gathers_0_cmd_valid, // @[:@8730.4]
  output [63:0] io_memStreams_gathers_0_cmd_bits_addr_0, // @[:@8730.4]
  output [63:0] io_memStreams_gathers_0_cmd_bits_addr_1, // @[:@8730.4]
  output [63:0] io_memStreams_gathers_0_cmd_bits_addr_2, // @[:@8730.4]
  output [63:0] io_memStreams_gathers_0_cmd_bits_addr_3, // @[:@8730.4]
  output [63:0] io_memStreams_gathers_0_cmd_bits_addr_4, // @[:@8730.4]
  output [63:0] io_memStreams_gathers_0_cmd_bits_addr_5, // @[:@8730.4]
  output [63:0] io_memStreams_gathers_0_cmd_bits_addr_6, // @[:@8730.4]
  output [63:0] io_memStreams_gathers_0_cmd_bits_addr_7, // @[:@8730.4]
  output [63:0] io_memStreams_gathers_0_cmd_bits_addr_8, // @[:@8730.4]
  output [63:0] io_memStreams_gathers_0_cmd_bits_addr_9, // @[:@8730.4]
  output [63:0] io_memStreams_gathers_0_cmd_bits_addr_10, // @[:@8730.4]
  output [63:0] io_memStreams_gathers_0_cmd_bits_addr_11, // @[:@8730.4]
  output [63:0] io_memStreams_gathers_0_cmd_bits_addr_12, // @[:@8730.4]
  output [63:0] io_memStreams_gathers_0_cmd_bits_addr_13, // @[:@8730.4]
  output [63:0] io_memStreams_gathers_0_cmd_bits_addr_14, // @[:@8730.4]
  output [63:0] io_memStreams_gathers_0_cmd_bits_addr_15, // @[:@8730.4]
  output        io_memStreams_gathers_0_data_ready, // @[:@8730.4]
  input         io_memStreams_gathers_0_data_valid, // @[:@8730.4]
  input  [31:0] io_memStreams_gathers_0_data_bits_0, // @[:@8730.4]
  input  [31:0] io_memStreams_gathers_0_data_bits_1, // @[:@8730.4]
  input  [31:0] io_memStreams_gathers_0_data_bits_2, // @[:@8730.4]
  input  [31:0] io_memStreams_gathers_0_data_bits_3, // @[:@8730.4]
  input  [31:0] io_memStreams_gathers_0_data_bits_4, // @[:@8730.4]
  input  [31:0] io_memStreams_gathers_0_data_bits_5, // @[:@8730.4]
  input  [31:0] io_memStreams_gathers_0_data_bits_6, // @[:@8730.4]
  input  [31:0] io_memStreams_gathers_0_data_bits_7, // @[:@8730.4]
  input  [31:0] io_memStreams_gathers_0_data_bits_8, // @[:@8730.4]
  input  [31:0] io_memStreams_gathers_0_data_bits_9, // @[:@8730.4]
  input  [31:0] io_memStreams_gathers_0_data_bits_10, // @[:@8730.4]
  input  [31:0] io_memStreams_gathers_0_data_bits_11, // @[:@8730.4]
  input  [31:0] io_memStreams_gathers_0_data_bits_12, // @[:@8730.4]
  input  [31:0] io_memStreams_gathers_0_data_bits_13, // @[:@8730.4]
  input  [31:0] io_memStreams_gathers_0_data_bits_14, // @[:@8730.4]
  input  [31:0] io_memStreams_gathers_0_data_bits_15, // @[:@8730.4]
  input         io_memStreams_scatters_0_cmd_ready, // @[:@8730.4]
  output        io_memStreams_scatters_0_cmd_valid, // @[:@8730.4]
  output [63:0] io_memStreams_scatters_0_cmd_bits_addr_addr_0, // @[:@8730.4]
  output [63:0] io_memStreams_scatters_0_cmd_bits_addr_addr_1, // @[:@8730.4]
  output [63:0] io_memStreams_scatters_0_cmd_bits_addr_addr_2, // @[:@8730.4]
  output [63:0] io_memStreams_scatters_0_cmd_bits_addr_addr_3, // @[:@8730.4]
  output [63:0] io_memStreams_scatters_0_cmd_bits_addr_addr_4, // @[:@8730.4]
  output [63:0] io_memStreams_scatters_0_cmd_bits_addr_addr_5, // @[:@8730.4]
  output [63:0] io_memStreams_scatters_0_cmd_bits_addr_addr_6, // @[:@8730.4]
  output [63:0] io_memStreams_scatters_0_cmd_bits_addr_addr_7, // @[:@8730.4]
  output [63:0] io_memStreams_scatters_0_cmd_bits_addr_addr_8, // @[:@8730.4]
  output [63:0] io_memStreams_scatters_0_cmd_bits_addr_addr_9, // @[:@8730.4]
  output [63:0] io_memStreams_scatters_0_cmd_bits_addr_addr_10, // @[:@8730.4]
  output [63:0] io_memStreams_scatters_0_cmd_bits_addr_addr_11, // @[:@8730.4]
  output [63:0] io_memStreams_scatters_0_cmd_bits_addr_addr_12, // @[:@8730.4]
  output [63:0] io_memStreams_scatters_0_cmd_bits_addr_addr_13, // @[:@8730.4]
  output [63:0] io_memStreams_scatters_0_cmd_bits_addr_addr_14, // @[:@8730.4]
  output [63:0] io_memStreams_scatters_0_cmd_bits_addr_addr_15, // @[:@8730.4]
  output [31:0] io_memStreams_scatters_0_cmd_bits_wdata_0, // @[:@8730.4]
  output [31:0] io_memStreams_scatters_0_cmd_bits_wdata_1, // @[:@8730.4]
  output [31:0] io_memStreams_scatters_0_cmd_bits_wdata_2, // @[:@8730.4]
  output [31:0] io_memStreams_scatters_0_cmd_bits_wdata_3, // @[:@8730.4]
  output [31:0] io_memStreams_scatters_0_cmd_bits_wdata_4, // @[:@8730.4]
  output [31:0] io_memStreams_scatters_0_cmd_bits_wdata_5, // @[:@8730.4]
  output [31:0] io_memStreams_scatters_0_cmd_bits_wdata_6, // @[:@8730.4]
  output [31:0] io_memStreams_scatters_0_cmd_bits_wdata_7, // @[:@8730.4]
  output [31:0] io_memStreams_scatters_0_cmd_bits_wdata_8, // @[:@8730.4]
  output [31:0] io_memStreams_scatters_0_cmd_bits_wdata_9, // @[:@8730.4]
  output [31:0] io_memStreams_scatters_0_cmd_bits_wdata_10, // @[:@8730.4]
  output [31:0] io_memStreams_scatters_0_cmd_bits_wdata_11, // @[:@8730.4]
  output [31:0] io_memStreams_scatters_0_cmd_bits_wdata_12, // @[:@8730.4]
  output [31:0] io_memStreams_scatters_0_cmd_bits_wdata_13, // @[:@8730.4]
  output [31:0] io_memStreams_scatters_0_cmd_bits_wdata_14, // @[:@8730.4]
  output [31:0] io_memStreams_scatters_0_cmd_bits_wdata_15, // @[:@8730.4]
  output        io_memStreams_scatters_0_wresp_ready, // @[:@8730.4]
  input         io_memStreams_scatters_0_wresp_valid, // @[:@8730.4]
  input         io_memStreams_scatters_0_wresp_bits, // @[:@8730.4]
  output        io_heap_0_req_valid, // @[:@8730.4]
  output        io_heap_0_req_bits_allocDealloc, // @[:@8730.4]
  output [63:0] io_heap_0_req_bits_sizeAddr, // @[:@8730.4]
  input         io_heap_0_resp_valid, // @[:@8730.4]
  input         io_heap_0_resp_bits_allocDealloc, // @[:@8730.4]
  input  [63:0] io_heap_0_resp_bits_sizeAddr, // @[:@8730.4]
  input  [63:0] io_argIns_0, // @[:@8730.4]
  input         io_argOuts_0_port_ready, // @[:@8730.4]
  output        io_argOuts_0_port_valid, // @[:@8730.4]
  output [63:0] io_argOuts_0_port_bits, // @[:@8730.4]
  input  [63:0] io_argOuts_0_echo, // @[:@8730.4]
  input         io_argOuts_1_port_ready, // @[:@8730.4]
  output        io_argOuts_1_port_valid, // @[:@8730.4]
  output [63:0] io_argOuts_1_port_bits, // @[:@8730.4]
  input  [63:0] io_argOuts_1_echo, // @[:@8730.4]
  input         io_argOuts_2_port_ready, // @[:@8730.4]
  output        io_argOuts_2_port_valid, // @[:@8730.4]
  output [63:0] io_argOuts_2_port_bits, // @[:@8730.4]
  input  [63:0] io_argOuts_2_echo, // @[:@8730.4]
  input         io_argOuts_3_port_ready, // @[:@8730.4]
  output        io_argOuts_3_port_valid, // @[:@8730.4]
  output [63:0] io_argOuts_3_port_bits, // @[:@8730.4]
  input  [63:0] io_argOuts_3_echo, // @[:@8730.4]
  input         io_argOuts_4_port_ready, // @[:@8730.4]
  output        io_argOuts_4_port_valid, // @[:@8730.4]
  output [63:0] io_argOuts_4_port_bits, // @[:@8730.4]
  input  [63:0] io_argOuts_4_echo, // @[:@8730.4]
  input         io_argOuts_5_port_ready, // @[:@8730.4]
  output        io_argOuts_5_port_valid, // @[:@8730.4]
  output [63:0] io_argOuts_5_port_bits, // @[:@8730.4]
  input  [63:0] io_argOuts_5_echo, // @[:@8730.4]
  input         io_argOuts_6_port_ready, // @[:@8730.4]
  output        io_argOuts_6_port_valid, // @[:@8730.4]
  output [63:0] io_argOuts_6_port_bits, // @[:@8730.4]
  input  [63:0] io_argOuts_6_echo, // @[:@8730.4]
  input         io_argOuts_7_port_ready, // @[:@8730.4]
  output        io_argOuts_7_port_valid, // @[:@8730.4]
  output [63:0] io_argOuts_7_port_bits, // @[:@8730.4]
  input  [63:0] io_argOuts_7_echo, // @[:@8730.4]
  input         io_argOuts_8_port_ready, // @[:@8730.4]
  output        io_argOuts_8_port_valid, // @[:@8730.4]
  output [63:0] io_argOuts_8_port_bits, // @[:@8730.4]
  input  [63:0] io_argOuts_8_echo, // @[:@8730.4]
  input         io_argOuts_9_port_ready, // @[:@8730.4]
  output        io_argOuts_9_port_valid, // @[:@8730.4]
  output [63:0] io_argOuts_9_port_bits, // @[:@8730.4]
  input  [63:0] io_argOuts_9_echo, // @[:@8730.4]
  input         io_argOuts_10_port_ready, // @[:@8730.4]
  output        io_argOuts_10_port_valid, // @[:@8730.4]
  output [63:0] io_argOuts_10_port_bits, // @[:@8730.4]
  input  [63:0] io_argOuts_10_echo, // @[:@8730.4]
  input         io_argOuts_11_port_ready, // @[:@8730.4]
  output        io_argOuts_11_port_valid, // @[:@8730.4]
  output [63:0] io_argOuts_11_port_bits, // @[:@8730.4]
  input  [63:0] io_argOuts_11_echo, // @[:@8730.4]
  input         io_argOuts_12_port_ready, // @[:@8730.4]
  output        io_argOuts_12_port_valid, // @[:@8730.4]
  output [63:0] io_argOuts_12_port_bits, // @[:@8730.4]
  input  [63:0] io_argOuts_12_echo, // @[:@8730.4]
  input         io_argOuts_13_port_ready, // @[:@8730.4]
  output        io_argOuts_13_port_valid, // @[:@8730.4]
  output [63:0] io_argOuts_13_port_bits, // @[:@8730.4]
  input  [63:0] io_argOuts_13_echo, // @[:@8730.4]
  input         io_argOuts_14_port_ready, // @[:@8730.4]
  output        io_argOuts_14_port_valid, // @[:@8730.4]
  output [63:0] io_argOuts_14_port_bits, // @[:@8730.4]
  input  [63:0] io_argOuts_14_echo, // @[:@8730.4]
  input         io_argOuts_15_port_ready, // @[:@8730.4]
  output        io_argOuts_15_port_valid, // @[:@8730.4]
  output [63:0] io_argOuts_15_port_bits, // @[:@8730.4]
  input  [63:0] io_argOuts_15_echo // @[:@8730.4]
);
  wire  SingleCounter_clock; // @[Main.scala 113:32:@9045.4]
  wire  SingleCounter_reset; // @[Main.scala 113:32:@9045.4]
  wire  SingleCounter_io_input_reset; // @[Main.scala 113:32:@9045.4]
  wire  SingleCounter_io_output_done; // @[Main.scala 113:32:@9045.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@9063.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@9063.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@9063.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@9063.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@9063.4]
  wire  SRFF_clock; // @[Main.scala 117:28:@9072.4]
  wire  SRFF_reset; // @[Main.scala 117:28:@9072.4]
  wire  SRFF_io_input_set; // @[Main.scala 117:28:@9072.4]
  wire  SRFF_io_input_reset; // @[Main.scala 117:28:@9072.4]
  wire  SRFF_io_input_asyn_reset; // @[Main.scala 117:28:@9072.4]
  wire  SRFF_io_output; // @[Main.scala 117:28:@9072.4]
  wire  RootController_sm_clock; // @[sm_RootController.scala 34:18:@9115.4]
  wire  RootController_sm_reset; // @[sm_RootController.scala 34:18:@9115.4]
  wire  RootController_sm_io_enable; // @[sm_RootController.scala 34:18:@9115.4]
  wire  RootController_sm_io_done; // @[sm_RootController.scala 34:18:@9115.4]
  wire  RootController_sm_io_rst; // @[sm_RootController.scala 34:18:@9115.4]
  wire  RootController_sm_io_ctrDone; // @[sm_RootController.scala 34:18:@9115.4]
  wire  RootController_sm_io_ctrInc; // @[sm_RootController.scala 34:18:@9115.4]
  wire  RootController_sm_io_doneIn_0; // @[sm_RootController.scala 34:18:@9115.4]
  wire  RootController_sm_io_doneIn_1; // @[sm_RootController.scala 34:18:@9115.4]
  wire  RootController_sm_io_enableOut_0; // @[sm_RootController.scala 34:18:@9115.4]
  wire  RootController_sm_io_enableOut_1; // @[sm_RootController.scala 34:18:@9115.4]
  wire  RootController_sm_io_childAck_0; // @[sm_RootController.scala 34:18:@9115.4]
  wire  RootController_sm_io_childAck_1; // @[sm_RootController.scala 34:18:@9115.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@9152.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@9152.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@9152.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@9152.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@9152.4]
  wire  RootController_kernelRootController_concrete1_clock; // @[sm_RootController.scala 165:24:@9216.4]
  wire  RootController_kernelRootController_concrete1_reset; // @[sm_RootController.scala 165:24:@9216.4]
  wire  RootController_kernelRootController_concrete1_io_in_x269_argOut_port_0_valid; // @[sm_RootController.scala 165:24:@9216.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x269_argOut_port_0_bits; // @[sm_RootController.scala 165:24:@9216.4]
  wire  RootController_kernelRootController_concrete1_io_in_x257_argOut_port_0_valid; // @[sm_RootController.scala 165:24:@9216.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x257_argOut_port_0_bits; // @[sm_RootController.scala 165:24:@9216.4]
  wire  RootController_kernelRootController_concrete1_io_in_x261_argOut_port_0_valid; // @[sm_RootController.scala 165:24:@9216.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x261_argOut_port_0_bits; // @[sm_RootController.scala 165:24:@9216.4]
  wire  RootController_kernelRootController_concrete1_io_in_x265_argOut_port_0_valid; // @[sm_RootController.scala 165:24:@9216.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x265_argOut_port_0_bits; // @[sm_RootController.scala 165:24:@9216.4]
  wire  RootController_kernelRootController_concrete1_io_in_x270_argOut_port_0_valid; // @[sm_RootController.scala 165:24:@9216.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x270_argOut_port_0_bits; // @[sm_RootController.scala 165:24:@9216.4]
  wire  RootController_kernelRootController_concrete1_io_in_x260_argOut_port_0_valid; // @[sm_RootController.scala 165:24:@9216.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x260_argOut_port_0_bits; // @[sm_RootController.scala 165:24:@9216.4]
  wire  RootController_kernelRootController_concrete1_io_in_x275_ready; // @[sm_RootController.scala 165:24:@9216.4]
  wire  RootController_kernelRootController_concrete1_io_in_x275_valid; // @[sm_RootController.scala 165:24:@9216.4]
  wire [31:0] RootController_kernelRootController_concrete1_io_in_x275_bits_rdata_0; // @[sm_RootController.scala 165:24:@9216.4]
  wire  RootController_kernelRootController_concrete1_io_in_x256_argOut_port_0_valid; // @[sm_RootController.scala 165:24:@9216.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x256_argOut_port_0_bits; // @[sm_RootController.scala 165:24:@9216.4]
  wire  RootController_kernelRootController_concrete1_io_in_x266_argOut_port_0_valid; // @[sm_RootController.scala 165:24:@9216.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x266_argOut_port_0_bits; // @[sm_RootController.scala 165:24:@9216.4]
  wire  RootController_kernelRootController_concrete1_io_in_x264_argOut_port_0_valid; // @[sm_RootController.scala 165:24:@9216.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x264_argOut_port_0_bits; // @[sm_RootController.scala 165:24:@9216.4]
  wire  RootController_kernelRootController_concrete1_io_in_x259_argOut_port_0_valid; // @[sm_RootController.scala 165:24:@9216.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x259_argOut_port_0_bits; // @[sm_RootController.scala 165:24:@9216.4]
  wire  RootController_kernelRootController_concrete1_io_in_x274_ready; // @[sm_RootController.scala 165:24:@9216.4]
  wire  RootController_kernelRootController_concrete1_io_in_x274_valid; // @[sm_RootController.scala 165:24:@9216.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x274_bits_addr; // @[sm_RootController.scala 165:24:@9216.4]
  wire [31:0] RootController_kernelRootController_concrete1_io_in_x274_bits_size; // @[sm_RootController.scala 165:24:@9216.4]
  wire  RootController_kernelRootController_concrete1_io_in_x267_argOut_port_0_valid; // @[sm_RootController.scala 165:24:@9216.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x267_argOut_port_0_bits; // @[sm_RootController.scala 165:24:@9216.4]
  wire  RootController_kernelRootController_concrete1_io_in_x255_argOut_port_0_valid; // @[sm_RootController.scala 165:24:@9216.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x255_argOut_port_0_bits; // @[sm_RootController.scala 165:24:@9216.4]
  wire  RootController_kernelRootController_concrete1_io_in_x263_argOut_port_0_valid; // @[sm_RootController.scala 165:24:@9216.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x263_argOut_port_0_bits; // @[sm_RootController.scala 165:24:@9216.4]
  wire  RootController_kernelRootController_concrete1_io_in_x258_argOut_port_0_valid; // @[sm_RootController.scala 165:24:@9216.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x258_argOut_port_0_bits; // @[sm_RootController.scala 165:24:@9216.4]
  wire  RootController_kernelRootController_concrete1_io_in_x262_argOut_port_0_valid; // @[sm_RootController.scala 165:24:@9216.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x262_argOut_port_0_bits; // @[sm_RootController.scala 165:24:@9216.4]
  wire  RootController_kernelRootController_concrete1_io_in_x268_argOut_port_0_valid; // @[sm_RootController.scala 165:24:@9216.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x268_argOut_port_0_bits; // @[sm_RootController.scala 165:24:@9216.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x254_in_number; // @[sm_RootController.scala 165:24:@9216.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_RootController.scala 165:24:@9216.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_RootController.scala 165:24:@9216.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0; // @[sm_RootController.scala 165:24:@9216.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_1; // @[sm_RootController.scala 165:24:@9216.4]
  wire  RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[sm_RootController.scala 165:24:@9216.4]
  wire  RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_1; // @[sm_RootController.scala 165:24:@9216.4]
  wire  RootController_kernelRootController_concrete1_io_rr; // @[sm_RootController.scala 165:24:@9216.4]
  wire  _T_1007; // @[package.scala 96:25:@9068.4 package.scala 96:25:@9069.4]
  wire  _T_1072; // @[Main.scala 119:44:@9148.4]
  wire  _T_1073; // @[Main.scala 119:53:@9149.4]
  wire  _T_1085; // @[package.scala 100:49:@9169.4]
  reg  _T_1088; // @[package.scala 48:56:@9170.4]
  reg [31:0] _RAND_0;
  SingleCounter SingleCounter ( // @[Main.scala 113:32:@9045.4]
    .clock(SingleCounter_clock),
    .reset(SingleCounter_reset),
    .io_input_reset(SingleCounter_io_input_reset),
    .io_output_done(SingleCounter_io_output_done)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@9063.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  SRFF SRFF ( // @[Main.scala 117:28:@9072.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  RootController_sm RootController_sm ( // @[sm_RootController.scala 34:18:@9115.4]
    .clock(RootController_sm_clock),
    .reset(RootController_sm_reset),
    .io_enable(RootController_sm_io_enable),
    .io_done(RootController_sm_io_done),
    .io_rst(RootController_sm_io_rst),
    .io_ctrDone(RootController_sm_io_ctrDone),
    .io_ctrInc(RootController_sm_io_ctrInc),
    .io_doneIn_0(RootController_sm_io_doneIn_0),
    .io_doneIn_1(RootController_sm_io_doneIn_1),
    .io_enableOut_0(RootController_sm_io_enableOut_0),
    .io_enableOut_1(RootController_sm_io_enableOut_1),
    .io_childAck_0(RootController_sm_io_childAck_0),
    .io_childAck_1(RootController_sm_io_childAck_1)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@9152.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RootController_kernelRootController_concrete1 RootController_kernelRootController_concrete1 ( // @[sm_RootController.scala 165:24:@9216.4]
    .clock(RootController_kernelRootController_concrete1_clock),
    .reset(RootController_kernelRootController_concrete1_reset),
    .io_in_x269_argOut_port_0_valid(RootController_kernelRootController_concrete1_io_in_x269_argOut_port_0_valid),
    .io_in_x269_argOut_port_0_bits(RootController_kernelRootController_concrete1_io_in_x269_argOut_port_0_bits),
    .io_in_x257_argOut_port_0_valid(RootController_kernelRootController_concrete1_io_in_x257_argOut_port_0_valid),
    .io_in_x257_argOut_port_0_bits(RootController_kernelRootController_concrete1_io_in_x257_argOut_port_0_bits),
    .io_in_x261_argOut_port_0_valid(RootController_kernelRootController_concrete1_io_in_x261_argOut_port_0_valid),
    .io_in_x261_argOut_port_0_bits(RootController_kernelRootController_concrete1_io_in_x261_argOut_port_0_bits),
    .io_in_x265_argOut_port_0_valid(RootController_kernelRootController_concrete1_io_in_x265_argOut_port_0_valid),
    .io_in_x265_argOut_port_0_bits(RootController_kernelRootController_concrete1_io_in_x265_argOut_port_0_bits),
    .io_in_x270_argOut_port_0_valid(RootController_kernelRootController_concrete1_io_in_x270_argOut_port_0_valid),
    .io_in_x270_argOut_port_0_bits(RootController_kernelRootController_concrete1_io_in_x270_argOut_port_0_bits),
    .io_in_x260_argOut_port_0_valid(RootController_kernelRootController_concrete1_io_in_x260_argOut_port_0_valid),
    .io_in_x260_argOut_port_0_bits(RootController_kernelRootController_concrete1_io_in_x260_argOut_port_0_bits),
    .io_in_x275_ready(RootController_kernelRootController_concrete1_io_in_x275_ready),
    .io_in_x275_valid(RootController_kernelRootController_concrete1_io_in_x275_valid),
    .io_in_x275_bits_rdata_0(RootController_kernelRootController_concrete1_io_in_x275_bits_rdata_0),
    .io_in_x256_argOut_port_0_valid(RootController_kernelRootController_concrete1_io_in_x256_argOut_port_0_valid),
    .io_in_x256_argOut_port_0_bits(RootController_kernelRootController_concrete1_io_in_x256_argOut_port_0_bits),
    .io_in_x266_argOut_port_0_valid(RootController_kernelRootController_concrete1_io_in_x266_argOut_port_0_valid),
    .io_in_x266_argOut_port_0_bits(RootController_kernelRootController_concrete1_io_in_x266_argOut_port_0_bits),
    .io_in_x264_argOut_port_0_valid(RootController_kernelRootController_concrete1_io_in_x264_argOut_port_0_valid),
    .io_in_x264_argOut_port_0_bits(RootController_kernelRootController_concrete1_io_in_x264_argOut_port_0_bits),
    .io_in_x259_argOut_port_0_valid(RootController_kernelRootController_concrete1_io_in_x259_argOut_port_0_valid),
    .io_in_x259_argOut_port_0_bits(RootController_kernelRootController_concrete1_io_in_x259_argOut_port_0_bits),
    .io_in_x274_ready(RootController_kernelRootController_concrete1_io_in_x274_ready),
    .io_in_x274_valid(RootController_kernelRootController_concrete1_io_in_x274_valid),
    .io_in_x274_bits_addr(RootController_kernelRootController_concrete1_io_in_x274_bits_addr),
    .io_in_x274_bits_size(RootController_kernelRootController_concrete1_io_in_x274_bits_size),
    .io_in_x267_argOut_port_0_valid(RootController_kernelRootController_concrete1_io_in_x267_argOut_port_0_valid),
    .io_in_x267_argOut_port_0_bits(RootController_kernelRootController_concrete1_io_in_x267_argOut_port_0_bits),
    .io_in_x255_argOut_port_0_valid(RootController_kernelRootController_concrete1_io_in_x255_argOut_port_0_valid),
    .io_in_x255_argOut_port_0_bits(RootController_kernelRootController_concrete1_io_in_x255_argOut_port_0_bits),
    .io_in_x263_argOut_port_0_valid(RootController_kernelRootController_concrete1_io_in_x263_argOut_port_0_valid),
    .io_in_x263_argOut_port_0_bits(RootController_kernelRootController_concrete1_io_in_x263_argOut_port_0_bits),
    .io_in_x258_argOut_port_0_valid(RootController_kernelRootController_concrete1_io_in_x258_argOut_port_0_valid),
    .io_in_x258_argOut_port_0_bits(RootController_kernelRootController_concrete1_io_in_x258_argOut_port_0_bits),
    .io_in_x262_argOut_port_0_valid(RootController_kernelRootController_concrete1_io_in_x262_argOut_port_0_valid),
    .io_in_x262_argOut_port_0_bits(RootController_kernelRootController_concrete1_io_in_x262_argOut_port_0_bits),
    .io_in_x268_argOut_port_0_valid(RootController_kernelRootController_concrete1_io_in_x268_argOut_port_0_valid),
    .io_in_x268_argOut_port_0_bits(RootController_kernelRootController_concrete1_io_in_x268_argOut_port_0_bits),
    .io_in_x254_in_number(RootController_kernelRootController_concrete1_io_in_x254_in_number),
    .io_sigsIn_smEnableOuts_0(RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smChildAcks_0(RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsOut_smDoneIn_0(RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_1),
    .io_rr(RootController_kernelRootController_concrete1_io_rr)
  );
  assign _T_1007 = RetimeWrapper_io_out; // @[package.scala 96:25:@9068.4 package.scala 96:25:@9069.4]
  assign _T_1072 = io_enable & _T_1007; // @[Main.scala 119:44:@9148.4]
  assign _T_1073 = ~ SRFF_io_output; // @[Main.scala 119:53:@9149.4]
  assign _T_1085 = RootController_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@9169.4]
  assign io_done = SRFF_io_output; // @[Main.scala 126:17:@9168.4]
  assign io_memStreams_loads_0_cmd_valid = RootController_kernelRootController_concrete1_io_in_x274_valid; // @[sm_RootController.scala 105:23:@9378.4]
  assign io_memStreams_loads_0_cmd_bits_addr = RootController_kernelRootController_concrete1_io_in_x274_bits_addr; // @[sm_RootController.scala 105:23:@9377.4]
  assign io_memStreams_loads_0_cmd_bits_size = RootController_kernelRootController_concrete1_io_in_x274_bits_size; // @[sm_RootController.scala 105:23:@9376.4]
  assign io_memStreams_loads_0_data_ready = RootController_kernelRootController_concrete1_io_in_x275_ready; // @[sm_RootController.scala 96:23:@9355.4]
  assign io_memStreams_stores_0_cmd_valid = 1'h0;
  assign io_memStreams_stores_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_stores_0_cmd_bits_size = 32'h0;
  assign io_memStreams_stores_0_data_valid = 1'h0;
  assign io_memStreams_stores_0_data_bits_wdata_0 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_1 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_2 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_3 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_4 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_5 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_6 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_7 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_8 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_9 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_10 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_11 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_12 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_13 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_14 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_15 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wstrb = 16'h0;
  assign io_memStreams_stores_0_wresp_ready = 1'h0;
  assign io_memStreams_gathers_0_cmd_valid = 1'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_0 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_1 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_2 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_3 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_4 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_5 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_6 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_7 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_8 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_9 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_10 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_11 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_12 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_13 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_14 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_15 = 64'h0;
  assign io_memStreams_gathers_0_data_ready = 1'h0;
  assign io_memStreams_scatters_0_cmd_valid = 1'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_0 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_1 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_2 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_3 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_4 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_5 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_6 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_7 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_8 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_9 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_10 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_11 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_12 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_13 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_14 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_15 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_0 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_1 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_2 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_3 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_4 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_5 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_6 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_7 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_8 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_9 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_10 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_11 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_12 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_13 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_14 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_15 = 32'h0;
  assign io_memStreams_scatters_0_wresp_ready = 1'h0;
  assign io_heap_0_req_valid = 1'h0;
  assign io_heap_0_req_bits_allocDealloc = 1'h0;
  assign io_heap_0_req_bits_sizeAddr = 64'h0;
  assign io_argOuts_0_port_valid = RootController_kernelRootController_concrete1_io_in_x255_argOut_port_0_valid; // @[Main.scala 34:57:@8921.4]
  assign io_argOuts_0_port_bits = RootController_kernelRootController_concrete1_io_in_x255_argOut_port_0_bits; // @[Main.scala 35:56:@8922.4]
  assign io_argOuts_1_port_valid = RootController_kernelRootController_concrete1_io_in_x256_argOut_port_0_valid; // @[Main.scala 39:57:@8929.4]
  assign io_argOuts_1_port_bits = RootController_kernelRootController_concrete1_io_in_x256_argOut_port_0_bits; // @[Main.scala 40:56:@8930.4]
  assign io_argOuts_2_port_valid = RootController_kernelRootController_concrete1_io_in_x257_argOut_port_0_valid; // @[Main.scala 44:57:@8937.4]
  assign io_argOuts_2_port_bits = RootController_kernelRootController_concrete1_io_in_x257_argOut_port_0_bits; // @[Main.scala 45:56:@8938.4]
  assign io_argOuts_3_port_valid = RootController_kernelRootController_concrete1_io_in_x258_argOut_port_0_valid; // @[Main.scala 49:57:@8945.4]
  assign io_argOuts_3_port_bits = RootController_kernelRootController_concrete1_io_in_x258_argOut_port_0_bits; // @[Main.scala 50:56:@8946.4]
  assign io_argOuts_4_port_valid = RootController_kernelRootController_concrete1_io_in_x259_argOut_port_0_valid; // @[Main.scala 54:57:@8953.4]
  assign io_argOuts_4_port_bits = RootController_kernelRootController_concrete1_io_in_x259_argOut_port_0_bits; // @[Main.scala 55:56:@8954.4]
  assign io_argOuts_5_port_valid = RootController_kernelRootController_concrete1_io_in_x260_argOut_port_0_valid; // @[Main.scala 59:57:@8961.4]
  assign io_argOuts_5_port_bits = RootController_kernelRootController_concrete1_io_in_x260_argOut_port_0_bits; // @[Main.scala 60:56:@8962.4]
  assign io_argOuts_6_port_valid = RootController_kernelRootController_concrete1_io_in_x261_argOut_port_0_valid; // @[Main.scala 64:57:@8969.4]
  assign io_argOuts_6_port_bits = RootController_kernelRootController_concrete1_io_in_x261_argOut_port_0_bits; // @[Main.scala 65:56:@8970.4]
  assign io_argOuts_7_port_valid = RootController_kernelRootController_concrete1_io_in_x262_argOut_port_0_valid; // @[Main.scala 69:57:@8977.4]
  assign io_argOuts_7_port_bits = RootController_kernelRootController_concrete1_io_in_x262_argOut_port_0_bits; // @[Main.scala 70:56:@8978.4]
  assign io_argOuts_8_port_valid = RootController_kernelRootController_concrete1_io_in_x263_argOut_port_0_valid; // @[Main.scala 74:57:@8985.4]
  assign io_argOuts_8_port_bits = RootController_kernelRootController_concrete1_io_in_x263_argOut_port_0_bits; // @[Main.scala 75:56:@8986.4]
  assign io_argOuts_9_port_valid = RootController_kernelRootController_concrete1_io_in_x264_argOut_port_0_valid; // @[Main.scala 79:57:@8993.4]
  assign io_argOuts_9_port_bits = RootController_kernelRootController_concrete1_io_in_x264_argOut_port_0_bits; // @[Main.scala 80:56:@8994.4]
  assign io_argOuts_10_port_valid = RootController_kernelRootController_concrete1_io_in_x265_argOut_port_0_valid; // @[Main.scala 84:58:@9001.4]
  assign io_argOuts_10_port_bits = RootController_kernelRootController_concrete1_io_in_x265_argOut_port_0_bits; // @[Main.scala 85:57:@9002.4]
  assign io_argOuts_11_port_valid = RootController_kernelRootController_concrete1_io_in_x266_argOut_port_0_valid; // @[Main.scala 89:58:@9009.4]
  assign io_argOuts_11_port_bits = RootController_kernelRootController_concrete1_io_in_x266_argOut_port_0_bits; // @[Main.scala 90:57:@9010.4]
  assign io_argOuts_12_port_valid = RootController_kernelRootController_concrete1_io_in_x267_argOut_port_0_valid; // @[Main.scala 94:58:@9017.4]
  assign io_argOuts_12_port_bits = RootController_kernelRootController_concrete1_io_in_x267_argOut_port_0_bits; // @[Main.scala 95:57:@9018.4]
  assign io_argOuts_13_port_valid = RootController_kernelRootController_concrete1_io_in_x268_argOut_port_0_valid; // @[Main.scala 99:58:@9025.4]
  assign io_argOuts_13_port_bits = RootController_kernelRootController_concrete1_io_in_x268_argOut_port_0_bits; // @[Main.scala 100:57:@9026.4]
  assign io_argOuts_14_port_valid = RootController_kernelRootController_concrete1_io_in_x269_argOut_port_0_valid; // @[Main.scala 104:58:@9033.4]
  assign io_argOuts_14_port_bits = RootController_kernelRootController_concrete1_io_in_x269_argOut_port_0_bits; // @[Main.scala 105:57:@9034.4]
  assign io_argOuts_15_port_valid = RootController_kernelRootController_concrete1_io_in_x270_argOut_port_0_valid; // @[Main.scala 109:58:@9041.4]
  assign io_argOuts_15_port_bits = RootController_kernelRootController_concrete1_io_in_x270_argOut_port_0_bits; // @[Main.scala 110:57:@9042.4]
  assign SingleCounter_clock = clock; // @[:@9046.4]
  assign SingleCounter_reset = reset; // @[:@9047.4]
  assign SingleCounter_io_input_reset = reset; // @[Main.scala 114:79:@9061.4]
  assign RetimeWrapper_clock = clock; // @[:@9064.4]
  assign RetimeWrapper_reset = reset; // @[:@9065.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@9067.4]
  assign RetimeWrapper_io_in = SingleCounter_io_output_done; // @[package.scala 94:16:@9066.4]
  assign SRFF_clock = clock; // @[:@9073.4]
  assign SRFF_reset = reset; // @[:@9074.4]
  assign SRFF_io_input_set = RootController_sm_io_done; // @[Main.scala 135:29:@9442.4]
  assign SRFF_io_input_reset = RetimeWrapper_1_io_out; // @[Main.scala 124:31:@9166.4]
  assign SRFF_io_input_asyn_reset = RetimeWrapper_1_io_out; // @[Main.scala 125:36:@9167.4]
  assign RootController_sm_clock = clock; // @[:@9116.4]
  assign RootController_sm_reset = reset; // @[:@9117.4]
  assign RootController_sm_io_enable = _T_1072 & _T_1073; // @[Main.scala 123:33:@9165.4 SpatialBlocks.scala 112:18:@9204.4]
  assign RootController_sm_io_rst = RetimeWrapper_1_io_out; // @[SpatialBlocks.scala 106:15:@9198.4]
  assign RootController_sm_io_ctrDone = RootController_sm_io_ctrInc & _T_1088; // @[Main.scala 127:34:@9173.4]
  assign RootController_sm_io_doneIn_0 = RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 102:67:@9193.4]
  assign RootController_sm_io_doneIn_1 = RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 102:67:@9194.4]
  assign RetimeWrapper_1_clock = clock; // @[:@9153.4]
  assign RetimeWrapper_1_reset = reset; // @[:@9154.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@9156.4]
  assign RetimeWrapper_1_io_in = reset | io_reset; // @[package.scala 94:16:@9155.4]
  assign RootController_kernelRootController_concrete1_clock = clock; // @[:@9217.4]
  assign RootController_kernelRootController_concrete1_reset = reset; // @[:@9218.4]
  assign RootController_kernelRootController_concrete1_io_in_x275_valid = io_memStreams_loads_0_data_valid; // @[sm_RootController.scala 96:23:@9354.4]
  assign RootController_kernelRootController_concrete1_io_in_x275_bits_rdata_0 = io_memStreams_loads_0_data_bits_rdata_0; // @[sm_RootController.scala 96:23:@9353.4]
  assign RootController_kernelRootController_concrete1_io_in_x274_ready = io_memStreams_loads_0_cmd_ready; // @[sm_RootController.scala 105:23:@9379.4]
  assign RootController_kernelRootController_concrete1_io_in_x254_in_number = io_argIns_0; // @[sm_RootController.scala 118:26:@9410.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0 = RootController_sm_io_enableOut_0; // @[sm_RootController.scala 169:22:@9421.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_1 = RootController_sm_io_enableOut_1; // @[sm_RootController.scala 169:22:@9422.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0 = RootController_sm_io_childAck_0; // @[sm_RootController.scala 169:22:@9417.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_1 = RootController_sm_io_childAck_1; // @[sm_RootController.scala 169:22:@9418.4]
  assign RootController_kernelRootController_concrete1_io_rr = RetimeWrapper_io_out; // @[sm_RootController.scala 168:18:@9411.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1088 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_1088 <= 1'h0;
    end else begin
      _T_1088 <= _T_1085;
    end
  end
endmodule
module Counter( // @[:@9444.2]
  input        clock, // @[:@9445.4]
  input        reset, // @[:@9446.4]
  input        io_enable, // @[:@9447.4]
  output [5:0] io_out, // @[:@9447.4]
  output [5:0] io_next // @[:@9447.4]
);
  reg [5:0] count; // @[Counter.scala 15:22:@9449.4]
  reg [31:0] _RAND_0;
  wire [6:0] _T_17; // @[Counter.scala 17:24:@9450.4]
  wire [5:0] newCount; // @[Counter.scala 17:24:@9451.4]
  wire [5:0] _GEN_0; // @[Counter.scala 21:26:@9456.6]
  assign _T_17 = count + 6'h1; // @[Counter.scala 17:24:@9450.4]
  assign newCount = count + 6'h1; // @[Counter.scala 17:24:@9451.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@9456.6]
  assign io_out = count; // @[Counter.scala 25:10:@9459.4]
  assign io_next = count + 6'h1; // @[Counter.scala 26:11:@9460.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[5:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 6'h0;
    end else begin
      if (io_enable) begin
        count <= newCount;
      end
    end
  end
endmodule
module SRAM( // @[:@9496.2]
  input         clock, // @[:@9497.4]
  input         reset, // @[:@9498.4]
  input  [5:0]  io_raddr, // @[:@9499.4]
  input         io_wen, // @[:@9499.4]
  input  [5:0]  io_waddr, // @[:@9499.4]
  input  [63:0] io_wdata_addr, // @[:@9499.4]
  input  [31:0] io_wdata_size, // @[:@9499.4]
  output [63:0] io_rdata_addr, // @[:@9499.4]
  output [31:0] io_rdata_size // @[:@9499.4]
);
  wire [95:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 124:30:@9501.4]
  wire [95:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 124:30:@9501.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 124:30:@9501.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 124:30:@9501.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 124:30:@9501.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 124:30:@9501.4]
  wire [5:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 124:30:@9501.4]
  wire [5:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 124:30:@9501.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 124:30:@9501.4]
  wire [95:0] _T_17; // @[SRAM.scala 130:38:@9515.4]
  wire  _T_20; // @[SRAM.scala 137:49:@9520.4]
  wire  _T_21; // @[SRAM.scala 137:37:@9521.4]
  reg  _T_24; // @[SRAM.scala 137:29:@9522.4]
  reg [31:0] _RAND_0;
  reg [95:0] _T_28; // @[SRAM.scala 138:29:@9525.4]
  reg [95:0] _RAND_1;
  wire [95:0] _T_29; // @[SRAM.scala 139:22:@9527.4]
  SRAMVerilogAWS #(.DWIDTH(96), .WORDS(64), .AWIDTH(6)) SRAMVerilogAWS ( // @[SRAM.scala 124:30:@9501.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_17 = {io_wdata_addr,io_wdata_size}; // @[SRAM.scala 130:38:@9515.4]
  assign _T_20 = io_raddr == io_waddr; // @[SRAM.scala 137:49:@9520.4]
  assign _T_21 = io_wen & _T_20; // @[SRAM.scala 137:37:@9521.4]
  assign _T_29 = _T_24 ? _T_28 : SRAMVerilogAWS_rdata; // @[SRAM.scala 139:22:@9527.4]
  assign io_rdata_addr = _T_29[95:32]; // @[SRAM.scala 139:16:@9536.4]
  assign io_rdata_size = _T_29[31:0]; // @[SRAM.scala 139:16:@9535.4]
  assign SRAMVerilogAWS_wdata = {io_wdata_addr,io_wdata_size}; // @[SRAM.scala 130:20:@9516.4]
  assign SRAMVerilogAWS_backpressure = 1'h1; // @[SRAM.scala 131:27:@9517.4]
  assign SRAMVerilogAWS_wen = io_wen; // @[SRAM.scala 128:18:@9513.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 133:22:@9519.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 132:22:@9518.4]
  assign SRAMVerilogAWS_waddr = io_waddr; // @[SRAM.scala 129:20:@9514.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 127:20:@9512.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 126:18:@9511.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_24 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {3{`RANDOM}};
  _T_28 = _RAND_1[95:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_24 <= 1'h0;
    end else begin
      _T_24 <= _T_21;
    end
    if (reset) begin
      _T_28 <= 96'h0;
    end else begin
      _T_28 <= _T_17;
    end
  end
endmodule
module FIFO( // @[:@9538.2]
  input         clock, // @[:@9539.4]
  input         reset, // @[:@9540.4]
  output        io_in_ready, // @[:@9541.4]
  input         io_in_valid, // @[:@9541.4]
  input  [63:0] io_in_bits_addr, // @[:@9541.4]
  input  [31:0] io_in_bits_size, // @[:@9541.4]
  input         io_out_ready, // @[:@9541.4]
  output        io_out_valid, // @[:@9541.4]
  output [63:0] io_out_bits_addr, // @[:@9541.4]
  output [31:0] io_out_bits_size // @[:@9541.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@9937.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@9937.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@9937.4]
  wire [5:0] enqCounter_io_out; // @[FIFO.scala 34:26:@9937.4]
  wire [5:0] enqCounter_io_next; // @[FIFO.scala 34:26:@9937.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@9947.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@9947.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@9947.4]
  wire [5:0] deqCounter_io_out; // @[FIFO.scala 38:26:@9947.4]
  wire [5:0] deqCounter_io_next; // @[FIFO.scala 38:26:@9947.4]
  wire  SRAM_clock; // @[FIFO.scala 73:19:@9962.4]
  wire  SRAM_reset; // @[FIFO.scala 73:19:@9962.4]
  wire [5:0] SRAM_io_raddr; // @[FIFO.scala 73:19:@9962.4]
  wire  SRAM_io_wen; // @[FIFO.scala 73:19:@9962.4]
  wire [5:0] SRAM_io_waddr; // @[FIFO.scala 73:19:@9962.4]
  wire [63:0] SRAM_io_wdata_addr; // @[FIFO.scala 73:19:@9962.4]
  wire [31:0] SRAM_io_wdata_size; // @[FIFO.scala 73:19:@9962.4]
  wire [63:0] SRAM_io_rdata_addr; // @[FIFO.scala 73:19:@9962.4]
  wire [31:0] SRAM_io_rdata_size; // @[FIFO.scala 73:19:@9962.4]
  wire  writeEn; // @[FIFO.scala 30:29:@9935.4]
  wire  readEn; // @[FIFO.scala 31:29:@9936.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@9957.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@9958.4]
  wire  _T_824; // @[FIFO.scala 45:27:@9959.4]
  wire  empty; // @[FIFO.scala 45:24:@9960.4]
  wire  full; // @[FIFO.scala 46:23:@9961.4]
  wire  _T_827; // @[FIFO.scala 83:17:@9974.4]
  wire  _GEN_0; // @[FIFO.scala 83:29:@9975.4]
  Counter enqCounter ( // @[FIFO.scala 34:26:@9937.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter deqCounter ( // @[FIFO.scala 38:26:@9947.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  SRAM SRAM ( // @[FIFO.scala 73:19:@9962.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata_addr(SRAM_io_wdata_addr),
    .io_wdata_size(SRAM_io_wdata_size),
    .io_rdata_addr(SRAM_io_rdata_addr),
    .io_rdata_size(SRAM_io_rdata_size)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@9935.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@9936.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@9958.4]
  assign _T_824 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@9959.4]
  assign empty = ptrMatch & _T_824; // @[FIFO.scala 45:24:@9960.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@9961.4]
  assign _T_827 = writeEn != readEn; // @[FIFO.scala 83:17:@9974.4]
  assign _GEN_0 = _T_827 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@9975.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@9981.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@9979.4]
  assign io_out_bits_addr = SRAM_io_rdata_addr; // @[FIFO.scala 79:17:@9972.4]
  assign io_out_bits_size = SRAM_io_rdata_size; // @[FIFO.scala 79:17:@9971.4]
  assign enqCounter_clock = clock; // @[:@9938.4]
  assign enqCounter_reset = reset; // @[:@9939.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@9945.4]
  assign deqCounter_clock = clock; // @[:@9948.4]
  assign deqCounter_reset = reset; // @[:@9949.4]
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@9955.4]
  assign SRAM_clock = clock; // @[:@9963.4]
  assign SRAM_reset = reset; // @[:@9964.4]
  assign SRAM_io_raddr = readEn ? deqCounter_io_next : deqCounter_io_out; // @[FIFO.scala 75:16:@9966.4]
  assign SRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 76:14:@9967.4]
  assign SRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 77:16:@9968.4]
  assign SRAM_io_wdata_addr = io_in_bits_addr; // @[FIFO.scala 78:16:@9970.4]
  assign SRAM_io_wdata_size = io_in_bits_size; // @[FIFO.scala 78:16:@9969.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_827) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module Counter_2( // @[:@9983.2]
  input        clock, // @[:@9984.4]
  input        reset, // @[:@9985.4]
  input        io_enable, // @[:@9986.4]
  output [3:0] io_out // @[:@9986.4]
);
  reg [3:0] count; // @[Counter.scala 15:22:@9988.4]
  reg [31:0] _RAND_0;
  wire [4:0] _T_17; // @[Counter.scala 17:24:@9989.4]
  wire [3:0] newCount; // @[Counter.scala 17:24:@9990.4]
  wire [3:0] _GEN_0; // @[Counter.scala 21:26:@9995.6]
  assign _T_17 = count + 4'h1; // @[Counter.scala 17:24:@9989.4]
  assign newCount = count + 4'h1; // @[Counter.scala 17:24:@9990.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@9995.6]
  assign io_out = count; // @[Counter.scala 25:10:@9998.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 4'h0;
    end else begin
      if (io_enable) begin
        count <= newCount;
      end
    end
  end
endmodule
module Counter_4( // @[:@10019.2]
  input        clock, // @[:@10020.4]
  input        reset, // @[:@10021.4]
  input        io_reset, // @[:@10022.4]
  input        io_enable, // @[:@10022.4]
  input  [1:0] io_stride, // @[:@10022.4]
  output [1:0] io_out, // @[:@10022.4]
  output [1:0] io_next // @[:@10022.4]
);
  reg [1:0] count; // @[Counter.scala 15:22:@10024.4]
  reg [31:0] _RAND_0;
  wire [2:0] _T_17; // @[Counter.scala 17:24:@10025.4]
  wire [1:0] newCount; // @[Counter.scala 17:24:@10026.4]
  wire [1:0] _GEN_0; // @[Counter.scala 21:26:@10031.6]
  wire [1:0] _GEN_1; // @[Counter.scala 19:18:@10027.4]
  assign _T_17 = count + io_stride; // @[Counter.scala 17:24:@10025.4]
  assign newCount = count + io_stride; // @[Counter.scala 17:24:@10026.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@10031.6]
  assign _GEN_1 = io_reset ? 2'h0 : _GEN_0; // @[Counter.scala 19:18:@10027.4]
  assign io_out = count; // @[Counter.scala 25:10:@10034.4]
  assign io_next = count + io_stride; // @[Counter.scala 26:11:@10035.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 2'h0;
    end else begin
      if (io_reset) begin
        count <= 2'h0;
      end else begin
        if (io_enable) begin
          count <= newCount;
        end
      end
    end
  end
endmodule
module SRAM_1( // @[:@10071.2]
  input         clock, // @[:@10072.4]
  input         reset, // @[:@10073.4]
  input  [1:0]  io_raddr, // @[:@10074.4]
  input         io_wen, // @[:@10074.4]
  input  [1:0]  io_waddr, // @[:@10074.4]
  input  [31:0] io_wdata, // @[:@10074.4]
  output [31:0] io_rdata, // @[:@10074.4]
  input         io_backpressure // @[:@10074.4]
);
  wire [31:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 124:30:@10076.4]
  wire [31:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 124:30:@10076.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 124:30:@10076.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 124:30:@10076.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 124:30:@10076.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 124:30:@10076.4]
  wire [1:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 124:30:@10076.4]
  wire [1:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 124:30:@10076.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 124:30:@10076.4]
  wire  _T_19; // @[SRAM.scala 137:49:@10094.4]
  wire  _T_20; // @[SRAM.scala 137:37:@10095.4]
  reg  _T_23; // @[SRAM.scala 137:29:@10096.4]
  reg [31:0] _RAND_0;
  reg [31:0] _T_26; // @[SRAM.scala 138:29:@10098.4]
  reg [31:0] _RAND_1;
  SRAMVerilogAWS #(.DWIDTH(32), .WORDS(4), .AWIDTH(2)) SRAMVerilogAWS ( // @[SRAM.scala 124:30:@10076.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_19 = io_raddr == io_waddr; // @[SRAM.scala 137:49:@10094.4]
  assign _T_20 = io_wen & _T_19; // @[SRAM.scala 137:37:@10095.4]
  assign io_rdata = _T_23 ? _T_26 : SRAMVerilogAWS_rdata; // @[SRAM.scala 139:16:@10103.4]
  assign SRAMVerilogAWS_wdata = io_wdata; // @[SRAM.scala 130:20:@10090.4]
  assign SRAMVerilogAWS_backpressure = io_backpressure; // @[SRAM.scala 131:27:@10091.4]
  assign SRAMVerilogAWS_wen = io_wen; // @[SRAM.scala 128:18:@10088.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 133:22:@10093.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 132:22:@10092.4]
  assign SRAMVerilogAWS_waddr = io_waddr; // @[SRAM.scala 129:20:@10089.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 127:20:@10087.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 126:18:@10086.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_23 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_26 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_23 <= 1'h0;
    end else begin
      _T_23 <= _T_20;
    end
    if (reset) begin
      _T_26 <= 32'h0;
    end else begin
      _T_26 <= io_wdata;
    end
  end
endmodule
module FIFO_1( // @[:@10105.2]
  input         clock, // @[:@10106.4]
  input         reset, // @[:@10107.4]
  output        io_in_ready, // @[:@10108.4]
  input         io_in_valid, // @[:@10108.4]
  input  [31:0] io_in_bits, // @[:@10108.4]
  input         io_out_ready, // @[:@10108.4]
  output        io_out_valid, // @[:@10108.4]
  output [31:0] io_out_bits // @[:@10108.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@10134.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@10134.4]
  wire  enqCounter_io_reset; // @[FIFO.scala 34:26:@10134.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@10134.4]
  wire [1:0] enqCounter_io_stride; // @[FIFO.scala 34:26:@10134.4]
  wire [1:0] enqCounter_io_out; // @[FIFO.scala 34:26:@10134.4]
  wire [1:0] enqCounter_io_next; // @[FIFO.scala 34:26:@10134.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@10144.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@10144.4]
  wire  deqCounter_io_reset; // @[FIFO.scala 38:26:@10144.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@10144.4]
  wire [1:0] deqCounter_io_stride; // @[FIFO.scala 38:26:@10144.4]
  wire [1:0] deqCounter_io_out; // @[FIFO.scala 38:26:@10144.4]
  wire [1:0] deqCounter_io_next; // @[FIFO.scala 38:26:@10144.4]
  wire  SRAM_clock; // @[FIFO.scala 73:19:@10159.4]
  wire  SRAM_reset; // @[FIFO.scala 73:19:@10159.4]
  wire [1:0] SRAM_io_raddr; // @[FIFO.scala 73:19:@10159.4]
  wire  SRAM_io_wen; // @[FIFO.scala 73:19:@10159.4]
  wire [1:0] SRAM_io_waddr; // @[FIFO.scala 73:19:@10159.4]
  wire [31:0] SRAM_io_wdata; // @[FIFO.scala 73:19:@10159.4]
  wire [31:0] SRAM_io_rdata; // @[FIFO.scala 73:19:@10159.4]
  wire  SRAM_io_backpressure; // @[FIFO.scala 73:19:@10159.4]
  wire  writeEn; // @[FIFO.scala 30:29:@10132.4]
  wire  readEn; // @[FIFO.scala 31:29:@10133.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@10154.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@10155.4]
  wire  _T_104; // @[FIFO.scala 45:27:@10156.4]
  wire  empty; // @[FIFO.scala 45:24:@10157.4]
  wire  full; // @[FIFO.scala 46:23:@10158.4]
  wire  _T_107; // @[FIFO.scala 83:17:@10169.4]
  wire  _GEN_0; // @[FIFO.scala 83:29:@10170.4]
  Counter_4 enqCounter ( // @[FIFO.scala 34:26:@10134.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_reset(enqCounter_io_reset),
    .io_enable(enqCounter_io_enable),
    .io_stride(enqCounter_io_stride),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter_4 deqCounter ( // @[FIFO.scala 38:26:@10144.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_reset(deqCounter_io_reset),
    .io_enable(deqCounter_io_enable),
    .io_stride(deqCounter_io_stride),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  SRAM_1 SRAM ( // @[FIFO.scala 73:19:@10159.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata(SRAM_io_wdata),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@10132.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@10133.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@10155.4]
  assign _T_104 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@10156.4]
  assign empty = ptrMatch & _T_104; // @[FIFO.scala 45:24:@10157.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@10158.4]
  assign _T_107 = writeEn != readEn; // @[FIFO.scala 83:17:@10169.4]
  assign _GEN_0 = _T_107 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@10170.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@10176.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@10174.4]
  assign io_out_bits = SRAM_io_rdata; // @[FIFO.scala 79:17:@10167.4]
  assign enqCounter_clock = clock; // @[:@10135.4]
  assign enqCounter_reset = reset; // @[:@10136.4]
  assign enqCounter_io_reset = 1'h0;
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@10142.4]
  assign enqCounter_io_stride = 2'h1; // @[FIFO.scala 37:24:@10143.4]
  assign deqCounter_clock = clock; // @[:@10145.4]
  assign deqCounter_reset = reset; // @[:@10146.4]
  assign deqCounter_io_reset = 1'h0;
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@10152.4]
  assign deqCounter_io_stride = 2'h1; // @[FIFO.scala 41:24:@10153.4]
  assign SRAM_clock = clock; // @[:@10160.4]
  assign SRAM_reset = reset; // @[:@10161.4]
  assign SRAM_io_raddr = readEn ? deqCounter_io_next : deqCounter_io_out; // @[FIFO.scala 75:16:@10163.4]
  assign SRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 76:14:@10164.4]
  assign SRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 77:16:@10165.4]
  assign SRAM_io_wdata = io_in_bits; // @[FIFO.scala 78:16:@10166.4]
  assign SRAM_io_backpressure = 1'h1; // @[FIFO.scala 80:23:@10168.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_107) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module FIFOVec( // @[:@12563.2]
  input         clock, // @[:@12564.4]
  input         reset, // @[:@12565.4]
  output        io_in_ready, // @[:@12566.4]
  input         io_in_valid, // @[:@12566.4]
  input  [31:0] io_in_bits_0, // @[:@12566.4]
  input  [31:0] io_in_bits_1, // @[:@12566.4]
  input  [31:0] io_in_bits_2, // @[:@12566.4]
  input  [31:0] io_in_bits_3, // @[:@12566.4]
  input  [31:0] io_in_bits_4, // @[:@12566.4]
  input  [31:0] io_in_bits_5, // @[:@12566.4]
  input  [31:0] io_in_bits_6, // @[:@12566.4]
  input  [31:0] io_in_bits_7, // @[:@12566.4]
  input  [31:0] io_in_bits_8, // @[:@12566.4]
  input  [31:0] io_in_bits_9, // @[:@12566.4]
  input  [31:0] io_in_bits_10, // @[:@12566.4]
  input  [31:0] io_in_bits_11, // @[:@12566.4]
  input  [31:0] io_in_bits_12, // @[:@12566.4]
  input  [31:0] io_in_bits_13, // @[:@12566.4]
  input  [31:0] io_in_bits_14, // @[:@12566.4]
  input  [31:0] io_in_bits_15, // @[:@12566.4]
  input         io_out_ready, // @[:@12566.4]
  output        io_out_valid, // @[:@12566.4]
  output [31:0] io_out_bits_0 // @[:@12566.4]
);
  wire  enqCounter_clock; // @[FIFOVec.scala 24:26:@12570.4]
  wire  enqCounter_reset; // @[FIFOVec.scala 24:26:@12570.4]
  wire  enqCounter_io_enable; // @[FIFOVec.scala 24:26:@12570.4]
  wire [3:0] enqCounter_io_out; // @[FIFOVec.scala 24:26:@12570.4]
  wire  deqCounter_clock; // @[FIFOVec.scala 28:26:@12581.4]
  wire  deqCounter_reset; // @[FIFOVec.scala 28:26:@12581.4]
  wire  deqCounter_io_enable; // @[FIFOVec.scala 28:26:@12581.4]
  wire [3:0] deqCounter_io_out; // @[FIFOVec.scala 28:26:@12581.4]
  wire  fifos_0_clock; // @[FIFOVec.scala 40:19:@12594.4]
  wire  fifos_0_reset; // @[FIFOVec.scala 40:19:@12594.4]
  wire  fifos_0_io_in_ready; // @[FIFOVec.scala 40:19:@12594.4]
  wire  fifos_0_io_in_valid; // @[FIFOVec.scala 40:19:@12594.4]
  wire [31:0] fifos_0_io_in_bits; // @[FIFOVec.scala 40:19:@12594.4]
  wire  fifos_0_io_out_ready; // @[FIFOVec.scala 40:19:@12594.4]
  wire  fifos_0_io_out_valid; // @[FIFOVec.scala 40:19:@12594.4]
  wire [31:0] fifos_0_io_out_bits; // @[FIFOVec.scala 40:19:@12594.4]
  wire  fifos_1_clock; // @[FIFOVec.scala 40:19:@12629.4]
  wire  fifos_1_reset; // @[FIFOVec.scala 40:19:@12629.4]
  wire  fifos_1_io_in_ready; // @[FIFOVec.scala 40:19:@12629.4]
  wire  fifos_1_io_in_valid; // @[FIFOVec.scala 40:19:@12629.4]
  wire [31:0] fifos_1_io_in_bits; // @[FIFOVec.scala 40:19:@12629.4]
  wire  fifos_1_io_out_ready; // @[FIFOVec.scala 40:19:@12629.4]
  wire  fifos_1_io_out_valid; // @[FIFOVec.scala 40:19:@12629.4]
  wire [31:0] fifos_1_io_out_bits; // @[FIFOVec.scala 40:19:@12629.4]
  wire  fifos_2_clock; // @[FIFOVec.scala 40:19:@12664.4]
  wire  fifos_2_reset; // @[FIFOVec.scala 40:19:@12664.4]
  wire  fifos_2_io_in_ready; // @[FIFOVec.scala 40:19:@12664.4]
  wire  fifos_2_io_in_valid; // @[FIFOVec.scala 40:19:@12664.4]
  wire [31:0] fifos_2_io_in_bits; // @[FIFOVec.scala 40:19:@12664.4]
  wire  fifos_2_io_out_ready; // @[FIFOVec.scala 40:19:@12664.4]
  wire  fifos_2_io_out_valid; // @[FIFOVec.scala 40:19:@12664.4]
  wire [31:0] fifos_2_io_out_bits; // @[FIFOVec.scala 40:19:@12664.4]
  wire  fifos_3_clock; // @[FIFOVec.scala 40:19:@12699.4]
  wire  fifos_3_reset; // @[FIFOVec.scala 40:19:@12699.4]
  wire  fifos_3_io_in_ready; // @[FIFOVec.scala 40:19:@12699.4]
  wire  fifos_3_io_in_valid; // @[FIFOVec.scala 40:19:@12699.4]
  wire [31:0] fifos_3_io_in_bits; // @[FIFOVec.scala 40:19:@12699.4]
  wire  fifos_3_io_out_ready; // @[FIFOVec.scala 40:19:@12699.4]
  wire  fifos_3_io_out_valid; // @[FIFOVec.scala 40:19:@12699.4]
  wire [31:0] fifos_3_io_out_bits; // @[FIFOVec.scala 40:19:@12699.4]
  wire  fifos_4_clock; // @[FIFOVec.scala 40:19:@12734.4]
  wire  fifos_4_reset; // @[FIFOVec.scala 40:19:@12734.4]
  wire  fifos_4_io_in_ready; // @[FIFOVec.scala 40:19:@12734.4]
  wire  fifos_4_io_in_valid; // @[FIFOVec.scala 40:19:@12734.4]
  wire [31:0] fifos_4_io_in_bits; // @[FIFOVec.scala 40:19:@12734.4]
  wire  fifos_4_io_out_ready; // @[FIFOVec.scala 40:19:@12734.4]
  wire  fifos_4_io_out_valid; // @[FIFOVec.scala 40:19:@12734.4]
  wire [31:0] fifos_4_io_out_bits; // @[FIFOVec.scala 40:19:@12734.4]
  wire  fifos_5_clock; // @[FIFOVec.scala 40:19:@12769.4]
  wire  fifos_5_reset; // @[FIFOVec.scala 40:19:@12769.4]
  wire  fifos_5_io_in_ready; // @[FIFOVec.scala 40:19:@12769.4]
  wire  fifos_5_io_in_valid; // @[FIFOVec.scala 40:19:@12769.4]
  wire [31:0] fifos_5_io_in_bits; // @[FIFOVec.scala 40:19:@12769.4]
  wire  fifos_5_io_out_ready; // @[FIFOVec.scala 40:19:@12769.4]
  wire  fifos_5_io_out_valid; // @[FIFOVec.scala 40:19:@12769.4]
  wire [31:0] fifos_5_io_out_bits; // @[FIFOVec.scala 40:19:@12769.4]
  wire  fifos_6_clock; // @[FIFOVec.scala 40:19:@12804.4]
  wire  fifos_6_reset; // @[FIFOVec.scala 40:19:@12804.4]
  wire  fifos_6_io_in_ready; // @[FIFOVec.scala 40:19:@12804.4]
  wire  fifos_6_io_in_valid; // @[FIFOVec.scala 40:19:@12804.4]
  wire [31:0] fifos_6_io_in_bits; // @[FIFOVec.scala 40:19:@12804.4]
  wire  fifos_6_io_out_ready; // @[FIFOVec.scala 40:19:@12804.4]
  wire  fifos_6_io_out_valid; // @[FIFOVec.scala 40:19:@12804.4]
  wire [31:0] fifos_6_io_out_bits; // @[FIFOVec.scala 40:19:@12804.4]
  wire  fifos_7_clock; // @[FIFOVec.scala 40:19:@12839.4]
  wire  fifos_7_reset; // @[FIFOVec.scala 40:19:@12839.4]
  wire  fifos_7_io_in_ready; // @[FIFOVec.scala 40:19:@12839.4]
  wire  fifos_7_io_in_valid; // @[FIFOVec.scala 40:19:@12839.4]
  wire [31:0] fifos_7_io_in_bits; // @[FIFOVec.scala 40:19:@12839.4]
  wire  fifos_7_io_out_ready; // @[FIFOVec.scala 40:19:@12839.4]
  wire  fifos_7_io_out_valid; // @[FIFOVec.scala 40:19:@12839.4]
  wire [31:0] fifos_7_io_out_bits; // @[FIFOVec.scala 40:19:@12839.4]
  wire  fifos_8_clock; // @[FIFOVec.scala 40:19:@12874.4]
  wire  fifos_8_reset; // @[FIFOVec.scala 40:19:@12874.4]
  wire  fifos_8_io_in_ready; // @[FIFOVec.scala 40:19:@12874.4]
  wire  fifos_8_io_in_valid; // @[FIFOVec.scala 40:19:@12874.4]
  wire [31:0] fifos_8_io_in_bits; // @[FIFOVec.scala 40:19:@12874.4]
  wire  fifos_8_io_out_ready; // @[FIFOVec.scala 40:19:@12874.4]
  wire  fifos_8_io_out_valid; // @[FIFOVec.scala 40:19:@12874.4]
  wire [31:0] fifos_8_io_out_bits; // @[FIFOVec.scala 40:19:@12874.4]
  wire  fifos_9_clock; // @[FIFOVec.scala 40:19:@12909.4]
  wire  fifos_9_reset; // @[FIFOVec.scala 40:19:@12909.4]
  wire  fifos_9_io_in_ready; // @[FIFOVec.scala 40:19:@12909.4]
  wire  fifos_9_io_in_valid; // @[FIFOVec.scala 40:19:@12909.4]
  wire [31:0] fifos_9_io_in_bits; // @[FIFOVec.scala 40:19:@12909.4]
  wire  fifos_9_io_out_ready; // @[FIFOVec.scala 40:19:@12909.4]
  wire  fifos_9_io_out_valid; // @[FIFOVec.scala 40:19:@12909.4]
  wire [31:0] fifos_9_io_out_bits; // @[FIFOVec.scala 40:19:@12909.4]
  wire  fifos_10_clock; // @[FIFOVec.scala 40:19:@12944.4]
  wire  fifos_10_reset; // @[FIFOVec.scala 40:19:@12944.4]
  wire  fifos_10_io_in_ready; // @[FIFOVec.scala 40:19:@12944.4]
  wire  fifos_10_io_in_valid; // @[FIFOVec.scala 40:19:@12944.4]
  wire [31:0] fifos_10_io_in_bits; // @[FIFOVec.scala 40:19:@12944.4]
  wire  fifos_10_io_out_ready; // @[FIFOVec.scala 40:19:@12944.4]
  wire  fifos_10_io_out_valid; // @[FIFOVec.scala 40:19:@12944.4]
  wire [31:0] fifos_10_io_out_bits; // @[FIFOVec.scala 40:19:@12944.4]
  wire  fifos_11_clock; // @[FIFOVec.scala 40:19:@12979.4]
  wire  fifos_11_reset; // @[FIFOVec.scala 40:19:@12979.4]
  wire  fifos_11_io_in_ready; // @[FIFOVec.scala 40:19:@12979.4]
  wire  fifos_11_io_in_valid; // @[FIFOVec.scala 40:19:@12979.4]
  wire [31:0] fifos_11_io_in_bits; // @[FIFOVec.scala 40:19:@12979.4]
  wire  fifos_11_io_out_ready; // @[FIFOVec.scala 40:19:@12979.4]
  wire  fifos_11_io_out_valid; // @[FIFOVec.scala 40:19:@12979.4]
  wire [31:0] fifos_11_io_out_bits; // @[FIFOVec.scala 40:19:@12979.4]
  wire  fifos_12_clock; // @[FIFOVec.scala 40:19:@13014.4]
  wire  fifos_12_reset; // @[FIFOVec.scala 40:19:@13014.4]
  wire  fifos_12_io_in_ready; // @[FIFOVec.scala 40:19:@13014.4]
  wire  fifos_12_io_in_valid; // @[FIFOVec.scala 40:19:@13014.4]
  wire [31:0] fifos_12_io_in_bits; // @[FIFOVec.scala 40:19:@13014.4]
  wire  fifos_12_io_out_ready; // @[FIFOVec.scala 40:19:@13014.4]
  wire  fifos_12_io_out_valid; // @[FIFOVec.scala 40:19:@13014.4]
  wire [31:0] fifos_12_io_out_bits; // @[FIFOVec.scala 40:19:@13014.4]
  wire  fifos_13_clock; // @[FIFOVec.scala 40:19:@13049.4]
  wire  fifos_13_reset; // @[FIFOVec.scala 40:19:@13049.4]
  wire  fifos_13_io_in_ready; // @[FIFOVec.scala 40:19:@13049.4]
  wire  fifos_13_io_in_valid; // @[FIFOVec.scala 40:19:@13049.4]
  wire [31:0] fifos_13_io_in_bits; // @[FIFOVec.scala 40:19:@13049.4]
  wire  fifos_13_io_out_ready; // @[FIFOVec.scala 40:19:@13049.4]
  wire  fifos_13_io_out_valid; // @[FIFOVec.scala 40:19:@13049.4]
  wire [31:0] fifos_13_io_out_bits; // @[FIFOVec.scala 40:19:@13049.4]
  wire  fifos_14_clock; // @[FIFOVec.scala 40:19:@13084.4]
  wire  fifos_14_reset; // @[FIFOVec.scala 40:19:@13084.4]
  wire  fifos_14_io_in_ready; // @[FIFOVec.scala 40:19:@13084.4]
  wire  fifos_14_io_in_valid; // @[FIFOVec.scala 40:19:@13084.4]
  wire [31:0] fifos_14_io_in_bits; // @[FIFOVec.scala 40:19:@13084.4]
  wire  fifos_14_io_out_ready; // @[FIFOVec.scala 40:19:@13084.4]
  wire  fifos_14_io_out_valid; // @[FIFOVec.scala 40:19:@13084.4]
  wire [31:0] fifos_14_io_out_bits; // @[FIFOVec.scala 40:19:@13084.4]
  wire  fifos_15_clock; // @[FIFOVec.scala 40:19:@13119.4]
  wire  fifos_15_reset; // @[FIFOVec.scala 40:19:@13119.4]
  wire  fifos_15_io_in_ready; // @[FIFOVec.scala 40:19:@13119.4]
  wire  fifos_15_io_in_valid; // @[FIFOVec.scala 40:19:@13119.4]
  wire [31:0] fifos_15_io_in_bits; // @[FIFOVec.scala 40:19:@13119.4]
  wire  fifos_15_io_out_ready; // @[FIFOVec.scala 40:19:@13119.4]
  wire  fifos_15_io_out_valid; // @[FIFOVec.scala 40:19:@13119.4]
  wire [31:0] fifos_15_io_out_bits; // @[FIFOVec.scala 40:19:@13119.4]
  wire  readEn; // @[FIFOVec.scala 20:29:@12568.4]
  wire [15:0] deqDecoder; // @[OneHot.scala 45:35:@12593.4]
  wire  _T_154; // @[FIFOVec.scala 44:50:@12625.4]
  wire  _T_163; // @[FIFOVec.scala 44:50:@12660.4]
  wire  _T_172; // @[FIFOVec.scala 44:50:@12695.4]
  wire  _T_181; // @[FIFOVec.scala 44:50:@12730.4]
  wire  _T_190; // @[FIFOVec.scala 44:50:@12765.4]
  wire  _T_199; // @[FIFOVec.scala 44:50:@12800.4]
  wire  _T_208; // @[FIFOVec.scala 44:50:@12835.4]
  wire  _T_217; // @[FIFOVec.scala 44:50:@12870.4]
  wire  _T_226; // @[FIFOVec.scala 44:50:@12905.4]
  wire  _T_235; // @[FIFOVec.scala 44:50:@12940.4]
  wire  _T_244; // @[FIFOVec.scala 44:50:@12975.4]
  wire  _T_253; // @[FIFOVec.scala 44:50:@13010.4]
  wire  _T_262; // @[FIFOVec.scala 44:50:@13045.4]
  wire  _T_271; // @[FIFOVec.scala 44:50:@13080.4]
  wire  _T_280; // @[FIFOVec.scala 44:50:@13115.4]
  wire  _T_289; // @[FIFOVec.scala 44:50:@13150.4]
  wire  _T_316; // @[FIFOVec.scala 49:90:@13171.4]
  wire  _T_317; // @[FIFOVec.scala 49:90:@13172.4]
  wire  _T_318; // @[FIFOVec.scala 49:90:@13173.4]
  wire  _T_319; // @[FIFOVec.scala 49:90:@13174.4]
  wire  _T_320; // @[FIFOVec.scala 49:90:@13175.4]
  wire  _T_321; // @[FIFOVec.scala 49:90:@13176.4]
  wire  _T_322; // @[FIFOVec.scala 49:90:@13177.4]
  wire  _T_323; // @[FIFOVec.scala 49:90:@13178.4]
  wire  _T_324; // @[FIFOVec.scala 49:90:@13179.4]
  wire  _T_325; // @[FIFOVec.scala 49:90:@13180.4]
  wire  _T_326; // @[FIFOVec.scala 49:90:@13181.4]
  wire  _T_327; // @[FIFOVec.scala 49:90:@13182.4]
  wire  _T_328; // @[FIFOVec.scala 49:90:@13183.4]
  wire  _T_329; // @[FIFOVec.scala 49:90:@13184.4]
  wire  _T_335_0; // @[FIFOVec.scala 51:43:@13188.4 FIFOVec.scala 51:43:@13189.4]
  wire  _T_335_1; // @[FIFOVec.scala 51:43:@13188.4 FIFOVec.scala 51:43:@13190.4]
  wire  _GEN_17; // @[FIFOVec.scala 51:22:@13220.4]
  wire  _T_335_2; // @[FIFOVec.scala 51:43:@13188.4 FIFOVec.scala 51:43:@13191.4]
  wire  _GEN_18; // @[FIFOVec.scala 51:22:@13220.4]
  wire  _T_335_3; // @[FIFOVec.scala 51:43:@13188.4 FIFOVec.scala 51:43:@13192.4]
  wire  _GEN_19; // @[FIFOVec.scala 51:22:@13220.4]
  wire  _T_335_4; // @[FIFOVec.scala 51:43:@13188.4 FIFOVec.scala 51:43:@13193.4]
  wire  _GEN_20; // @[FIFOVec.scala 51:22:@13220.4]
  wire  _T_335_5; // @[FIFOVec.scala 51:43:@13188.4 FIFOVec.scala 51:43:@13194.4]
  wire  _GEN_21; // @[FIFOVec.scala 51:22:@13220.4]
  wire  _T_335_6; // @[FIFOVec.scala 51:43:@13188.4 FIFOVec.scala 51:43:@13195.4]
  wire  _GEN_22; // @[FIFOVec.scala 51:22:@13220.4]
  wire  _T_335_7; // @[FIFOVec.scala 51:43:@13188.4 FIFOVec.scala 51:43:@13196.4]
  wire  _GEN_23; // @[FIFOVec.scala 51:22:@13220.4]
  wire  _T_335_8; // @[FIFOVec.scala 51:43:@13188.4 FIFOVec.scala 51:43:@13197.4]
  wire  _GEN_24; // @[FIFOVec.scala 51:22:@13220.4]
  wire  _T_335_9; // @[FIFOVec.scala 51:43:@13188.4 FIFOVec.scala 51:43:@13198.4]
  wire  _GEN_25; // @[FIFOVec.scala 51:22:@13220.4]
  wire  _T_335_10; // @[FIFOVec.scala 51:43:@13188.4 FIFOVec.scala 51:43:@13199.4]
  wire  _GEN_26; // @[FIFOVec.scala 51:22:@13220.4]
  wire  _T_335_11; // @[FIFOVec.scala 51:43:@13188.4 FIFOVec.scala 51:43:@13200.4]
  wire  _GEN_27; // @[FIFOVec.scala 51:22:@13220.4]
  wire  _T_335_12; // @[FIFOVec.scala 51:43:@13188.4 FIFOVec.scala 51:43:@13201.4]
  wire  _GEN_28; // @[FIFOVec.scala 51:22:@13220.4]
  wire  _T_335_13; // @[FIFOVec.scala 51:43:@13188.4 FIFOVec.scala 51:43:@13202.4]
  wire  _GEN_29; // @[FIFOVec.scala 51:22:@13220.4]
  wire  _T_335_14; // @[FIFOVec.scala 51:43:@13188.4 FIFOVec.scala 51:43:@13203.4]
  wire  _GEN_30; // @[FIFOVec.scala 51:22:@13220.4]
  wire  _T_335_15; // @[FIFOVec.scala 51:43:@13188.4 FIFOVec.scala 51:43:@13204.4]
  wire [31:0] _T_374_0; // @[FIFOVec.scala 53:65:@13222.4 FIFOVec.scala 53:65:@13223.4]
  wire [31:0] _T_374_1; // @[FIFOVec.scala 53:65:@13222.4 FIFOVec.scala 53:65:@13224.4]
  wire [31:0] _GEN_33; // @[FIFOVec.scala 53:42:@13495.4]
  wire [31:0] _T_374_2; // @[FIFOVec.scala 53:65:@13222.4 FIFOVec.scala 53:65:@13225.4]
  wire [31:0] _GEN_34; // @[FIFOVec.scala 53:42:@13495.4]
  wire [31:0] _T_374_3; // @[FIFOVec.scala 53:65:@13222.4 FIFOVec.scala 53:65:@13226.4]
  wire [31:0] _GEN_35; // @[FIFOVec.scala 53:42:@13495.4]
  wire [31:0] _T_374_4; // @[FIFOVec.scala 53:65:@13222.4 FIFOVec.scala 53:65:@13227.4]
  wire [31:0] _GEN_36; // @[FIFOVec.scala 53:42:@13495.4]
  wire [31:0] _T_374_5; // @[FIFOVec.scala 53:65:@13222.4 FIFOVec.scala 53:65:@13228.4]
  wire [31:0] _GEN_37; // @[FIFOVec.scala 53:42:@13495.4]
  wire [31:0] _T_374_6; // @[FIFOVec.scala 53:65:@13222.4 FIFOVec.scala 53:65:@13229.4]
  wire [31:0] _GEN_38; // @[FIFOVec.scala 53:42:@13495.4]
  wire [31:0] _T_374_7; // @[FIFOVec.scala 53:65:@13222.4 FIFOVec.scala 53:65:@13230.4]
  wire [31:0] _GEN_39; // @[FIFOVec.scala 53:42:@13495.4]
  wire [31:0] _T_374_8; // @[FIFOVec.scala 53:65:@13222.4 FIFOVec.scala 53:65:@13231.4]
  wire [31:0] _GEN_40; // @[FIFOVec.scala 53:42:@13495.4]
  wire [31:0] _T_374_9; // @[FIFOVec.scala 53:65:@13222.4 FIFOVec.scala 53:65:@13232.4]
  wire [31:0] _GEN_41; // @[FIFOVec.scala 53:42:@13495.4]
  wire [31:0] _T_374_10; // @[FIFOVec.scala 53:65:@13222.4 FIFOVec.scala 53:65:@13233.4]
  wire [31:0] _GEN_42; // @[FIFOVec.scala 53:42:@13495.4]
  wire [31:0] _T_374_11; // @[FIFOVec.scala 53:65:@13222.4 FIFOVec.scala 53:65:@13234.4]
  wire [31:0] _GEN_43; // @[FIFOVec.scala 53:42:@13495.4]
  wire [31:0] _T_374_12; // @[FIFOVec.scala 53:65:@13222.4 FIFOVec.scala 53:65:@13235.4]
  wire [31:0] _GEN_44; // @[FIFOVec.scala 53:42:@13495.4]
  wire [31:0] _T_374_13; // @[FIFOVec.scala 53:65:@13222.4 FIFOVec.scala 53:65:@13236.4]
  wire [31:0] _GEN_45; // @[FIFOVec.scala 53:42:@13495.4]
  wire [31:0] _T_374_14; // @[FIFOVec.scala 53:65:@13222.4 FIFOVec.scala 53:65:@13237.4]
  wire [31:0] _GEN_46; // @[FIFOVec.scala 53:42:@13495.4]
  wire [31:0] _T_374_15; // @[FIFOVec.scala 53:65:@13222.4 FIFOVec.scala 53:65:@13238.4]
  Counter_2 enqCounter ( // @[FIFOVec.scala 24:26:@12570.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out)
  );
  Counter_2 deqCounter ( // @[FIFOVec.scala 28:26:@12581.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out)
  );
  FIFO_1 fifos_0 ( // @[FIFOVec.scala 40:19:@12594.4]
    .clock(fifos_0_clock),
    .reset(fifos_0_reset),
    .io_in_ready(fifos_0_io_in_ready),
    .io_in_valid(fifos_0_io_in_valid),
    .io_in_bits(fifos_0_io_in_bits),
    .io_out_ready(fifos_0_io_out_ready),
    .io_out_valid(fifos_0_io_out_valid),
    .io_out_bits(fifos_0_io_out_bits)
  );
  FIFO_1 fifos_1 ( // @[FIFOVec.scala 40:19:@12629.4]
    .clock(fifos_1_clock),
    .reset(fifos_1_reset),
    .io_in_ready(fifos_1_io_in_ready),
    .io_in_valid(fifos_1_io_in_valid),
    .io_in_bits(fifos_1_io_in_bits),
    .io_out_ready(fifos_1_io_out_ready),
    .io_out_valid(fifos_1_io_out_valid),
    .io_out_bits(fifos_1_io_out_bits)
  );
  FIFO_1 fifos_2 ( // @[FIFOVec.scala 40:19:@12664.4]
    .clock(fifos_2_clock),
    .reset(fifos_2_reset),
    .io_in_ready(fifos_2_io_in_ready),
    .io_in_valid(fifos_2_io_in_valid),
    .io_in_bits(fifos_2_io_in_bits),
    .io_out_ready(fifos_2_io_out_ready),
    .io_out_valid(fifos_2_io_out_valid),
    .io_out_bits(fifos_2_io_out_bits)
  );
  FIFO_1 fifos_3 ( // @[FIFOVec.scala 40:19:@12699.4]
    .clock(fifos_3_clock),
    .reset(fifos_3_reset),
    .io_in_ready(fifos_3_io_in_ready),
    .io_in_valid(fifos_3_io_in_valid),
    .io_in_bits(fifos_3_io_in_bits),
    .io_out_ready(fifos_3_io_out_ready),
    .io_out_valid(fifos_3_io_out_valid),
    .io_out_bits(fifos_3_io_out_bits)
  );
  FIFO_1 fifos_4 ( // @[FIFOVec.scala 40:19:@12734.4]
    .clock(fifos_4_clock),
    .reset(fifos_4_reset),
    .io_in_ready(fifos_4_io_in_ready),
    .io_in_valid(fifos_4_io_in_valid),
    .io_in_bits(fifos_4_io_in_bits),
    .io_out_ready(fifos_4_io_out_ready),
    .io_out_valid(fifos_4_io_out_valid),
    .io_out_bits(fifos_4_io_out_bits)
  );
  FIFO_1 fifos_5 ( // @[FIFOVec.scala 40:19:@12769.4]
    .clock(fifos_5_clock),
    .reset(fifos_5_reset),
    .io_in_ready(fifos_5_io_in_ready),
    .io_in_valid(fifos_5_io_in_valid),
    .io_in_bits(fifos_5_io_in_bits),
    .io_out_ready(fifos_5_io_out_ready),
    .io_out_valid(fifos_5_io_out_valid),
    .io_out_bits(fifos_5_io_out_bits)
  );
  FIFO_1 fifos_6 ( // @[FIFOVec.scala 40:19:@12804.4]
    .clock(fifos_6_clock),
    .reset(fifos_6_reset),
    .io_in_ready(fifos_6_io_in_ready),
    .io_in_valid(fifos_6_io_in_valid),
    .io_in_bits(fifos_6_io_in_bits),
    .io_out_ready(fifos_6_io_out_ready),
    .io_out_valid(fifos_6_io_out_valid),
    .io_out_bits(fifos_6_io_out_bits)
  );
  FIFO_1 fifos_7 ( // @[FIFOVec.scala 40:19:@12839.4]
    .clock(fifos_7_clock),
    .reset(fifos_7_reset),
    .io_in_ready(fifos_7_io_in_ready),
    .io_in_valid(fifos_7_io_in_valid),
    .io_in_bits(fifos_7_io_in_bits),
    .io_out_ready(fifos_7_io_out_ready),
    .io_out_valid(fifos_7_io_out_valid),
    .io_out_bits(fifos_7_io_out_bits)
  );
  FIFO_1 fifos_8 ( // @[FIFOVec.scala 40:19:@12874.4]
    .clock(fifos_8_clock),
    .reset(fifos_8_reset),
    .io_in_ready(fifos_8_io_in_ready),
    .io_in_valid(fifos_8_io_in_valid),
    .io_in_bits(fifos_8_io_in_bits),
    .io_out_ready(fifos_8_io_out_ready),
    .io_out_valid(fifos_8_io_out_valid),
    .io_out_bits(fifos_8_io_out_bits)
  );
  FIFO_1 fifos_9 ( // @[FIFOVec.scala 40:19:@12909.4]
    .clock(fifos_9_clock),
    .reset(fifos_9_reset),
    .io_in_ready(fifos_9_io_in_ready),
    .io_in_valid(fifos_9_io_in_valid),
    .io_in_bits(fifos_9_io_in_bits),
    .io_out_ready(fifos_9_io_out_ready),
    .io_out_valid(fifos_9_io_out_valid),
    .io_out_bits(fifos_9_io_out_bits)
  );
  FIFO_1 fifos_10 ( // @[FIFOVec.scala 40:19:@12944.4]
    .clock(fifos_10_clock),
    .reset(fifos_10_reset),
    .io_in_ready(fifos_10_io_in_ready),
    .io_in_valid(fifos_10_io_in_valid),
    .io_in_bits(fifos_10_io_in_bits),
    .io_out_ready(fifos_10_io_out_ready),
    .io_out_valid(fifos_10_io_out_valid),
    .io_out_bits(fifos_10_io_out_bits)
  );
  FIFO_1 fifos_11 ( // @[FIFOVec.scala 40:19:@12979.4]
    .clock(fifos_11_clock),
    .reset(fifos_11_reset),
    .io_in_ready(fifos_11_io_in_ready),
    .io_in_valid(fifos_11_io_in_valid),
    .io_in_bits(fifos_11_io_in_bits),
    .io_out_ready(fifos_11_io_out_ready),
    .io_out_valid(fifos_11_io_out_valid),
    .io_out_bits(fifos_11_io_out_bits)
  );
  FIFO_1 fifos_12 ( // @[FIFOVec.scala 40:19:@13014.4]
    .clock(fifos_12_clock),
    .reset(fifos_12_reset),
    .io_in_ready(fifos_12_io_in_ready),
    .io_in_valid(fifos_12_io_in_valid),
    .io_in_bits(fifos_12_io_in_bits),
    .io_out_ready(fifos_12_io_out_ready),
    .io_out_valid(fifos_12_io_out_valid),
    .io_out_bits(fifos_12_io_out_bits)
  );
  FIFO_1 fifos_13 ( // @[FIFOVec.scala 40:19:@13049.4]
    .clock(fifos_13_clock),
    .reset(fifos_13_reset),
    .io_in_ready(fifos_13_io_in_ready),
    .io_in_valid(fifos_13_io_in_valid),
    .io_in_bits(fifos_13_io_in_bits),
    .io_out_ready(fifos_13_io_out_ready),
    .io_out_valid(fifos_13_io_out_valid),
    .io_out_bits(fifos_13_io_out_bits)
  );
  FIFO_1 fifos_14 ( // @[FIFOVec.scala 40:19:@13084.4]
    .clock(fifos_14_clock),
    .reset(fifos_14_reset),
    .io_in_ready(fifos_14_io_in_ready),
    .io_in_valid(fifos_14_io_in_valid),
    .io_in_bits(fifos_14_io_in_bits),
    .io_out_ready(fifos_14_io_out_ready),
    .io_out_valid(fifos_14_io_out_valid),
    .io_out_bits(fifos_14_io_out_bits)
  );
  FIFO_1 fifos_15 ( // @[FIFOVec.scala 40:19:@13119.4]
    .clock(fifos_15_clock),
    .reset(fifos_15_reset),
    .io_in_ready(fifos_15_io_in_ready),
    .io_in_valid(fifos_15_io_in_valid),
    .io_in_bits(fifos_15_io_in_bits),
    .io_out_ready(fifos_15_io_out_ready),
    .io_out_valid(fifos_15_io_out_valid),
    .io_out_bits(fifos_15_io_out_bits)
  );
  assign readEn = io_out_valid & io_out_ready; // @[FIFOVec.scala 20:29:@12568.4]
  assign deqDecoder = 16'h1 << deqCounter_io_out; // @[OneHot.scala 45:35:@12593.4]
  assign _T_154 = deqDecoder[0]; // @[FIFOVec.scala 44:50:@12625.4]
  assign _T_163 = deqDecoder[1]; // @[FIFOVec.scala 44:50:@12660.4]
  assign _T_172 = deqDecoder[2]; // @[FIFOVec.scala 44:50:@12695.4]
  assign _T_181 = deqDecoder[3]; // @[FIFOVec.scala 44:50:@12730.4]
  assign _T_190 = deqDecoder[4]; // @[FIFOVec.scala 44:50:@12765.4]
  assign _T_199 = deqDecoder[5]; // @[FIFOVec.scala 44:50:@12800.4]
  assign _T_208 = deqDecoder[6]; // @[FIFOVec.scala 44:50:@12835.4]
  assign _T_217 = deqDecoder[7]; // @[FIFOVec.scala 44:50:@12870.4]
  assign _T_226 = deqDecoder[8]; // @[FIFOVec.scala 44:50:@12905.4]
  assign _T_235 = deqDecoder[9]; // @[FIFOVec.scala 44:50:@12940.4]
  assign _T_244 = deqDecoder[10]; // @[FIFOVec.scala 44:50:@12975.4]
  assign _T_253 = deqDecoder[11]; // @[FIFOVec.scala 44:50:@13010.4]
  assign _T_262 = deqDecoder[12]; // @[FIFOVec.scala 44:50:@13045.4]
  assign _T_271 = deqDecoder[13]; // @[FIFOVec.scala 44:50:@13080.4]
  assign _T_280 = deqDecoder[14]; // @[FIFOVec.scala 44:50:@13115.4]
  assign _T_289 = deqDecoder[15]; // @[FIFOVec.scala 44:50:@13150.4]
  assign _T_316 = fifos_0_io_in_ready & fifos_1_io_in_ready; // @[FIFOVec.scala 49:90:@13171.4]
  assign _T_317 = _T_316 & fifos_2_io_in_ready; // @[FIFOVec.scala 49:90:@13172.4]
  assign _T_318 = _T_317 & fifos_3_io_in_ready; // @[FIFOVec.scala 49:90:@13173.4]
  assign _T_319 = _T_318 & fifos_4_io_in_ready; // @[FIFOVec.scala 49:90:@13174.4]
  assign _T_320 = _T_319 & fifos_5_io_in_ready; // @[FIFOVec.scala 49:90:@13175.4]
  assign _T_321 = _T_320 & fifos_6_io_in_ready; // @[FIFOVec.scala 49:90:@13176.4]
  assign _T_322 = _T_321 & fifos_7_io_in_ready; // @[FIFOVec.scala 49:90:@13177.4]
  assign _T_323 = _T_322 & fifos_8_io_in_ready; // @[FIFOVec.scala 49:90:@13178.4]
  assign _T_324 = _T_323 & fifos_9_io_in_ready; // @[FIFOVec.scala 49:90:@13179.4]
  assign _T_325 = _T_324 & fifos_10_io_in_ready; // @[FIFOVec.scala 49:90:@13180.4]
  assign _T_326 = _T_325 & fifos_11_io_in_ready; // @[FIFOVec.scala 49:90:@13181.4]
  assign _T_327 = _T_326 & fifos_12_io_in_ready; // @[FIFOVec.scala 49:90:@13182.4]
  assign _T_328 = _T_327 & fifos_13_io_in_ready; // @[FIFOVec.scala 49:90:@13183.4]
  assign _T_329 = _T_328 & fifos_14_io_in_ready; // @[FIFOVec.scala 49:90:@13184.4]
  assign _T_335_0 = fifos_0_io_out_valid; // @[FIFOVec.scala 51:43:@13188.4 FIFOVec.scala 51:43:@13189.4]
  assign _T_335_1 = fifos_1_io_out_valid; // @[FIFOVec.scala 51:43:@13188.4 FIFOVec.scala 51:43:@13190.4]
  assign _GEN_17 = 4'h1 == deqCounter_io_out ? _T_335_1 : _T_335_0; // @[FIFOVec.scala 51:22:@13220.4]
  assign _T_335_2 = fifos_2_io_out_valid; // @[FIFOVec.scala 51:43:@13188.4 FIFOVec.scala 51:43:@13191.4]
  assign _GEN_18 = 4'h2 == deqCounter_io_out ? _T_335_2 : _GEN_17; // @[FIFOVec.scala 51:22:@13220.4]
  assign _T_335_3 = fifos_3_io_out_valid; // @[FIFOVec.scala 51:43:@13188.4 FIFOVec.scala 51:43:@13192.4]
  assign _GEN_19 = 4'h3 == deqCounter_io_out ? _T_335_3 : _GEN_18; // @[FIFOVec.scala 51:22:@13220.4]
  assign _T_335_4 = fifos_4_io_out_valid; // @[FIFOVec.scala 51:43:@13188.4 FIFOVec.scala 51:43:@13193.4]
  assign _GEN_20 = 4'h4 == deqCounter_io_out ? _T_335_4 : _GEN_19; // @[FIFOVec.scala 51:22:@13220.4]
  assign _T_335_5 = fifos_5_io_out_valid; // @[FIFOVec.scala 51:43:@13188.4 FIFOVec.scala 51:43:@13194.4]
  assign _GEN_21 = 4'h5 == deqCounter_io_out ? _T_335_5 : _GEN_20; // @[FIFOVec.scala 51:22:@13220.4]
  assign _T_335_6 = fifos_6_io_out_valid; // @[FIFOVec.scala 51:43:@13188.4 FIFOVec.scala 51:43:@13195.4]
  assign _GEN_22 = 4'h6 == deqCounter_io_out ? _T_335_6 : _GEN_21; // @[FIFOVec.scala 51:22:@13220.4]
  assign _T_335_7 = fifos_7_io_out_valid; // @[FIFOVec.scala 51:43:@13188.4 FIFOVec.scala 51:43:@13196.4]
  assign _GEN_23 = 4'h7 == deqCounter_io_out ? _T_335_7 : _GEN_22; // @[FIFOVec.scala 51:22:@13220.4]
  assign _T_335_8 = fifos_8_io_out_valid; // @[FIFOVec.scala 51:43:@13188.4 FIFOVec.scala 51:43:@13197.4]
  assign _GEN_24 = 4'h8 == deqCounter_io_out ? _T_335_8 : _GEN_23; // @[FIFOVec.scala 51:22:@13220.4]
  assign _T_335_9 = fifos_9_io_out_valid; // @[FIFOVec.scala 51:43:@13188.4 FIFOVec.scala 51:43:@13198.4]
  assign _GEN_25 = 4'h9 == deqCounter_io_out ? _T_335_9 : _GEN_24; // @[FIFOVec.scala 51:22:@13220.4]
  assign _T_335_10 = fifos_10_io_out_valid; // @[FIFOVec.scala 51:43:@13188.4 FIFOVec.scala 51:43:@13199.4]
  assign _GEN_26 = 4'ha == deqCounter_io_out ? _T_335_10 : _GEN_25; // @[FIFOVec.scala 51:22:@13220.4]
  assign _T_335_11 = fifos_11_io_out_valid; // @[FIFOVec.scala 51:43:@13188.4 FIFOVec.scala 51:43:@13200.4]
  assign _GEN_27 = 4'hb == deqCounter_io_out ? _T_335_11 : _GEN_26; // @[FIFOVec.scala 51:22:@13220.4]
  assign _T_335_12 = fifos_12_io_out_valid; // @[FIFOVec.scala 51:43:@13188.4 FIFOVec.scala 51:43:@13201.4]
  assign _GEN_28 = 4'hc == deqCounter_io_out ? _T_335_12 : _GEN_27; // @[FIFOVec.scala 51:22:@13220.4]
  assign _T_335_13 = fifos_13_io_out_valid; // @[FIFOVec.scala 51:43:@13188.4 FIFOVec.scala 51:43:@13202.4]
  assign _GEN_29 = 4'hd == deqCounter_io_out ? _T_335_13 : _GEN_28; // @[FIFOVec.scala 51:22:@13220.4]
  assign _T_335_14 = fifos_14_io_out_valid; // @[FIFOVec.scala 51:43:@13188.4 FIFOVec.scala 51:43:@13203.4]
  assign _GEN_30 = 4'he == deqCounter_io_out ? _T_335_14 : _GEN_29; // @[FIFOVec.scala 51:22:@13220.4]
  assign _T_335_15 = fifos_15_io_out_valid; // @[FIFOVec.scala 51:43:@13188.4 FIFOVec.scala 51:43:@13204.4]
  assign _T_374_0 = fifos_0_io_out_bits; // @[FIFOVec.scala 53:65:@13222.4 FIFOVec.scala 53:65:@13223.4]
  assign _T_374_1 = fifos_1_io_out_bits; // @[FIFOVec.scala 53:65:@13222.4 FIFOVec.scala 53:65:@13224.4]
  assign _GEN_33 = 4'h1 == deqCounter_io_out ? _T_374_1 : _T_374_0; // @[FIFOVec.scala 53:42:@13495.4]
  assign _T_374_2 = fifos_2_io_out_bits; // @[FIFOVec.scala 53:65:@13222.4 FIFOVec.scala 53:65:@13225.4]
  assign _GEN_34 = 4'h2 == deqCounter_io_out ? _T_374_2 : _GEN_33; // @[FIFOVec.scala 53:42:@13495.4]
  assign _T_374_3 = fifos_3_io_out_bits; // @[FIFOVec.scala 53:65:@13222.4 FIFOVec.scala 53:65:@13226.4]
  assign _GEN_35 = 4'h3 == deqCounter_io_out ? _T_374_3 : _GEN_34; // @[FIFOVec.scala 53:42:@13495.4]
  assign _T_374_4 = fifos_4_io_out_bits; // @[FIFOVec.scala 53:65:@13222.4 FIFOVec.scala 53:65:@13227.4]
  assign _GEN_36 = 4'h4 == deqCounter_io_out ? _T_374_4 : _GEN_35; // @[FIFOVec.scala 53:42:@13495.4]
  assign _T_374_5 = fifos_5_io_out_bits; // @[FIFOVec.scala 53:65:@13222.4 FIFOVec.scala 53:65:@13228.4]
  assign _GEN_37 = 4'h5 == deqCounter_io_out ? _T_374_5 : _GEN_36; // @[FIFOVec.scala 53:42:@13495.4]
  assign _T_374_6 = fifos_6_io_out_bits; // @[FIFOVec.scala 53:65:@13222.4 FIFOVec.scala 53:65:@13229.4]
  assign _GEN_38 = 4'h6 == deqCounter_io_out ? _T_374_6 : _GEN_37; // @[FIFOVec.scala 53:42:@13495.4]
  assign _T_374_7 = fifos_7_io_out_bits; // @[FIFOVec.scala 53:65:@13222.4 FIFOVec.scala 53:65:@13230.4]
  assign _GEN_39 = 4'h7 == deqCounter_io_out ? _T_374_7 : _GEN_38; // @[FIFOVec.scala 53:42:@13495.4]
  assign _T_374_8 = fifos_8_io_out_bits; // @[FIFOVec.scala 53:65:@13222.4 FIFOVec.scala 53:65:@13231.4]
  assign _GEN_40 = 4'h8 == deqCounter_io_out ? _T_374_8 : _GEN_39; // @[FIFOVec.scala 53:42:@13495.4]
  assign _T_374_9 = fifos_9_io_out_bits; // @[FIFOVec.scala 53:65:@13222.4 FIFOVec.scala 53:65:@13232.4]
  assign _GEN_41 = 4'h9 == deqCounter_io_out ? _T_374_9 : _GEN_40; // @[FIFOVec.scala 53:42:@13495.4]
  assign _T_374_10 = fifos_10_io_out_bits; // @[FIFOVec.scala 53:65:@13222.4 FIFOVec.scala 53:65:@13233.4]
  assign _GEN_42 = 4'ha == deqCounter_io_out ? _T_374_10 : _GEN_41; // @[FIFOVec.scala 53:42:@13495.4]
  assign _T_374_11 = fifos_11_io_out_bits; // @[FIFOVec.scala 53:65:@13222.4 FIFOVec.scala 53:65:@13234.4]
  assign _GEN_43 = 4'hb == deqCounter_io_out ? _T_374_11 : _GEN_42; // @[FIFOVec.scala 53:42:@13495.4]
  assign _T_374_12 = fifos_12_io_out_bits; // @[FIFOVec.scala 53:65:@13222.4 FIFOVec.scala 53:65:@13235.4]
  assign _GEN_44 = 4'hc == deqCounter_io_out ? _T_374_12 : _GEN_43; // @[FIFOVec.scala 53:42:@13495.4]
  assign _T_374_13 = fifos_13_io_out_bits; // @[FIFOVec.scala 53:65:@13222.4 FIFOVec.scala 53:65:@13236.4]
  assign _GEN_45 = 4'hd == deqCounter_io_out ? _T_374_13 : _GEN_44; // @[FIFOVec.scala 53:42:@13495.4]
  assign _T_374_14 = fifos_14_io_out_bits; // @[FIFOVec.scala 53:65:@13222.4 FIFOVec.scala 53:65:@13237.4]
  assign _GEN_46 = 4'he == deqCounter_io_out ? _T_374_14 : _GEN_45; // @[FIFOVec.scala 53:42:@13495.4]
  assign _T_374_15 = fifos_15_io_out_bits; // @[FIFOVec.scala 53:65:@13222.4 FIFOVec.scala 53:65:@13238.4]
  assign io_in_ready = _T_329 & fifos_15_io_in_ready; // @[FIFOVec.scala 49:15:@13187.4]
  assign io_out_valid = 4'hf == deqCounter_io_out ? _T_335_15 : _GEN_30; // @[FIFOVec.scala 51:16:@13221.4]
  assign io_out_bits_0 = 4'hf == deqCounter_io_out ? _T_374_15 : _GEN_46; // @[FIFOVec.scala 53:15:@13529.4]
  assign enqCounter_clock = clock; // @[:@12571.4]
  assign enqCounter_reset = reset; // @[:@12572.4]
  assign enqCounter_io_enable = 1'h0; // @[FIFOVec.scala 26:24:@12579.4]
  assign deqCounter_clock = clock; // @[:@12582.4]
  assign deqCounter_reset = reset; // @[:@12583.4]
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFOVec.scala 30:24:@12590.4]
  assign fifos_0_clock = clock; // @[:@12595.4]
  assign fifos_0_reset = reset; // @[:@12596.4]
  assign fifos_0_io_in_valid = io_in_valid & io_in_ready; // @[FIFOVec.scala 42:19:@12622.4]
  assign fifos_0_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@12624.4]
  assign fifos_0_io_out_ready = _T_154 & readEn; // @[FIFOVec.scala 44:20:@12628.4]
  assign fifos_1_clock = clock; // @[:@12630.4]
  assign fifos_1_reset = reset; // @[:@12631.4]
  assign fifos_1_io_in_valid = io_in_valid & io_in_ready; // @[FIFOVec.scala 42:19:@12657.4]
  assign fifos_1_io_in_bits = io_in_bits_1; // @[FIFOVec.scala 43:18:@12659.4]
  assign fifos_1_io_out_ready = _T_163 & readEn; // @[FIFOVec.scala 44:20:@12663.4]
  assign fifos_2_clock = clock; // @[:@12665.4]
  assign fifos_2_reset = reset; // @[:@12666.4]
  assign fifos_2_io_in_valid = io_in_valid & io_in_ready; // @[FIFOVec.scala 42:19:@12692.4]
  assign fifos_2_io_in_bits = io_in_bits_2; // @[FIFOVec.scala 43:18:@12694.4]
  assign fifos_2_io_out_ready = _T_172 & readEn; // @[FIFOVec.scala 44:20:@12698.4]
  assign fifos_3_clock = clock; // @[:@12700.4]
  assign fifos_3_reset = reset; // @[:@12701.4]
  assign fifos_3_io_in_valid = io_in_valid & io_in_ready; // @[FIFOVec.scala 42:19:@12727.4]
  assign fifos_3_io_in_bits = io_in_bits_3; // @[FIFOVec.scala 43:18:@12729.4]
  assign fifos_3_io_out_ready = _T_181 & readEn; // @[FIFOVec.scala 44:20:@12733.4]
  assign fifos_4_clock = clock; // @[:@12735.4]
  assign fifos_4_reset = reset; // @[:@12736.4]
  assign fifos_4_io_in_valid = io_in_valid & io_in_ready; // @[FIFOVec.scala 42:19:@12762.4]
  assign fifos_4_io_in_bits = io_in_bits_4; // @[FIFOVec.scala 43:18:@12764.4]
  assign fifos_4_io_out_ready = _T_190 & readEn; // @[FIFOVec.scala 44:20:@12768.4]
  assign fifos_5_clock = clock; // @[:@12770.4]
  assign fifos_5_reset = reset; // @[:@12771.4]
  assign fifos_5_io_in_valid = io_in_valid & io_in_ready; // @[FIFOVec.scala 42:19:@12797.4]
  assign fifos_5_io_in_bits = io_in_bits_5; // @[FIFOVec.scala 43:18:@12799.4]
  assign fifos_5_io_out_ready = _T_199 & readEn; // @[FIFOVec.scala 44:20:@12803.4]
  assign fifos_6_clock = clock; // @[:@12805.4]
  assign fifos_6_reset = reset; // @[:@12806.4]
  assign fifos_6_io_in_valid = io_in_valid & io_in_ready; // @[FIFOVec.scala 42:19:@12832.4]
  assign fifos_6_io_in_bits = io_in_bits_6; // @[FIFOVec.scala 43:18:@12834.4]
  assign fifos_6_io_out_ready = _T_208 & readEn; // @[FIFOVec.scala 44:20:@12838.4]
  assign fifos_7_clock = clock; // @[:@12840.4]
  assign fifos_7_reset = reset; // @[:@12841.4]
  assign fifos_7_io_in_valid = io_in_valid & io_in_ready; // @[FIFOVec.scala 42:19:@12867.4]
  assign fifos_7_io_in_bits = io_in_bits_7; // @[FIFOVec.scala 43:18:@12869.4]
  assign fifos_7_io_out_ready = _T_217 & readEn; // @[FIFOVec.scala 44:20:@12873.4]
  assign fifos_8_clock = clock; // @[:@12875.4]
  assign fifos_8_reset = reset; // @[:@12876.4]
  assign fifos_8_io_in_valid = io_in_valid & io_in_ready; // @[FIFOVec.scala 42:19:@12902.4]
  assign fifos_8_io_in_bits = io_in_bits_8; // @[FIFOVec.scala 43:18:@12904.4]
  assign fifos_8_io_out_ready = _T_226 & readEn; // @[FIFOVec.scala 44:20:@12908.4]
  assign fifos_9_clock = clock; // @[:@12910.4]
  assign fifos_9_reset = reset; // @[:@12911.4]
  assign fifos_9_io_in_valid = io_in_valid & io_in_ready; // @[FIFOVec.scala 42:19:@12937.4]
  assign fifos_9_io_in_bits = io_in_bits_9; // @[FIFOVec.scala 43:18:@12939.4]
  assign fifos_9_io_out_ready = _T_235 & readEn; // @[FIFOVec.scala 44:20:@12943.4]
  assign fifos_10_clock = clock; // @[:@12945.4]
  assign fifos_10_reset = reset; // @[:@12946.4]
  assign fifos_10_io_in_valid = io_in_valid & io_in_ready; // @[FIFOVec.scala 42:19:@12972.4]
  assign fifos_10_io_in_bits = io_in_bits_10; // @[FIFOVec.scala 43:18:@12974.4]
  assign fifos_10_io_out_ready = _T_244 & readEn; // @[FIFOVec.scala 44:20:@12978.4]
  assign fifos_11_clock = clock; // @[:@12980.4]
  assign fifos_11_reset = reset; // @[:@12981.4]
  assign fifos_11_io_in_valid = io_in_valid & io_in_ready; // @[FIFOVec.scala 42:19:@13007.4]
  assign fifos_11_io_in_bits = io_in_bits_11; // @[FIFOVec.scala 43:18:@13009.4]
  assign fifos_11_io_out_ready = _T_253 & readEn; // @[FIFOVec.scala 44:20:@13013.4]
  assign fifos_12_clock = clock; // @[:@13015.4]
  assign fifos_12_reset = reset; // @[:@13016.4]
  assign fifos_12_io_in_valid = io_in_valid & io_in_ready; // @[FIFOVec.scala 42:19:@13042.4]
  assign fifos_12_io_in_bits = io_in_bits_12; // @[FIFOVec.scala 43:18:@13044.4]
  assign fifos_12_io_out_ready = _T_262 & readEn; // @[FIFOVec.scala 44:20:@13048.4]
  assign fifos_13_clock = clock; // @[:@13050.4]
  assign fifos_13_reset = reset; // @[:@13051.4]
  assign fifos_13_io_in_valid = io_in_valid & io_in_ready; // @[FIFOVec.scala 42:19:@13077.4]
  assign fifos_13_io_in_bits = io_in_bits_13; // @[FIFOVec.scala 43:18:@13079.4]
  assign fifos_13_io_out_ready = _T_271 & readEn; // @[FIFOVec.scala 44:20:@13083.4]
  assign fifos_14_clock = clock; // @[:@13085.4]
  assign fifos_14_reset = reset; // @[:@13086.4]
  assign fifos_14_io_in_valid = io_in_valid & io_in_ready; // @[FIFOVec.scala 42:19:@13112.4]
  assign fifos_14_io_in_bits = io_in_bits_14; // @[FIFOVec.scala 43:18:@13114.4]
  assign fifos_14_io_out_ready = _T_280 & readEn; // @[FIFOVec.scala 44:20:@13118.4]
  assign fifos_15_clock = clock; // @[:@13120.4]
  assign fifos_15_reset = reset; // @[:@13121.4]
  assign fifos_15_io_in_valid = io_in_valid & io_in_ready; // @[FIFOVec.scala 42:19:@13147.4]
  assign fifos_15_io_in_bits = io_in_bits_15; // @[FIFOVec.scala 43:18:@13149.4]
  assign fifos_15_io_out_ready = _T_289 & readEn; // @[FIFOVec.scala 44:20:@13153.4]
endmodule
module SRAM_17( // @[:@13634.2]
  input        clock, // @[:@13635.4]
  input  [5:0] io_raddr, // @[:@13637.4]
  input        io_wen, // @[:@13637.4]
  input  [5:0] io_waddr // @[:@13637.4]
);
  wire [15:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 124:30:@13639.4]
  wire [15:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 124:30:@13639.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 124:30:@13639.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 124:30:@13639.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 124:30:@13639.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 124:30:@13639.4]
  wire [5:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 124:30:@13639.4]
  wire [5:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 124:30:@13639.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 124:30:@13639.4]
  SRAMVerilogAWS #(.DWIDTH(16), .WORDS(64), .AWIDTH(6)) SRAMVerilogAWS ( // @[SRAM.scala 124:30:@13639.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign SRAMVerilogAWS_wdata = 16'h0; // @[SRAM.scala 130:20:@13653.4]
  assign SRAMVerilogAWS_backpressure = 1'h1; // @[SRAM.scala 131:27:@13654.4]
  assign SRAMVerilogAWS_wen = io_wen; // @[SRAM.scala 128:18:@13651.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 133:22:@13656.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 132:22:@13655.4]
  assign SRAMVerilogAWS_waddr = io_waddr; // @[SRAM.scala 129:20:@13652.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 127:20:@13650.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 126:18:@13649.4]
endmodule
module FIFO_17( // @[:@13668.2]
  input   clock, // @[:@13669.4]
  input   reset, // @[:@13670.4]
  output  io_in_ready, // @[:@13671.4]
  input   io_in_valid // @[:@13671.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@13937.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@13937.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@13937.4]
  wire [5:0] enqCounter_io_out; // @[FIFO.scala 34:26:@13937.4]
  wire [5:0] enqCounter_io_next; // @[FIFO.scala 34:26:@13937.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@13947.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@13947.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@13947.4]
  wire [5:0] deqCounter_io_out; // @[FIFO.scala 38:26:@13947.4]
  wire [5:0] deqCounter_io_next; // @[FIFO.scala 38:26:@13947.4]
  wire  SRAM_clock; // @[FIFO.scala 73:19:@13962.4]
  wire [5:0] SRAM_io_raddr; // @[FIFO.scala 73:19:@13962.4]
  wire  SRAM_io_wen; // @[FIFO.scala 73:19:@13962.4]
  wire [5:0] SRAM_io_waddr; // @[FIFO.scala 73:19:@13962.4]
  wire  writeEn; // @[FIFO.scala 30:29:@13935.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@13957.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@13958.4]
  wire  full; // @[FIFO.scala 46:23:@13961.4]
  wire  _GEN_0; // @[FIFO.scala 83:29:@13973.4]
  Counter enqCounter ( // @[FIFO.scala 34:26:@13937.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter deqCounter ( // @[FIFO.scala 38:26:@13947.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  SRAM_17 SRAM ( // @[FIFO.scala 73:19:@13962.4]
    .clock(SRAM_clock),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@13935.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@13958.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@13961.4]
  assign _GEN_0 = writeEn ? writeEn : maybeFull; // @[FIFO.scala 83:29:@13973.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@13979.4]
  assign enqCounter_clock = clock; // @[:@13938.4]
  assign enqCounter_reset = reset; // @[:@13939.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@13945.4]
  assign deqCounter_clock = clock; // @[:@13948.4]
  assign deqCounter_reset = reset; // @[:@13949.4]
  assign deqCounter_io_enable = 1'h0; // @[FIFO.scala 40:24:@13955.4]
  assign SRAM_clock = clock; // @[:@13963.4]
  assign SRAM_io_raddr = deqCounter_io_out; // @[FIFO.scala 75:16:@13966.4]
  assign SRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 76:14:@13967.4]
  assign SRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 77:16:@13968.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (writeEn) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module FIFOVec_1( // @[:@13981.2]
  input   clock, // @[:@13982.4]
  input   reset, // @[:@13983.4]
  output  io_in_ready, // @[:@13984.4]
  input   io_in_valid // @[:@13984.4]
);
  wire  fifos_0_clock; // @[FIFOVec.scala 40:19:@14012.4]
  wire  fifos_0_reset; // @[FIFOVec.scala 40:19:@14012.4]
  wire  fifos_0_io_in_ready; // @[FIFOVec.scala 40:19:@14012.4]
  wire  fifos_0_io_in_valid; // @[FIFOVec.scala 40:19:@14012.4]
  FIFO_17 fifos_0 ( // @[FIFOVec.scala 40:19:@14012.4]
    .clock(fifos_0_clock),
    .reset(fifos_0_reset),
    .io_in_ready(fifos_0_io_in_ready),
    .io_in_valid(fifos_0_io_in_valid)
  );
  assign io_in_ready = fifos_0_io_in_ready; // @[FIFOVec.scala 49:15:@14290.4]
  assign fifos_0_clock = clock; // @[:@14013.4]
  assign fifos_0_reset = reset; // @[:@14014.4]
  assign fifos_0_io_in_valid = io_in_valid & io_in_ready; // @[FIFOVec.scala 42:19:@14280.4]
endmodule
module FIFOWidthConvert( // @[:@14304.2]
  input         clock, // @[:@14305.4]
  input         reset, // @[:@14306.4]
  output        io_in_ready, // @[:@14307.4]
  input         io_in_valid, // @[:@14307.4]
  input  [31:0] io_in_bits_data_0, // @[:@14307.4]
  input  [31:0] io_in_bits_data_1, // @[:@14307.4]
  input  [31:0] io_in_bits_data_2, // @[:@14307.4]
  input  [31:0] io_in_bits_data_3, // @[:@14307.4]
  input  [31:0] io_in_bits_data_4, // @[:@14307.4]
  input  [31:0] io_in_bits_data_5, // @[:@14307.4]
  input  [31:0] io_in_bits_data_6, // @[:@14307.4]
  input  [31:0] io_in_bits_data_7, // @[:@14307.4]
  input  [31:0] io_in_bits_data_8, // @[:@14307.4]
  input  [31:0] io_in_bits_data_9, // @[:@14307.4]
  input  [31:0] io_in_bits_data_10, // @[:@14307.4]
  input  [31:0] io_in_bits_data_11, // @[:@14307.4]
  input  [31:0] io_in_bits_data_12, // @[:@14307.4]
  input  [31:0] io_in_bits_data_13, // @[:@14307.4]
  input  [31:0] io_in_bits_data_14, // @[:@14307.4]
  input  [31:0] io_in_bits_data_15, // @[:@14307.4]
  input         io_out_ready, // @[:@14307.4]
  output        io_out_valid, // @[:@14307.4]
  output [31:0] io_out_bits_data_0 // @[:@14307.4]
);
  wire  FIFOVec_clock; // @[FIFOWidthConvert.scala 82:22:@14309.4]
  wire  FIFOVec_reset; // @[FIFOWidthConvert.scala 82:22:@14309.4]
  wire  FIFOVec_io_in_ready; // @[FIFOWidthConvert.scala 82:22:@14309.4]
  wire  FIFOVec_io_in_valid; // @[FIFOWidthConvert.scala 82:22:@14309.4]
  wire [31:0] FIFOVec_io_in_bits_0; // @[FIFOWidthConvert.scala 82:22:@14309.4]
  wire [31:0] FIFOVec_io_in_bits_1; // @[FIFOWidthConvert.scala 82:22:@14309.4]
  wire [31:0] FIFOVec_io_in_bits_2; // @[FIFOWidthConvert.scala 82:22:@14309.4]
  wire [31:0] FIFOVec_io_in_bits_3; // @[FIFOWidthConvert.scala 82:22:@14309.4]
  wire [31:0] FIFOVec_io_in_bits_4; // @[FIFOWidthConvert.scala 82:22:@14309.4]
  wire [31:0] FIFOVec_io_in_bits_5; // @[FIFOWidthConvert.scala 82:22:@14309.4]
  wire [31:0] FIFOVec_io_in_bits_6; // @[FIFOWidthConvert.scala 82:22:@14309.4]
  wire [31:0] FIFOVec_io_in_bits_7; // @[FIFOWidthConvert.scala 82:22:@14309.4]
  wire [31:0] FIFOVec_io_in_bits_8; // @[FIFOWidthConvert.scala 82:22:@14309.4]
  wire [31:0] FIFOVec_io_in_bits_9; // @[FIFOWidthConvert.scala 82:22:@14309.4]
  wire [31:0] FIFOVec_io_in_bits_10; // @[FIFOWidthConvert.scala 82:22:@14309.4]
  wire [31:0] FIFOVec_io_in_bits_11; // @[FIFOWidthConvert.scala 82:22:@14309.4]
  wire [31:0] FIFOVec_io_in_bits_12; // @[FIFOWidthConvert.scala 82:22:@14309.4]
  wire [31:0] FIFOVec_io_in_bits_13; // @[FIFOWidthConvert.scala 82:22:@14309.4]
  wire [31:0] FIFOVec_io_in_bits_14; // @[FIFOWidthConvert.scala 82:22:@14309.4]
  wire [31:0] FIFOVec_io_in_bits_15; // @[FIFOWidthConvert.scala 82:22:@14309.4]
  wire  FIFOVec_io_out_ready; // @[FIFOWidthConvert.scala 82:22:@14309.4]
  wire  FIFOVec_io_out_valid; // @[FIFOWidthConvert.scala 82:22:@14309.4]
  wire [31:0] FIFOVec_io_out_bits_0; // @[FIFOWidthConvert.scala 82:22:@14309.4]
  wire  FIFOVec_1_clock; // @[FIFOWidthConvert.scala 83:26:@14350.4]
  wire  FIFOVec_1_reset; // @[FIFOWidthConvert.scala 83:26:@14350.4]
  wire  FIFOVec_1_io_in_ready; // @[FIFOWidthConvert.scala 83:26:@14350.4]
  wire  FIFOVec_1_io_in_valid; // @[FIFOWidthConvert.scala 83:26:@14350.4]
  wire [319:0] _T_55; // @[Cat.scala 30:58:@14375.4]
  wire [511:0] _T_61; // @[Cat.scala 30:58:@14381.4]
  FIFOVec FIFOVec ( // @[FIFOWidthConvert.scala 82:22:@14309.4]
    .clock(FIFOVec_clock),
    .reset(FIFOVec_reset),
    .io_in_ready(FIFOVec_io_in_ready),
    .io_in_valid(FIFOVec_io_in_valid),
    .io_in_bits_0(FIFOVec_io_in_bits_0),
    .io_in_bits_1(FIFOVec_io_in_bits_1),
    .io_in_bits_2(FIFOVec_io_in_bits_2),
    .io_in_bits_3(FIFOVec_io_in_bits_3),
    .io_in_bits_4(FIFOVec_io_in_bits_4),
    .io_in_bits_5(FIFOVec_io_in_bits_5),
    .io_in_bits_6(FIFOVec_io_in_bits_6),
    .io_in_bits_7(FIFOVec_io_in_bits_7),
    .io_in_bits_8(FIFOVec_io_in_bits_8),
    .io_in_bits_9(FIFOVec_io_in_bits_9),
    .io_in_bits_10(FIFOVec_io_in_bits_10),
    .io_in_bits_11(FIFOVec_io_in_bits_11),
    .io_in_bits_12(FIFOVec_io_in_bits_12),
    .io_in_bits_13(FIFOVec_io_in_bits_13),
    .io_in_bits_14(FIFOVec_io_in_bits_14),
    .io_in_bits_15(FIFOVec_io_in_bits_15),
    .io_out_ready(FIFOVec_io_out_ready),
    .io_out_valid(FIFOVec_io_out_valid),
    .io_out_bits_0(FIFOVec_io_out_bits_0)
  );
  FIFOVec_1 FIFOVec_1 ( // @[FIFOWidthConvert.scala 83:26:@14350.4]
    .clock(FIFOVec_1_clock),
    .reset(FIFOVec_1_reset),
    .io_in_ready(FIFOVec_1_io_in_ready),
    .io_in_valid(FIFOVec_1_io_in_valid)
  );
  assign _T_55 = {io_in_bits_data_15,io_in_bits_data_14,io_in_bits_data_13,io_in_bits_data_12,io_in_bits_data_11,io_in_bits_data_10,io_in_bits_data_9,io_in_bits_data_8,io_in_bits_data_7,io_in_bits_data_6}; // @[Cat.scala 30:58:@14375.4]
  assign _T_61 = {_T_55,io_in_bits_data_5,io_in_bits_data_4,io_in_bits_data_3,io_in_bits_data_2,io_in_bits_data_1,io_in_bits_data_0}; // @[Cat.scala 30:58:@14381.4]
  assign io_in_ready = FIFOVec_io_in_ready; // @[FIFOWidthConvert.scala 88:17:@14365.4]
  assign io_out_valid = FIFOVec_io_out_valid; // @[FIFOWidthConvert.scala 89:18:@14366.4]
  assign io_out_bits_data_0 = FIFOVec_io_out_bits_0; // @[FIFOWidthConvert.scala 96:22:@14439.4]
  assign FIFOVec_clock = clock; // @[:@14310.4]
  assign FIFOVec_reset = reset; // @[:@14311.4]
  assign FIFOVec_io_in_valid = io_in_valid; // @[FIFOWidthConvert.scala 92:22:@14431.4]
  assign FIFOVec_io_in_bits_0 = _T_61[31:0]; // @[FIFOWidthConvert.scala 91:21:@14415.4]
  assign FIFOVec_io_in_bits_1 = _T_61[63:32]; // @[FIFOWidthConvert.scala 91:21:@14416.4]
  assign FIFOVec_io_in_bits_2 = _T_61[95:64]; // @[FIFOWidthConvert.scala 91:21:@14417.4]
  assign FIFOVec_io_in_bits_3 = _T_61[127:96]; // @[FIFOWidthConvert.scala 91:21:@14418.4]
  assign FIFOVec_io_in_bits_4 = _T_61[159:128]; // @[FIFOWidthConvert.scala 91:21:@14419.4]
  assign FIFOVec_io_in_bits_5 = _T_61[191:160]; // @[FIFOWidthConvert.scala 91:21:@14420.4]
  assign FIFOVec_io_in_bits_6 = _T_61[223:192]; // @[FIFOWidthConvert.scala 91:21:@14421.4]
  assign FIFOVec_io_in_bits_7 = _T_61[255:224]; // @[FIFOWidthConvert.scala 91:21:@14422.4]
  assign FIFOVec_io_in_bits_8 = _T_61[287:256]; // @[FIFOWidthConvert.scala 91:21:@14423.4]
  assign FIFOVec_io_in_bits_9 = _T_61[319:288]; // @[FIFOWidthConvert.scala 91:21:@14424.4]
  assign FIFOVec_io_in_bits_10 = _T_61[351:320]; // @[FIFOWidthConvert.scala 91:21:@14425.4]
  assign FIFOVec_io_in_bits_11 = _T_61[383:352]; // @[FIFOWidthConvert.scala 91:21:@14426.4]
  assign FIFOVec_io_in_bits_12 = _T_61[415:384]; // @[FIFOWidthConvert.scala 91:21:@14427.4]
  assign FIFOVec_io_in_bits_13 = _T_61[447:416]; // @[FIFOWidthConvert.scala 91:21:@14428.4]
  assign FIFOVec_io_in_bits_14 = _T_61[479:448]; // @[FIFOWidthConvert.scala 91:21:@14429.4]
  assign FIFOVec_io_in_bits_15 = _T_61[511:480]; // @[FIFOWidthConvert.scala 91:21:@14430.4]
  assign FIFOVec_io_out_ready = io_out_ready; // @[FIFOWidthConvert.scala 98:23:@14453.4]
  assign FIFOVec_1_clock = clock; // @[:@14351.4]
  assign FIFOVec_1_reset = reset; // @[:@14352.4]
  assign FIFOVec_1_io_in_valid = io_in_valid; // @[FIFOWidthConvert.scala 94:26:@14433.4]
endmodule
module StreamControllerLoad( // @[:@14455.2]
  input         clock, // @[:@14456.4]
  input         reset, // @[:@14457.4]
  input         io_dram_cmd_ready, // @[:@14458.4]
  output        io_dram_cmd_valid, // @[:@14458.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@14458.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@14458.4]
  output        io_dram_rresp_ready, // @[:@14458.4]
  input         io_dram_rresp_valid, // @[:@14458.4]
  input  [31:0] io_dram_rresp_bits_rdata_0, // @[:@14458.4]
  input  [31:0] io_dram_rresp_bits_rdata_1, // @[:@14458.4]
  input  [31:0] io_dram_rresp_bits_rdata_2, // @[:@14458.4]
  input  [31:0] io_dram_rresp_bits_rdata_3, // @[:@14458.4]
  input  [31:0] io_dram_rresp_bits_rdata_4, // @[:@14458.4]
  input  [31:0] io_dram_rresp_bits_rdata_5, // @[:@14458.4]
  input  [31:0] io_dram_rresp_bits_rdata_6, // @[:@14458.4]
  input  [31:0] io_dram_rresp_bits_rdata_7, // @[:@14458.4]
  input  [31:0] io_dram_rresp_bits_rdata_8, // @[:@14458.4]
  input  [31:0] io_dram_rresp_bits_rdata_9, // @[:@14458.4]
  input  [31:0] io_dram_rresp_bits_rdata_10, // @[:@14458.4]
  input  [31:0] io_dram_rresp_bits_rdata_11, // @[:@14458.4]
  input  [31:0] io_dram_rresp_bits_rdata_12, // @[:@14458.4]
  input  [31:0] io_dram_rresp_bits_rdata_13, // @[:@14458.4]
  input  [31:0] io_dram_rresp_bits_rdata_14, // @[:@14458.4]
  input  [31:0] io_dram_rresp_bits_rdata_15, // @[:@14458.4]
  output        io_load_cmd_ready, // @[:@14458.4]
  input         io_load_cmd_valid, // @[:@14458.4]
  input  [63:0] io_load_cmd_bits_addr, // @[:@14458.4]
  input  [31:0] io_load_cmd_bits_size, // @[:@14458.4]
  input         io_load_data_ready, // @[:@14458.4]
  output        io_load_data_valid, // @[:@14458.4]
  output [31:0] io_load_data_bits_rdata_0 // @[:@14458.4]
);
  wire  cmd_clock; // @[StreamController.scala 38:19:@14579.4]
  wire  cmd_reset; // @[StreamController.scala 38:19:@14579.4]
  wire  cmd_io_in_ready; // @[StreamController.scala 38:19:@14579.4]
  wire  cmd_io_in_valid; // @[StreamController.scala 38:19:@14579.4]
  wire [63:0] cmd_io_in_bits_addr; // @[StreamController.scala 38:19:@14579.4]
  wire [31:0] cmd_io_in_bits_size; // @[StreamController.scala 38:19:@14579.4]
  wire  cmd_io_out_ready; // @[StreamController.scala 38:19:@14579.4]
  wire  cmd_io_out_valid; // @[StreamController.scala 38:19:@14579.4]
  wire [63:0] cmd_io_out_bits_addr; // @[StreamController.scala 38:19:@14579.4]
  wire [31:0] cmd_io_out_bits_size; // @[StreamController.scala 38:19:@14579.4]
  wire  rdata_clock; // @[StreamController.scala 51:21:@14985.4]
  wire  rdata_reset; // @[StreamController.scala 51:21:@14985.4]
  wire  rdata_io_in_ready; // @[StreamController.scala 51:21:@14985.4]
  wire  rdata_io_in_valid; // @[StreamController.scala 51:21:@14985.4]
  wire [31:0] rdata_io_in_bits_data_0; // @[StreamController.scala 51:21:@14985.4]
  wire [31:0] rdata_io_in_bits_data_1; // @[StreamController.scala 51:21:@14985.4]
  wire [31:0] rdata_io_in_bits_data_2; // @[StreamController.scala 51:21:@14985.4]
  wire [31:0] rdata_io_in_bits_data_3; // @[StreamController.scala 51:21:@14985.4]
  wire [31:0] rdata_io_in_bits_data_4; // @[StreamController.scala 51:21:@14985.4]
  wire [31:0] rdata_io_in_bits_data_5; // @[StreamController.scala 51:21:@14985.4]
  wire [31:0] rdata_io_in_bits_data_6; // @[StreamController.scala 51:21:@14985.4]
  wire [31:0] rdata_io_in_bits_data_7; // @[StreamController.scala 51:21:@14985.4]
  wire [31:0] rdata_io_in_bits_data_8; // @[StreamController.scala 51:21:@14985.4]
  wire [31:0] rdata_io_in_bits_data_9; // @[StreamController.scala 51:21:@14985.4]
  wire [31:0] rdata_io_in_bits_data_10; // @[StreamController.scala 51:21:@14985.4]
  wire [31:0] rdata_io_in_bits_data_11; // @[StreamController.scala 51:21:@14985.4]
  wire [31:0] rdata_io_in_bits_data_12; // @[StreamController.scala 51:21:@14985.4]
  wire [31:0] rdata_io_in_bits_data_13; // @[StreamController.scala 51:21:@14985.4]
  wire [31:0] rdata_io_in_bits_data_14; // @[StreamController.scala 51:21:@14985.4]
  wire [31:0] rdata_io_in_bits_data_15; // @[StreamController.scala 51:21:@14985.4]
  wire  rdata_io_out_ready; // @[StreamController.scala 51:21:@14985.4]
  wire  rdata_io_out_valid; // @[StreamController.scala 51:21:@14985.4]
  wire [31:0] rdata_io_out_bits_data_0; // @[StreamController.scala 51:21:@14985.4]
  wire [25:0] _T_95; // @[StreamController.scala 21:10:@14982.4]
  FIFO cmd ( // @[StreamController.scala 38:19:@14579.4]
    .clock(cmd_clock),
    .reset(cmd_reset),
    .io_in_ready(cmd_io_in_ready),
    .io_in_valid(cmd_io_in_valid),
    .io_in_bits_addr(cmd_io_in_bits_addr),
    .io_in_bits_size(cmd_io_in_bits_size),
    .io_out_ready(cmd_io_out_ready),
    .io_out_valid(cmd_io_out_valid),
    .io_out_bits_addr(cmd_io_out_bits_addr),
    .io_out_bits_size(cmd_io_out_bits_size)
  );
  FIFOWidthConvert rdata ( // @[StreamController.scala 51:21:@14985.4]
    .clock(rdata_clock),
    .reset(rdata_reset),
    .io_in_ready(rdata_io_in_ready),
    .io_in_valid(rdata_io_in_valid),
    .io_in_bits_data_0(rdata_io_in_bits_data_0),
    .io_in_bits_data_1(rdata_io_in_bits_data_1),
    .io_in_bits_data_2(rdata_io_in_bits_data_2),
    .io_in_bits_data_3(rdata_io_in_bits_data_3),
    .io_in_bits_data_4(rdata_io_in_bits_data_4),
    .io_in_bits_data_5(rdata_io_in_bits_data_5),
    .io_in_bits_data_6(rdata_io_in_bits_data_6),
    .io_in_bits_data_7(rdata_io_in_bits_data_7),
    .io_in_bits_data_8(rdata_io_in_bits_data_8),
    .io_in_bits_data_9(rdata_io_in_bits_data_9),
    .io_in_bits_data_10(rdata_io_in_bits_data_10),
    .io_in_bits_data_11(rdata_io_in_bits_data_11),
    .io_in_bits_data_12(rdata_io_in_bits_data_12),
    .io_in_bits_data_13(rdata_io_in_bits_data_13),
    .io_in_bits_data_14(rdata_io_in_bits_data_14),
    .io_in_bits_data_15(rdata_io_in_bits_data_15),
    .io_out_ready(rdata_io_out_ready),
    .io_out_valid(rdata_io_out_valid),
    .io_out_bits_data_0(rdata_io_out_bits_data_0)
  );
  assign _T_95 = cmd_io_out_bits_size[31:6]; // @[StreamController.scala 21:10:@14982.4]
  assign io_dram_cmd_valid = cmd_io_out_valid; // @[StreamController.scala 44:21:@14979.4]
  assign io_dram_cmd_bits_addr = cmd_io_out_bits_addr; // @[StreamController.scala 46:25:@14980.4]
  assign io_dram_cmd_bits_size = {{6'd0}, _T_95}; // @[StreamController.scala 48:25:@14983.4]
  assign io_dram_rresp_ready = rdata_io_in_ready; // @[StreamController.scala 55:23:@15028.4]
  assign io_load_cmd_ready = cmd_io_in_ready; // @[StreamController.scala 42:21:@14977.4]
  assign io_load_data_valid = rdata_io_out_valid; // @[StreamController.scala 57:22:@15029.4]
  assign io_load_data_bits_rdata_0 = rdata_io_out_bits_data_0; // @[StreamController.scala 58:27:@15030.4]
  assign cmd_clock = clock; // @[:@14580.4]
  assign cmd_reset = reset; // @[:@14581.4]
  assign cmd_io_in_valid = io_load_cmd_valid; // @[StreamController.scala 40:19:@14974.4]
  assign cmd_io_in_bits_addr = io_load_cmd_bits_addr; // @[StreamController.scala 41:18:@14976.4]
  assign cmd_io_in_bits_size = io_load_cmd_bits_size; // @[StreamController.scala 41:18:@14975.4]
  assign cmd_io_out_ready = io_dram_cmd_ready; // @[StreamController.scala 43:20:@14978.4]
  assign rdata_clock = clock; // @[:@14986.4]
  assign rdata_reset = reset; // @[:@14987.4]
  assign rdata_io_in_valid = io_dram_rresp_valid; // @[StreamController.scala 54:21:@15027.4]
  assign rdata_io_in_bits_data_0 = io_dram_rresp_bits_rdata_0; // @[StreamController.scala 53:25:@15011.4]
  assign rdata_io_in_bits_data_1 = io_dram_rresp_bits_rdata_1; // @[StreamController.scala 53:25:@15012.4]
  assign rdata_io_in_bits_data_2 = io_dram_rresp_bits_rdata_2; // @[StreamController.scala 53:25:@15013.4]
  assign rdata_io_in_bits_data_3 = io_dram_rresp_bits_rdata_3; // @[StreamController.scala 53:25:@15014.4]
  assign rdata_io_in_bits_data_4 = io_dram_rresp_bits_rdata_4; // @[StreamController.scala 53:25:@15015.4]
  assign rdata_io_in_bits_data_5 = io_dram_rresp_bits_rdata_5; // @[StreamController.scala 53:25:@15016.4]
  assign rdata_io_in_bits_data_6 = io_dram_rresp_bits_rdata_6; // @[StreamController.scala 53:25:@15017.4]
  assign rdata_io_in_bits_data_7 = io_dram_rresp_bits_rdata_7; // @[StreamController.scala 53:25:@15018.4]
  assign rdata_io_in_bits_data_8 = io_dram_rresp_bits_rdata_8; // @[StreamController.scala 53:25:@15019.4]
  assign rdata_io_in_bits_data_9 = io_dram_rresp_bits_rdata_9; // @[StreamController.scala 53:25:@15020.4]
  assign rdata_io_in_bits_data_10 = io_dram_rresp_bits_rdata_10; // @[StreamController.scala 53:25:@15021.4]
  assign rdata_io_in_bits_data_11 = io_dram_rresp_bits_rdata_11; // @[StreamController.scala 53:25:@15022.4]
  assign rdata_io_in_bits_data_12 = io_dram_rresp_bits_rdata_12; // @[StreamController.scala 53:25:@15023.4]
  assign rdata_io_in_bits_data_13 = io_dram_rresp_bits_rdata_13; // @[StreamController.scala 53:25:@15024.4]
  assign rdata_io_in_bits_data_14 = io_dram_rresp_bits_rdata_14; // @[StreamController.scala 53:25:@15025.4]
  assign rdata_io_in_bits_data_15 = io_dram_rresp_bits_rdata_15; // @[StreamController.scala 53:25:@15026.4]
  assign rdata_io_out_ready = io_load_data_ready; // @[StreamController.scala 59:22:@15031.4]
endmodule
module MuxPipe( // @[:@15097.2]
  output        io_in_ready, // @[:@15100.4]
  input         io_in_valid, // @[:@15100.4]
  input  [63:0] io_in_bits_0_addr, // @[:@15100.4]
  input  [31:0] io_in_bits_0_size, // @[:@15100.4]
  input         io_out_ready, // @[:@15100.4]
  output        io_out_valid, // @[:@15100.4]
  output [63:0] io_out_bits_addr, // @[:@15100.4]
  output [31:0] io_out_bits_size // @[:@15100.4]
);
  wire  _T_42; // @[MuxN.scala 28:31:@15102.4]
  assign _T_42 = io_out_valid == 1'h0; // @[MuxN.scala 28:31:@15102.4]
  assign io_in_ready = io_out_ready | _T_42; // @[MuxN.scala 71:15:@15111.4]
  assign io_out_valid = io_in_valid; // @[MuxN.scala 70:16:@15110.4]
  assign io_out_bits_addr = io_in_bits_0_addr; // @[MuxN.scala 72:15:@15116.4]
  assign io_out_bits_size = io_in_bits_0_size; // @[MuxN.scala 72:15:@15115.4]
endmodule
module StreamArbiter( // @[:@15308.2]
  input         clock, // @[:@15309.4]
  input         reset, // @[:@15310.4]
  output        io_app_0_cmd_ready, // @[:@15311.4]
  input         io_app_0_cmd_valid, // @[:@15311.4]
  input  [63:0] io_app_0_cmd_bits_addr, // @[:@15311.4]
  input  [31:0] io_app_0_cmd_bits_size, // @[:@15311.4]
  input         io_app_0_rresp_ready, // @[:@15311.4]
  output        io_app_0_rresp_valid, // @[:@15311.4]
  output [31:0] io_app_0_rresp_bits_rdata_0, // @[:@15311.4]
  output [31:0] io_app_0_rresp_bits_rdata_1, // @[:@15311.4]
  output [31:0] io_app_0_rresp_bits_rdata_2, // @[:@15311.4]
  output [31:0] io_app_0_rresp_bits_rdata_3, // @[:@15311.4]
  output [31:0] io_app_0_rresp_bits_rdata_4, // @[:@15311.4]
  output [31:0] io_app_0_rresp_bits_rdata_5, // @[:@15311.4]
  output [31:0] io_app_0_rresp_bits_rdata_6, // @[:@15311.4]
  output [31:0] io_app_0_rresp_bits_rdata_7, // @[:@15311.4]
  output [31:0] io_app_0_rresp_bits_rdata_8, // @[:@15311.4]
  output [31:0] io_app_0_rresp_bits_rdata_9, // @[:@15311.4]
  output [31:0] io_app_0_rresp_bits_rdata_10, // @[:@15311.4]
  output [31:0] io_app_0_rresp_bits_rdata_11, // @[:@15311.4]
  output [31:0] io_app_0_rresp_bits_rdata_12, // @[:@15311.4]
  output [31:0] io_app_0_rresp_bits_rdata_13, // @[:@15311.4]
  output [31:0] io_app_0_rresp_bits_rdata_14, // @[:@15311.4]
  output [31:0] io_app_0_rresp_bits_rdata_15, // @[:@15311.4]
  input         io_dram_cmd_ready, // @[:@15311.4]
  output        io_dram_cmd_valid, // @[:@15311.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@15311.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@15311.4]
  output        io_dram_rresp_ready, // @[:@15311.4]
  input         io_dram_rresp_valid, // @[:@15311.4]
  input  [31:0] io_dram_rresp_bits_rdata_0, // @[:@15311.4]
  input  [31:0] io_dram_rresp_bits_rdata_1, // @[:@15311.4]
  input  [31:0] io_dram_rresp_bits_rdata_2, // @[:@15311.4]
  input  [31:0] io_dram_rresp_bits_rdata_3, // @[:@15311.4]
  input  [31:0] io_dram_rresp_bits_rdata_4, // @[:@15311.4]
  input  [31:0] io_dram_rresp_bits_rdata_5, // @[:@15311.4]
  input  [31:0] io_dram_rresp_bits_rdata_6, // @[:@15311.4]
  input  [31:0] io_dram_rresp_bits_rdata_7, // @[:@15311.4]
  input  [31:0] io_dram_rresp_bits_rdata_8, // @[:@15311.4]
  input  [31:0] io_dram_rresp_bits_rdata_9, // @[:@15311.4]
  input  [31:0] io_dram_rresp_bits_rdata_10, // @[:@15311.4]
  input  [31:0] io_dram_rresp_bits_rdata_11, // @[:@15311.4]
  input  [31:0] io_dram_rresp_bits_rdata_12, // @[:@15311.4]
  input  [31:0] io_dram_rresp_bits_rdata_13, // @[:@15311.4]
  input  [31:0] io_dram_rresp_bits_rdata_14, // @[:@15311.4]
  input  [31:0] io_dram_rresp_bits_rdata_15, // @[:@15311.4]
  input  [31:0] io_dram_rresp_bits_tag // @[:@15311.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@15540.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@15540.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@15540.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@15540.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@15540.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@15547.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@15547.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@15547.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@15547.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@15547.4]
  wire  cmdMux_io_in_ready; // @[StreamArbiter.scala 25:22:@15557.4]
  wire  cmdMux_io_in_valid; // @[StreamArbiter.scala 25:22:@15557.4]
  wire [63:0] cmdMux_io_in_bits_0_addr; // @[StreamArbiter.scala 25:22:@15557.4]
  wire [31:0] cmdMux_io_in_bits_0_size; // @[StreamArbiter.scala 25:22:@15557.4]
  wire  cmdMux_io_out_ready; // @[StreamArbiter.scala 25:22:@15557.4]
  wire  cmdMux_io_out_valid; // @[StreamArbiter.scala 25:22:@15557.4]
  wire [63:0] cmdMux_io_out_bits_addr; // @[StreamArbiter.scala 25:22:@15557.4]
  wire [31:0] cmdMux_io_out_bits_size; // @[StreamArbiter.scala 25:22:@15557.4]
  wire  _T_346; // @[package.scala 96:25:@15552.4 package.scala 96:25:@15553.4]
  wire  cmdIdx; // @[StreamArbiter.scala 21:16:@15554.4]
  wire [1:0] cmdInDecoder; // @[OneHot.scala 45:35:@15556.4]
  wire [7:0] _T_387; // @[FringeBundles.scala 132:28:@15780.4]
  wire [255:0] rrespDecoder; // @[OneHot.scala 45:35:@15795.4]
  wire  _T_400; // @[StreamArbiter.scala 61:55:@15801.4]
  wire  _T_407; // @[StreamArbiter.scala 64:58:@15810.4]
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@15540.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@15547.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  MuxPipe cmdMux ( // @[StreamArbiter.scala 25:22:@15557.4]
    .io_in_ready(cmdMux_io_in_ready),
    .io_in_valid(cmdMux_io_in_valid),
    .io_in_bits_0_addr(cmdMux_io_in_bits_0_addr),
    .io_in_bits_0_size(cmdMux_io_in_bits_0_size),
    .io_out_ready(cmdMux_io_out_ready),
    .io_out_valid(cmdMux_io_out_valid),
    .io_out_bits_addr(cmdMux_io_out_bits_addr),
    .io_out_bits_size(cmdMux_io_out_bits_size)
  );
  assign _T_346 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@15552.4 package.scala 96:25:@15553.4]
  assign cmdIdx = io_app_0_cmd_valid ? _T_346 : 1'h0; // @[StreamArbiter.scala 21:16:@15554.4]
  assign cmdInDecoder = 2'h1 << cmdIdx; // @[OneHot.scala 45:35:@15556.4]
  assign _T_387 = io_dram_rresp_bits_tag[7:0]; // @[FringeBundles.scala 132:28:@15780.4]
  assign rrespDecoder = 256'h1 << _T_387; // @[OneHot.scala 45:35:@15795.4]
  assign _T_400 = cmdInDecoder[0]; // @[StreamArbiter.scala 61:55:@15801.4]
  assign _T_407 = rrespDecoder[0]; // @[StreamArbiter.scala 64:58:@15810.4]
  assign io_app_0_cmd_ready = cmdMux_io_in_ready & _T_400; // @[StreamArbiter.scala 61:19:@15803.4]
  assign io_app_0_rresp_valid = io_dram_rresp_valid & _T_407; // @[StreamArbiter.scala 64:21:@15812.4]
  assign io_app_0_rresp_bits_rdata_0 = io_dram_rresp_bits_rdata_0; // @[StreamArbiter.scala 65:20:@15814.4]
  assign io_app_0_rresp_bits_rdata_1 = io_dram_rresp_bits_rdata_1; // @[StreamArbiter.scala 65:20:@15815.4]
  assign io_app_0_rresp_bits_rdata_2 = io_dram_rresp_bits_rdata_2; // @[StreamArbiter.scala 65:20:@15816.4]
  assign io_app_0_rresp_bits_rdata_3 = io_dram_rresp_bits_rdata_3; // @[StreamArbiter.scala 65:20:@15817.4]
  assign io_app_0_rresp_bits_rdata_4 = io_dram_rresp_bits_rdata_4; // @[StreamArbiter.scala 65:20:@15818.4]
  assign io_app_0_rresp_bits_rdata_5 = io_dram_rresp_bits_rdata_5; // @[StreamArbiter.scala 65:20:@15819.4]
  assign io_app_0_rresp_bits_rdata_6 = io_dram_rresp_bits_rdata_6; // @[StreamArbiter.scala 65:20:@15820.4]
  assign io_app_0_rresp_bits_rdata_7 = io_dram_rresp_bits_rdata_7; // @[StreamArbiter.scala 65:20:@15821.4]
  assign io_app_0_rresp_bits_rdata_8 = io_dram_rresp_bits_rdata_8; // @[StreamArbiter.scala 65:20:@15822.4]
  assign io_app_0_rresp_bits_rdata_9 = io_dram_rresp_bits_rdata_9; // @[StreamArbiter.scala 65:20:@15823.4]
  assign io_app_0_rresp_bits_rdata_10 = io_dram_rresp_bits_rdata_10; // @[StreamArbiter.scala 65:20:@15824.4]
  assign io_app_0_rresp_bits_rdata_11 = io_dram_rresp_bits_rdata_11; // @[StreamArbiter.scala 65:20:@15825.4]
  assign io_app_0_rresp_bits_rdata_12 = io_dram_rresp_bits_rdata_12; // @[StreamArbiter.scala 65:20:@15826.4]
  assign io_app_0_rresp_bits_rdata_13 = io_dram_rresp_bits_rdata_13; // @[StreamArbiter.scala 65:20:@15827.4]
  assign io_app_0_rresp_bits_rdata_14 = io_dram_rresp_bits_rdata_14; // @[StreamArbiter.scala 65:20:@15828.4]
  assign io_app_0_rresp_bits_rdata_15 = io_dram_rresp_bits_rdata_15; // @[StreamArbiter.scala 65:20:@15829.4]
  assign io_dram_cmd_valid = cmdMux_io_out_valid; // @[StreamArbiter.scala 46:15:@15692.4]
  assign io_dram_cmd_bits_addr = cmdMux_io_out_bits_addr; // @[StreamArbiter.scala 46:15:@15691.4]
  assign io_dram_cmd_bits_size = cmdMux_io_out_bits_size; // @[StreamArbiter.scala 46:15:@15690.4]
  assign io_dram_rresp_ready = io_app_0_rresp_ready; // @[StreamArbiter.scala 72:23:@15836.4]
  assign RetimeWrapper_clock = clock; // @[:@15541.4]
  assign RetimeWrapper_reset = reset; // @[:@15542.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@15544.4]
  assign RetimeWrapper_io_in = io_app_0_cmd_valid ? _T_346 : 1'h0; // @[package.scala 94:16:@15543.4]
  assign RetimeWrapper_1_clock = clock; // @[:@15548.4]
  assign RetimeWrapper_1_reset = reset; // @[:@15549.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@15551.4]
  assign RetimeWrapper_1_io_in = io_app_0_cmd_valid ? _T_346 : 1'h0; // @[package.scala 94:16:@15550.4]
  assign cmdMux_io_in_valid = io_app_0_cmd_valid; // @[StreamArbiter.scala 26:22:@15560.4]
  assign cmdMux_io_in_bits_0_addr = io_app_0_cmd_bits_addr; // @[StreamArbiter.scala 29:9:@15566.4]
  assign cmdMux_io_in_bits_0_size = io_app_0_cmd_bits_size; // @[StreamArbiter.scala 29:9:@15565.4]
  assign cmdMux_io_out_ready = io_dram_cmd_valid & io_dram_cmd_ready; // @[StreamArbiter.scala 46:15:@15693.4 StreamArbiter.scala 57:23:@15799.4]
endmodule
module Counter_40( // @[:@15841.2]
  input         clock, // @[:@15842.4]
  input         reset, // @[:@15843.4]
  input         io_reset, // @[:@15844.4]
  input         io_enable, // @[:@15844.4]
  input  [31:0] io_stride, // @[:@15844.4]
  output [31:0] io_out, // @[:@15844.4]
  output [31:0] io_next // @[:@15844.4]
);
  reg [31:0] count; // @[Counter.scala 15:22:@15846.4]
  reg [31:0] _RAND_0;
  wire [32:0] _T_17; // @[Counter.scala 17:24:@15847.4]
  wire [31:0] newCount; // @[Counter.scala 17:24:@15848.4]
  wire [31:0] _GEN_0; // @[Counter.scala 21:26:@15853.6]
  wire [31:0] _GEN_1; // @[Counter.scala 19:18:@15849.4]
  assign _T_17 = count + io_stride; // @[Counter.scala 17:24:@15847.4]
  assign newCount = count + io_stride; // @[Counter.scala 17:24:@15848.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@15853.6]
  assign _GEN_1 = io_reset ? 32'h0 : _GEN_0; // @[Counter.scala 19:18:@15849.4]
  assign io_out = count; // @[Counter.scala 25:10:@15856.4]
  assign io_next = count + io_stride; // @[Counter.scala 26:11:@15857.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 32'h0;
    end else begin
      if (io_reset) begin
        count <= 32'h0;
      end else begin
        if (io_enable) begin
          count <= newCount;
        end
      end
    end
  end
endmodule
module AXICmdSplit( // @[:@15859.2]
  input         clock, // @[:@15860.4]
  input         reset, // @[:@15861.4]
  output        io_in_cmd_ready, // @[:@15862.4]
  input         io_in_cmd_valid, // @[:@15862.4]
  input  [63:0] io_in_cmd_bits_addr, // @[:@15862.4]
  input  [31:0] io_in_cmd_bits_size, // @[:@15862.4]
  input         io_in_rresp_ready, // @[:@15862.4]
  output        io_in_rresp_valid, // @[:@15862.4]
  output [31:0] io_in_rresp_bits_rdata_0, // @[:@15862.4]
  output [31:0] io_in_rresp_bits_rdata_1, // @[:@15862.4]
  output [31:0] io_in_rresp_bits_rdata_2, // @[:@15862.4]
  output [31:0] io_in_rresp_bits_rdata_3, // @[:@15862.4]
  output [31:0] io_in_rresp_bits_rdata_4, // @[:@15862.4]
  output [31:0] io_in_rresp_bits_rdata_5, // @[:@15862.4]
  output [31:0] io_in_rresp_bits_rdata_6, // @[:@15862.4]
  output [31:0] io_in_rresp_bits_rdata_7, // @[:@15862.4]
  output [31:0] io_in_rresp_bits_rdata_8, // @[:@15862.4]
  output [31:0] io_in_rresp_bits_rdata_9, // @[:@15862.4]
  output [31:0] io_in_rresp_bits_rdata_10, // @[:@15862.4]
  output [31:0] io_in_rresp_bits_rdata_11, // @[:@15862.4]
  output [31:0] io_in_rresp_bits_rdata_12, // @[:@15862.4]
  output [31:0] io_in_rresp_bits_rdata_13, // @[:@15862.4]
  output [31:0] io_in_rresp_bits_rdata_14, // @[:@15862.4]
  output [31:0] io_in_rresp_bits_rdata_15, // @[:@15862.4]
  output [31:0] io_in_rresp_bits_tag, // @[:@15862.4]
  input         io_out_cmd_ready, // @[:@15862.4]
  output        io_out_cmd_valid, // @[:@15862.4]
  output [63:0] io_out_cmd_bits_addr, // @[:@15862.4]
  output [31:0] io_out_cmd_bits_size, // @[:@15862.4]
  output [31:0] io_out_cmd_bits_tag, // @[:@15862.4]
  output        io_out_rresp_ready, // @[:@15862.4]
  input         io_out_rresp_valid, // @[:@15862.4]
  input  [31:0] io_out_rresp_bits_rdata_0, // @[:@15862.4]
  input  [31:0] io_out_rresp_bits_rdata_1, // @[:@15862.4]
  input  [31:0] io_out_rresp_bits_rdata_2, // @[:@15862.4]
  input  [31:0] io_out_rresp_bits_rdata_3, // @[:@15862.4]
  input  [31:0] io_out_rresp_bits_rdata_4, // @[:@15862.4]
  input  [31:0] io_out_rresp_bits_rdata_5, // @[:@15862.4]
  input  [31:0] io_out_rresp_bits_rdata_6, // @[:@15862.4]
  input  [31:0] io_out_rresp_bits_rdata_7, // @[:@15862.4]
  input  [31:0] io_out_rresp_bits_rdata_8, // @[:@15862.4]
  input  [31:0] io_out_rresp_bits_rdata_9, // @[:@15862.4]
  input  [31:0] io_out_rresp_bits_rdata_10, // @[:@15862.4]
  input  [31:0] io_out_rresp_bits_rdata_11, // @[:@15862.4]
  input  [31:0] io_out_rresp_bits_rdata_12, // @[:@15862.4]
  input  [31:0] io_out_rresp_bits_rdata_13, // @[:@15862.4]
  input  [31:0] io_out_rresp_bits_rdata_14, // @[:@15862.4]
  input  [31:0] io_out_rresp_bits_rdata_15, // @[:@15862.4]
  input  [31:0] io_out_rresp_bits_tag, // @[:@15862.4]
  output        io_out_wresp_ready, // @[:@15862.4]
  input  [31:0] io_out_wresp_bits_tag // @[:@15862.4]
);
  wire  cmdSizeCounter_clock; // @[AXIProtocol.scala 18:30:@15976.4]
  wire  cmdSizeCounter_reset; // @[AXIProtocol.scala 18:30:@15976.4]
  wire  cmdSizeCounter_io_reset; // @[AXIProtocol.scala 18:30:@15976.4]
  wire  cmdSizeCounter_io_enable; // @[AXIProtocol.scala 18:30:@15976.4]
  wire [31:0] cmdSizeCounter_io_stride; // @[AXIProtocol.scala 18:30:@15976.4]
  wire [31:0] cmdSizeCounter_io_out; // @[AXIProtocol.scala 18:30:@15976.4]
  wire [31:0] cmdSizeCounter_io_next; // @[AXIProtocol.scala 18:30:@15976.4]
  wire [32:0] _T_199; // @[AXIProtocol.scala 20:46:@15979.4]
  wire [32:0] _T_200; // @[AXIProtocol.scala 20:46:@15980.4]
  wire [31:0] cmdSizeRemaining; // @[AXIProtocol.scala 20:46:@15981.4]
  wire  lastCmd; // @[AXIProtocol.scala 23:35:@15982.4]
  wire [37:0] _GEN_0; // @[AXIProtocol.scala 27:47:@15985.4]
  wire [37:0] addrOffsetBytes; // @[AXIProtocol.scala 27:47:@15985.4]
  wire [63:0] _GEN_1; // @[AXIProtocol.scala 28:49:@15986.4]
  wire [64:0] _T_201; // @[AXIProtocol.scala 28:49:@15986.4]
  wire [63:0] cmdAddr_bits; // @[AXIProtocol.scala 28:49:@15987.4]
  wire [57:0] _T_204; // @[FringeBundles.scala 158:22:@15990.4]
  wire [23:0] _T_214; // @[FringeBundles.scala 115:37:@16004.4]
  wire  cmdIssue; // @[AXIProtocol.scala 36:35:@16007.4]
  wire  _T_223; // @[FringeBundles.scala 140:28:@16018.4]
  Counter_40 cmdSizeCounter ( // @[AXIProtocol.scala 18:30:@15976.4]
    .clock(cmdSizeCounter_clock),
    .reset(cmdSizeCounter_reset),
    .io_reset(cmdSizeCounter_io_reset),
    .io_enable(cmdSizeCounter_io_enable),
    .io_stride(cmdSizeCounter_io_stride),
    .io_out(cmdSizeCounter_io_out),
    .io_next(cmdSizeCounter_io_next)
  );
  assign _T_199 = io_in_cmd_bits_size - cmdSizeCounter_io_out; // @[AXIProtocol.scala 20:46:@15979.4]
  assign _T_200 = $unsigned(_T_199); // @[AXIProtocol.scala 20:46:@15980.4]
  assign cmdSizeRemaining = _T_200[31:0]; // @[AXIProtocol.scala 20:46:@15981.4]
  assign lastCmd = cmdSizeRemaining <= 32'h100; // @[AXIProtocol.scala 23:35:@15982.4]
  assign _GEN_0 = {{6'd0}, cmdSizeCounter_io_out}; // @[AXIProtocol.scala 27:47:@15985.4]
  assign addrOffsetBytes = _GEN_0 << 6; // @[AXIProtocol.scala 27:47:@15985.4]
  assign _GEN_1 = {{26'd0}, addrOffsetBytes}; // @[AXIProtocol.scala 28:49:@15986.4]
  assign _T_201 = io_in_cmd_bits_addr + _GEN_1; // @[AXIProtocol.scala 28:49:@15986.4]
  assign cmdAddr_bits = io_in_cmd_bits_addr + _GEN_1; // @[AXIProtocol.scala 28:49:@15987.4]
  assign _T_204 = cmdAddr_bits[63:6]; // @[FringeBundles.scala 158:22:@15990.4]
  assign _T_214 = {23'h0,lastCmd}; // @[FringeBundles.scala 115:37:@16004.4]
  assign cmdIssue = io_out_cmd_valid & io_out_cmd_ready; // @[AXIProtocol.scala 36:35:@16007.4]
  assign _T_223 = io_out_wresp_bits_tag[8]; // @[FringeBundles.scala 140:28:@16018.4]
  assign io_in_cmd_ready = lastCmd & cmdIssue; // @[AXIProtocol.scala 15:10:@15975.4 AXIProtocol.scala 38:19:@16009.4]
  assign io_in_rresp_valid = io_out_rresp_valid; // @[AXIProtocol.scala 15:10:@15884.4]
  assign io_in_rresp_bits_rdata_0 = io_out_rresp_bits_rdata_0; // @[AXIProtocol.scala 15:10:@15868.4]
  assign io_in_rresp_bits_rdata_1 = io_out_rresp_bits_rdata_1; // @[AXIProtocol.scala 15:10:@15869.4]
  assign io_in_rresp_bits_rdata_2 = io_out_rresp_bits_rdata_2; // @[AXIProtocol.scala 15:10:@15870.4]
  assign io_in_rresp_bits_rdata_3 = io_out_rresp_bits_rdata_3; // @[AXIProtocol.scala 15:10:@15871.4]
  assign io_in_rresp_bits_rdata_4 = io_out_rresp_bits_rdata_4; // @[AXIProtocol.scala 15:10:@15872.4]
  assign io_in_rresp_bits_rdata_5 = io_out_rresp_bits_rdata_5; // @[AXIProtocol.scala 15:10:@15873.4]
  assign io_in_rresp_bits_rdata_6 = io_out_rresp_bits_rdata_6; // @[AXIProtocol.scala 15:10:@15874.4]
  assign io_in_rresp_bits_rdata_7 = io_out_rresp_bits_rdata_7; // @[AXIProtocol.scala 15:10:@15875.4]
  assign io_in_rresp_bits_rdata_8 = io_out_rresp_bits_rdata_8; // @[AXIProtocol.scala 15:10:@15876.4]
  assign io_in_rresp_bits_rdata_9 = io_out_rresp_bits_rdata_9; // @[AXIProtocol.scala 15:10:@15877.4]
  assign io_in_rresp_bits_rdata_10 = io_out_rresp_bits_rdata_10; // @[AXIProtocol.scala 15:10:@15878.4]
  assign io_in_rresp_bits_rdata_11 = io_out_rresp_bits_rdata_11; // @[AXIProtocol.scala 15:10:@15879.4]
  assign io_in_rresp_bits_rdata_12 = io_out_rresp_bits_rdata_12; // @[AXIProtocol.scala 15:10:@15880.4]
  assign io_in_rresp_bits_rdata_13 = io_out_rresp_bits_rdata_13; // @[AXIProtocol.scala 15:10:@15881.4]
  assign io_in_rresp_bits_rdata_14 = io_out_rresp_bits_rdata_14; // @[AXIProtocol.scala 15:10:@15882.4]
  assign io_in_rresp_bits_rdata_15 = io_out_rresp_bits_rdata_15; // @[AXIProtocol.scala 15:10:@15883.4]
  assign io_in_rresp_bits_tag = io_out_rresp_bits_tag; // @[AXIProtocol.scala 15:10:@15867.4]
  assign io_out_cmd_valid = io_in_cmd_valid; // @[AXIProtocol.scala 15:10:@15974.4]
  assign io_out_cmd_bits_addr = {_T_204,6'h0}; // @[AXIProtocol.scala 15:10:@15973.4 AXIProtocol.scala 29:24:@15992.4]
  assign io_out_cmd_bits_size = lastCmd ? cmdSizeRemaining : 32'h100; // @[AXIProtocol.scala 15:10:@15972.4 AXIProtocol.scala 25:24:@15984.4]
  assign io_out_cmd_bits_tag = {_T_214,8'h0}; // @[AXIProtocol.scala 15:10:@15969.4 FringeBundles.scala 115:32:@16006.4]
  assign io_out_rresp_ready = io_in_rresp_ready; // @[AXIProtocol.scala 15:10:@15885.4]
  assign io_out_wresp_ready = _T_223 ? 1'h0 : 1'h1; // @[AXIProtocol.scala 15:10:@15866.4 AXIProtocol.scala 47:22:@16025.4]
  assign cmdSizeCounter_clock = clock; // @[:@15977.4]
  assign cmdSizeCounter_reset = reset; // @[:@15978.4]
  assign cmdSizeCounter_io_reset = lastCmd & cmdIssue; // @[AXIProtocol.scala 40:27:@16010.4]
  assign cmdSizeCounter_io_enable = io_out_cmd_valid & io_out_cmd_ready; // @[AXIProtocol.scala 41:28:@16011.4]
  assign cmdSizeCounter_io_stride = 32'h100; // @[AXIProtocol.scala 42:28:@16012.4]
endmodule
module AXICmdIssue( // @[:@16045.2]
  input         clock, // @[:@16046.4]
  input         reset, // @[:@16047.4]
  output        io_in_cmd_ready, // @[:@16048.4]
  input         io_in_cmd_valid, // @[:@16048.4]
  input  [63:0] io_in_cmd_bits_addr, // @[:@16048.4]
  input  [31:0] io_in_cmd_bits_size, // @[:@16048.4]
  input  [31:0] io_in_cmd_bits_tag, // @[:@16048.4]
  input         io_in_rresp_ready, // @[:@16048.4]
  output        io_in_rresp_valid, // @[:@16048.4]
  output [31:0] io_in_rresp_bits_rdata_0, // @[:@16048.4]
  output [31:0] io_in_rresp_bits_rdata_1, // @[:@16048.4]
  output [31:0] io_in_rresp_bits_rdata_2, // @[:@16048.4]
  output [31:0] io_in_rresp_bits_rdata_3, // @[:@16048.4]
  output [31:0] io_in_rresp_bits_rdata_4, // @[:@16048.4]
  output [31:0] io_in_rresp_bits_rdata_5, // @[:@16048.4]
  output [31:0] io_in_rresp_bits_rdata_6, // @[:@16048.4]
  output [31:0] io_in_rresp_bits_rdata_7, // @[:@16048.4]
  output [31:0] io_in_rresp_bits_rdata_8, // @[:@16048.4]
  output [31:0] io_in_rresp_bits_rdata_9, // @[:@16048.4]
  output [31:0] io_in_rresp_bits_rdata_10, // @[:@16048.4]
  output [31:0] io_in_rresp_bits_rdata_11, // @[:@16048.4]
  output [31:0] io_in_rresp_bits_rdata_12, // @[:@16048.4]
  output [31:0] io_in_rresp_bits_rdata_13, // @[:@16048.4]
  output [31:0] io_in_rresp_bits_rdata_14, // @[:@16048.4]
  output [31:0] io_in_rresp_bits_rdata_15, // @[:@16048.4]
  output [31:0] io_in_rresp_bits_tag, // @[:@16048.4]
  input         io_in_wresp_ready, // @[:@16048.4]
  output [31:0] io_in_wresp_bits_tag, // @[:@16048.4]
  input         io_out_cmd_ready, // @[:@16048.4]
  output        io_out_cmd_valid, // @[:@16048.4]
  output [63:0] io_out_cmd_bits_addr, // @[:@16048.4]
  output [31:0] io_out_cmd_bits_size, // @[:@16048.4]
  output [31:0] io_out_cmd_bits_tag, // @[:@16048.4]
  input         io_out_wdata_ready, // @[:@16048.4]
  output        io_out_wdata_valid, // @[:@16048.4]
  output        io_out_wdata_bits_wlast, // @[:@16048.4]
  output        io_out_rresp_ready, // @[:@16048.4]
  input         io_out_rresp_valid, // @[:@16048.4]
  input  [31:0] io_out_rresp_bits_rdata_0, // @[:@16048.4]
  input  [31:0] io_out_rresp_bits_rdata_1, // @[:@16048.4]
  input  [31:0] io_out_rresp_bits_rdata_2, // @[:@16048.4]
  input  [31:0] io_out_rresp_bits_rdata_3, // @[:@16048.4]
  input  [31:0] io_out_rresp_bits_rdata_4, // @[:@16048.4]
  input  [31:0] io_out_rresp_bits_rdata_5, // @[:@16048.4]
  input  [31:0] io_out_rresp_bits_rdata_6, // @[:@16048.4]
  input  [31:0] io_out_rresp_bits_rdata_7, // @[:@16048.4]
  input  [31:0] io_out_rresp_bits_rdata_8, // @[:@16048.4]
  input  [31:0] io_out_rresp_bits_rdata_9, // @[:@16048.4]
  input  [31:0] io_out_rresp_bits_rdata_10, // @[:@16048.4]
  input  [31:0] io_out_rresp_bits_rdata_11, // @[:@16048.4]
  input  [31:0] io_out_rresp_bits_rdata_12, // @[:@16048.4]
  input  [31:0] io_out_rresp_bits_rdata_13, // @[:@16048.4]
  input  [31:0] io_out_rresp_bits_rdata_14, // @[:@16048.4]
  input  [31:0] io_out_rresp_bits_rdata_15, // @[:@16048.4]
  input  [31:0] io_out_rresp_bits_tag, // @[:@16048.4]
  output        io_out_wresp_ready, // @[:@16048.4]
  input  [31:0] io_out_wresp_bits_tag // @[:@16048.4]
);
  wire  wdataCounter_clock; // @[AXIProtocol.scala 59:28:@16162.4]
  wire  wdataCounter_reset; // @[AXIProtocol.scala 59:28:@16162.4]
  wire  wdataCounter_io_reset; // @[AXIProtocol.scala 59:28:@16162.4]
  wire  wdataCounter_io_enable; // @[AXIProtocol.scala 59:28:@16162.4]
  wire [31:0] wdataCounter_io_stride; // @[AXIProtocol.scala 59:28:@16162.4]
  wire [31:0] wdataCounter_io_out; // @[AXIProtocol.scala 59:28:@16162.4]
  wire [31:0] wdataCounter_io_next; // @[AXIProtocol.scala 59:28:@16162.4]
  wire  dramWriteIssue; // @[AXIProtocol.scala 64:43:@16167.4]
  wire  _T_201; // @[AXIProtocol.scala 68:54:@16168.4]
  Counter_40 wdataCounter ( // @[AXIProtocol.scala 59:28:@16162.4]
    .clock(wdataCounter_clock),
    .reset(wdataCounter_reset),
    .io_reset(wdataCounter_io_reset),
    .io_enable(wdataCounter_io_enable),
    .io_stride(wdataCounter_io_stride),
    .io_out(wdataCounter_io_out),
    .io_next(wdataCounter_io_next)
  );
  assign dramWriteIssue = io_out_wdata_valid & io_out_wdata_ready; // @[AXIProtocol.scala 64:43:@16167.4]
  assign _T_201 = wdataCounter_io_next == io_in_cmd_bits_size; // @[AXIProtocol.scala 68:54:@16168.4]
  assign io_in_cmd_ready = io_out_cmd_valid & io_out_cmd_ready; // @[AXIProtocol.scala 56:10:@16161.4 AXIProtocol.scala 81:19:@16183.4]
  assign io_in_rresp_valid = io_out_rresp_valid; // @[AXIProtocol.scala 56:10:@16070.4]
  assign io_in_rresp_bits_rdata_0 = io_out_rresp_bits_rdata_0; // @[AXIProtocol.scala 56:10:@16054.4]
  assign io_in_rresp_bits_rdata_1 = io_out_rresp_bits_rdata_1; // @[AXIProtocol.scala 56:10:@16055.4]
  assign io_in_rresp_bits_rdata_2 = io_out_rresp_bits_rdata_2; // @[AXIProtocol.scala 56:10:@16056.4]
  assign io_in_rresp_bits_rdata_3 = io_out_rresp_bits_rdata_3; // @[AXIProtocol.scala 56:10:@16057.4]
  assign io_in_rresp_bits_rdata_4 = io_out_rresp_bits_rdata_4; // @[AXIProtocol.scala 56:10:@16058.4]
  assign io_in_rresp_bits_rdata_5 = io_out_rresp_bits_rdata_5; // @[AXIProtocol.scala 56:10:@16059.4]
  assign io_in_rresp_bits_rdata_6 = io_out_rresp_bits_rdata_6; // @[AXIProtocol.scala 56:10:@16060.4]
  assign io_in_rresp_bits_rdata_7 = io_out_rresp_bits_rdata_7; // @[AXIProtocol.scala 56:10:@16061.4]
  assign io_in_rresp_bits_rdata_8 = io_out_rresp_bits_rdata_8; // @[AXIProtocol.scala 56:10:@16062.4]
  assign io_in_rresp_bits_rdata_9 = io_out_rresp_bits_rdata_9; // @[AXIProtocol.scala 56:10:@16063.4]
  assign io_in_rresp_bits_rdata_10 = io_out_rresp_bits_rdata_10; // @[AXIProtocol.scala 56:10:@16064.4]
  assign io_in_rresp_bits_rdata_11 = io_out_rresp_bits_rdata_11; // @[AXIProtocol.scala 56:10:@16065.4]
  assign io_in_rresp_bits_rdata_12 = io_out_rresp_bits_rdata_12; // @[AXIProtocol.scala 56:10:@16066.4]
  assign io_in_rresp_bits_rdata_13 = io_out_rresp_bits_rdata_13; // @[AXIProtocol.scala 56:10:@16067.4]
  assign io_in_rresp_bits_rdata_14 = io_out_rresp_bits_rdata_14; // @[AXIProtocol.scala 56:10:@16068.4]
  assign io_in_rresp_bits_rdata_15 = io_out_rresp_bits_rdata_15; // @[AXIProtocol.scala 56:10:@16069.4]
  assign io_in_rresp_bits_tag = io_out_rresp_bits_tag; // @[AXIProtocol.scala 56:10:@16053.4]
  assign io_in_wresp_bits_tag = io_out_wresp_bits_tag; // @[AXIProtocol.scala 56:10:@16050.4]
  assign io_out_cmd_valid = io_in_cmd_valid; // @[AXIProtocol.scala 56:10:@16160.4 AXIProtocol.scala 84:20:@16188.4]
  assign io_out_cmd_bits_addr = io_in_cmd_bits_addr; // @[AXIProtocol.scala 56:10:@16159.4]
  assign io_out_cmd_bits_size = io_in_cmd_bits_size; // @[AXIProtocol.scala 56:10:@16158.4]
  assign io_out_cmd_bits_tag = io_in_cmd_bits_tag; // @[AXIProtocol.scala 56:10:@16155.4]
  assign io_out_wdata_valid = 1'h0; // @[AXIProtocol.scala 56:10:@16153.4 AXIProtocol.scala 86:22:@16190.4]
  assign io_out_wdata_bits_wlast = dramWriteIssue & _T_201; // @[AXIProtocol.scala 56:10:@16072.4 AXIProtocol.scala 87:27:@16191.4]
  assign io_out_rresp_ready = io_in_rresp_ready; // @[AXIProtocol.scala 56:10:@16071.4]
  assign io_out_wresp_ready = io_in_wresp_ready; // @[AXIProtocol.scala 56:10:@16052.4]
  assign wdataCounter_clock = clock; // @[:@16163.4]
  assign wdataCounter_reset = reset; // @[:@16164.4]
  assign wdataCounter_io_reset = dramWriteIssue & _T_201; // @[AXIProtocol.scala 76:25:@16179.4]
  assign wdataCounter_io_enable = io_out_wdata_valid & io_out_wdata_ready; // @[AXIProtocol.scala 77:26:@16180.4]
  assign wdataCounter_io_stride = 32'h1; // @[AXIProtocol.scala 78:26:@16181.4]
endmodule
module DRAMArbiter( // @[:@16193.2]
  input         clock, // @[:@16194.4]
  input         reset, // @[:@16195.4]
  input         io_enable, // @[:@16196.4]
  output        io_app_loads_0_cmd_ready, // @[:@16196.4]
  input         io_app_loads_0_cmd_valid, // @[:@16196.4]
  input  [63:0] io_app_loads_0_cmd_bits_addr, // @[:@16196.4]
  input  [31:0] io_app_loads_0_cmd_bits_size, // @[:@16196.4]
  input         io_app_loads_0_data_ready, // @[:@16196.4]
  output        io_app_loads_0_data_valid, // @[:@16196.4]
  output [31:0] io_app_loads_0_data_bits_rdata_0, // @[:@16196.4]
  output        io_app_stores_0_cmd_ready, // @[:@16196.4]
  input         io_app_stores_0_cmd_valid, // @[:@16196.4]
  input  [63:0] io_app_stores_0_cmd_bits_addr, // @[:@16196.4]
  input  [31:0] io_app_stores_0_cmd_bits_size, // @[:@16196.4]
  output        io_app_stores_0_data_ready, // @[:@16196.4]
  input         io_app_stores_0_data_valid, // @[:@16196.4]
  input  [31:0] io_app_stores_0_data_bits_wdata_0, // @[:@16196.4]
  input  [15:0] io_app_stores_0_data_bits_wstrb, // @[:@16196.4]
  input         io_dram_cmd_ready, // @[:@16196.4]
  output        io_dram_cmd_valid, // @[:@16196.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@16196.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@16196.4]
  output        io_dram_cmd_bits_isWr, // @[:@16196.4]
  output [31:0] io_dram_cmd_bits_tag, // @[:@16196.4]
  input         io_dram_wdata_ready, // @[:@16196.4]
  output        io_dram_wdata_valid, // @[:@16196.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@16196.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@16196.4]
  output        io_dram_wdata_bits_wlast, // @[:@16196.4]
  output        io_dram_rresp_ready, // @[:@16196.4]
  input         io_dram_rresp_valid, // @[:@16196.4]
  input  [31:0] io_dram_rresp_bits_rdata_0, // @[:@16196.4]
  input  [31:0] io_dram_rresp_bits_rdata_1, // @[:@16196.4]
  input  [31:0] io_dram_rresp_bits_rdata_2, // @[:@16196.4]
  input  [31:0] io_dram_rresp_bits_rdata_3, // @[:@16196.4]
  input  [31:0] io_dram_rresp_bits_rdata_4, // @[:@16196.4]
  input  [31:0] io_dram_rresp_bits_rdata_5, // @[:@16196.4]
  input  [31:0] io_dram_rresp_bits_rdata_6, // @[:@16196.4]
  input  [31:0] io_dram_rresp_bits_rdata_7, // @[:@16196.4]
  input  [31:0] io_dram_rresp_bits_rdata_8, // @[:@16196.4]
  input  [31:0] io_dram_rresp_bits_rdata_9, // @[:@16196.4]
  input  [31:0] io_dram_rresp_bits_rdata_10, // @[:@16196.4]
  input  [31:0] io_dram_rresp_bits_rdata_11, // @[:@16196.4]
  input  [31:0] io_dram_rresp_bits_rdata_12, // @[:@16196.4]
  input  [31:0] io_dram_rresp_bits_rdata_13, // @[:@16196.4]
  input  [31:0] io_dram_rresp_bits_rdata_14, // @[:@16196.4]
  input  [31:0] io_dram_rresp_bits_rdata_15, // @[:@16196.4]
  input  [31:0] io_dram_rresp_bits_tag, // @[:@16196.4]
  output        io_dram_wresp_ready, // @[:@16196.4]
  input         io_dram_wresp_valid, // @[:@16196.4]
  input  [31:0] io_dram_wresp_bits_tag, // @[:@16196.4]
  output [31:0] io_debugSignals_0, // @[:@16196.4]
  output [31:0] io_debugSignals_1, // @[:@16196.4]
  output [31:0] io_debugSignals_2, // @[:@16196.4]
  output [31:0] io_debugSignals_3, // @[:@16196.4]
  output [31:0] io_debugSignals_4, // @[:@16196.4]
  output [31:0] io_debugSignals_5, // @[:@16196.4]
  output [31:0] io_debugSignals_6, // @[:@16196.4]
  output [31:0] io_debugSignals_7, // @[:@16196.4]
  output [31:0] io_debugSignals_8, // @[:@16196.4]
  output [31:0] io_debugSignals_9, // @[:@16196.4]
  output [31:0] io_debugSignals_10, // @[:@16196.4]
  output [31:0] io_debugSignals_11, // @[:@16196.4]
  output [31:0] io_debugSignals_12, // @[:@16196.4]
  output [31:0] io_debugSignals_13, // @[:@16196.4]
  output [31:0] io_debugSignals_14, // @[:@16196.4]
  output [31:0] io_debugSignals_15, // @[:@16196.4]
  output [31:0] io_debugSignals_16, // @[:@16196.4]
  output [31:0] io_debugSignals_17, // @[:@16196.4]
  output [31:0] io_debugSignals_18, // @[:@16196.4]
  output [31:0] io_debugSignals_19, // @[:@16196.4]
  output [31:0] io_debugSignals_20, // @[:@16196.4]
  output [31:0] io_debugSignals_21, // @[:@16196.4]
  output [31:0] io_debugSignals_22, // @[:@16196.4]
  output [31:0] io_debugSignals_23, // @[:@16196.4]
  output [31:0] io_debugSignals_24, // @[:@16196.4]
  output [31:0] io_debugSignals_25, // @[:@16196.4]
  output [31:0] io_debugSignals_26, // @[:@16196.4]
  output [31:0] io_debugSignals_27, // @[:@16196.4]
  output [31:0] io_debugSignals_28, // @[:@16196.4]
  output [31:0] io_debugSignals_29, // @[:@16196.4]
  output [31:0] io_debugSignals_40 // @[:@16196.4]
);
  wire  StreamControllerLoad_clock; // @[DRAMArbiter.scala 60:21:@17082.4]
  wire  StreamControllerLoad_reset; // @[DRAMArbiter.scala 60:21:@17082.4]
  wire  StreamControllerLoad_io_dram_cmd_ready; // @[DRAMArbiter.scala 60:21:@17082.4]
  wire  StreamControllerLoad_io_dram_cmd_valid; // @[DRAMArbiter.scala 60:21:@17082.4]
  wire [63:0] StreamControllerLoad_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 60:21:@17082.4]
  wire [31:0] StreamControllerLoad_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 60:21:@17082.4]
  wire  StreamControllerLoad_io_dram_rresp_ready; // @[DRAMArbiter.scala 60:21:@17082.4]
  wire  StreamControllerLoad_io_dram_rresp_valid; // @[DRAMArbiter.scala 60:21:@17082.4]
  wire [31:0] StreamControllerLoad_io_dram_rresp_bits_rdata_0; // @[DRAMArbiter.scala 60:21:@17082.4]
  wire [31:0] StreamControllerLoad_io_dram_rresp_bits_rdata_1; // @[DRAMArbiter.scala 60:21:@17082.4]
  wire [31:0] StreamControllerLoad_io_dram_rresp_bits_rdata_2; // @[DRAMArbiter.scala 60:21:@17082.4]
  wire [31:0] StreamControllerLoad_io_dram_rresp_bits_rdata_3; // @[DRAMArbiter.scala 60:21:@17082.4]
  wire [31:0] StreamControllerLoad_io_dram_rresp_bits_rdata_4; // @[DRAMArbiter.scala 60:21:@17082.4]
  wire [31:0] StreamControllerLoad_io_dram_rresp_bits_rdata_5; // @[DRAMArbiter.scala 60:21:@17082.4]
  wire [31:0] StreamControllerLoad_io_dram_rresp_bits_rdata_6; // @[DRAMArbiter.scala 60:21:@17082.4]
  wire [31:0] StreamControllerLoad_io_dram_rresp_bits_rdata_7; // @[DRAMArbiter.scala 60:21:@17082.4]
  wire [31:0] StreamControllerLoad_io_dram_rresp_bits_rdata_8; // @[DRAMArbiter.scala 60:21:@17082.4]
  wire [31:0] StreamControllerLoad_io_dram_rresp_bits_rdata_9; // @[DRAMArbiter.scala 60:21:@17082.4]
  wire [31:0] StreamControllerLoad_io_dram_rresp_bits_rdata_10; // @[DRAMArbiter.scala 60:21:@17082.4]
  wire [31:0] StreamControllerLoad_io_dram_rresp_bits_rdata_11; // @[DRAMArbiter.scala 60:21:@17082.4]
  wire [31:0] StreamControllerLoad_io_dram_rresp_bits_rdata_12; // @[DRAMArbiter.scala 60:21:@17082.4]
  wire [31:0] StreamControllerLoad_io_dram_rresp_bits_rdata_13; // @[DRAMArbiter.scala 60:21:@17082.4]
  wire [31:0] StreamControllerLoad_io_dram_rresp_bits_rdata_14; // @[DRAMArbiter.scala 60:21:@17082.4]
  wire [31:0] StreamControllerLoad_io_dram_rresp_bits_rdata_15; // @[DRAMArbiter.scala 60:21:@17082.4]
  wire  StreamControllerLoad_io_load_cmd_ready; // @[DRAMArbiter.scala 60:21:@17082.4]
  wire  StreamControllerLoad_io_load_cmd_valid; // @[DRAMArbiter.scala 60:21:@17082.4]
  wire [63:0] StreamControllerLoad_io_load_cmd_bits_addr; // @[DRAMArbiter.scala 60:21:@17082.4]
  wire [31:0] StreamControllerLoad_io_load_cmd_bits_size; // @[DRAMArbiter.scala 60:21:@17082.4]
  wire  StreamControllerLoad_io_load_data_ready; // @[DRAMArbiter.scala 60:21:@17082.4]
  wire  StreamControllerLoad_io_load_data_valid; // @[DRAMArbiter.scala 60:21:@17082.4]
  wire [31:0] StreamControllerLoad_io_load_data_bits_rdata_0; // @[DRAMArbiter.scala 60:21:@17082.4]
  wire  StreamArbiter_clock; // @[DRAMArbiter.scala 86:27:@17092.4]
  wire  StreamArbiter_reset; // @[DRAMArbiter.scala 86:27:@17092.4]
  wire  StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 86:27:@17092.4]
  wire  StreamArbiter_io_app_0_cmd_valid; // @[DRAMArbiter.scala 86:27:@17092.4]
  wire [63:0] StreamArbiter_io_app_0_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@17092.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@17092.4]
  wire  StreamArbiter_io_app_0_rresp_ready; // @[DRAMArbiter.scala 86:27:@17092.4]
  wire  StreamArbiter_io_app_0_rresp_valid; // @[DRAMArbiter.scala 86:27:@17092.4]
  wire [31:0] StreamArbiter_io_app_0_rresp_bits_rdata_0; // @[DRAMArbiter.scala 86:27:@17092.4]
  wire [31:0] StreamArbiter_io_app_0_rresp_bits_rdata_1; // @[DRAMArbiter.scala 86:27:@17092.4]
  wire [31:0] StreamArbiter_io_app_0_rresp_bits_rdata_2; // @[DRAMArbiter.scala 86:27:@17092.4]
  wire [31:0] StreamArbiter_io_app_0_rresp_bits_rdata_3; // @[DRAMArbiter.scala 86:27:@17092.4]
  wire [31:0] StreamArbiter_io_app_0_rresp_bits_rdata_4; // @[DRAMArbiter.scala 86:27:@17092.4]
  wire [31:0] StreamArbiter_io_app_0_rresp_bits_rdata_5; // @[DRAMArbiter.scala 86:27:@17092.4]
  wire [31:0] StreamArbiter_io_app_0_rresp_bits_rdata_6; // @[DRAMArbiter.scala 86:27:@17092.4]
  wire [31:0] StreamArbiter_io_app_0_rresp_bits_rdata_7; // @[DRAMArbiter.scala 86:27:@17092.4]
  wire [31:0] StreamArbiter_io_app_0_rresp_bits_rdata_8; // @[DRAMArbiter.scala 86:27:@17092.4]
  wire [31:0] StreamArbiter_io_app_0_rresp_bits_rdata_9; // @[DRAMArbiter.scala 86:27:@17092.4]
  wire [31:0] StreamArbiter_io_app_0_rresp_bits_rdata_10; // @[DRAMArbiter.scala 86:27:@17092.4]
  wire [31:0] StreamArbiter_io_app_0_rresp_bits_rdata_11; // @[DRAMArbiter.scala 86:27:@17092.4]
  wire [31:0] StreamArbiter_io_app_0_rresp_bits_rdata_12; // @[DRAMArbiter.scala 86:27:@17092.4]
  wire [31:0] StreamArbiter_io_app_0_rresp_bits_rdata_13; // @[DRAMArbiter.scala 86:27:@17092.4]
  wire [31:0] StreamArbiter_io_app_0_rresp_bits_rdata_14; // @[DRAMArbiter.scala 86:27:@17092.4]
  wire [31:0] StreamArbiter_io_app_0_rresp_bits_rdata_15; // @[DRAMArbiter.scala 86:27:@17092.4]
  wire  StreamArbiter_io_dram_cmd_ready; // @[DRAMArbiter.scala 86:27:@17092.4]
  wire  StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 86:27:@17092.4]
  wire [63:0] StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@17092.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@17092.4]
  wire  StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 86:27:@17092.4]
  wire  StreamArbiter_io_dram_rresp_valid; // @[DRAMArbiter.scala 86:27:@17092.4]
  wire [31:0] StreamArbiter_io_dram_rresp_bits_rdata_0; // @[DRAMArbiter.scala 86:27:@17092.4]
  wire [31:0] StreamArbiter_io_dram_rresp_bits_rdata_1; // @[DRAMArbiter.scala 86:27:@17092.4]
  wire [31:0] StreamArbiter_io_dram_rresp_bits_rdata_2; // @[DRAMArbiter.scala 86:27:@17092.4]
  wire [31:0] StreamArbiter_io_dram_rresp_bits_rdata_3; // @[DRAMArbiter.scala 86:27:@17092.4]
  wire [31:0] StreamArbiter_io_dram_rresp_bits_rdata_4; // @[DRAMArbiter.scala 86:27:@17092.4]
  wire [31:0] StreamArbiter_io_dram_rresp_bits_rdata_5; // @[DRAMArbiter.scala 86:27:@17092.4]
  wire [31:0] StreamArbiter_io_dram_rresp_bits_rdata_6; // @[DRAMArbiter.scala 86:27:@17092.4]
  wire [31:0] StreamArbiter_io_dram_rresp_bits_rdata_7; // @[DRAMArbiter.scala 86:27:@17092.4]
  wire [31:0] StreamArbiter_io_dram_rresp_bits_rdata_8; // @[DRAMArbiter.scala 86:27:@17092.4]
  wire [31:0] StreamArbiter_io_dram_rresp_bits_rdata_9; // @[DRAMArbiter.scala 86:27:@17092.4]
  wire [31:0] StreamArbiter_io_dram_rresp_bits_rdata_10; // @[DRAMArbiter.scala 86:27:@17092.4]
  wire [31:0] StreamArbiter_io_dram_rresp_bits_rdata_11; // @[DRAMArbiter.scala 86:27:@17092.4]
  wire [31:0] StreamArbiter_io_dram_rresp_bits_rdata_12; // @[DRAMArbiter.scala 86:27:@17092.4]
  wire [31:0] StreamArbiter_io_dram_rresp_bits_rdata_13; // @[DRAMArbiter.scala 86:27:@17092.4]
  wire [31:0] StreamArbiter_io_dram_rresp_bits_rdata_14; // @[DRAMArbiter.scala 86:27:@17092.4]
  wire [31:0] StreamArbiter_io_dram_rresp_bits_rdata_15; // @[DRAMArbiter.scala 86:27:@17092.4]
  wire [31:0] StreamArbiter_io_dram_rresp_bits_tag; // @[DRAMArbiter.scala 86:27:@17092.4]
  wire  AXICmdSplit_clock; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire  AXICmdSplit_reset; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire  AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire  AXICmdSplit_io_in_cmd_valid; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire [63:0] AXICmdSplit_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire  AXICmdSplit_io_in_rresp_ready; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire  AXICmdSplit_io_in_rresp_valid; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire [31:0] AXICmdSplit_io_in_rresp_bits_rdata_0; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire [31:0] AXICmdSplit_io_in_rresp_bits_rdata_1; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire [31:0] AXICmdSplit_io_in_rresp_bits_rdata_2; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire [31:0] AXICmdSplit_io_in_rresp_bits_rdata_3; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire [31:0] AXICmdSplit_io_in_rresp_bits_rdata_4; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire [31:0] AXICmdSplit_io_in_rresp_bits_rdata_5; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire [31:0] AXICmdSplit_io_in_rresp_bits_rdata_6; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire [31:0] AXICmdSplit_io_in_rresp_bits_rdata_7; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire [31:0] AXICmdSplit_io_in_rresp_bits_rdata_8; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire [31:0] AXICmdSplit_io_in_rresp_bits_rdata_9; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire [31:0] AXICmdSplit_io_in_rresp_bits_rdata_10; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire [31:0] AXICmdSplit_io_in_rresp_bits_rdata_11; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire [31:0] AXICmdSplit_io_in_rresp_bits_rdata_12; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire [31:0] AXICmdSplit_io_in_rresp_bits_rdata_13; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire [31:0] AXICmdSplit_io_in_rresp_bits_rdata_14; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire [31:0] AXICmdSplit_io_in_rresp_bits_rdata_15; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire [31:0] AXICmdSplit_io_in_rresp_bits_tag; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire  AXICmdSplit_io_out_cmd_ready; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire  AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire [63:0] AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire  AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire  AXICmdSplit_io_out_rresp_valid; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire [31:0] AXICmdSplit_io_out_rresp_bits_rdata_0; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire [31:0] AXICmdSplit_io_out_rresp_bits_rdata_1; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire [31:0] AXICmdSplit_io_out_rresp_bits_rdata_2; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire [31:0] AXICmdSplit_io_out_rresp_bits_rdata_3; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire [31:0] AXICmdSplit_io_out_rresp_bits_rdata_4; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire [31:0] AXICmdSplit_io_out_rresp_bits_rdata_5; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire [31:0] AXICmdSplit_io_out_rresp_bits_rdata_6; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire [31:0] AXICmdSplit_io_out_rresp_bits_rdata_7; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire [31:0] AXICmdSplit_io_out_rresp_bits_rdata_8; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire [31:0] AXICmdSplit_io_out_rresp_bits_rdata_9; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire [31:0] AXICmdSplit_io_out_rresp_bits_rdata_10; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire [31:0] AXICmdSplit_io_out_rresp_bits_rdata_11; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire [31:0] AXICmdSplit_io_out_rresp_bits_rdata_12; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire [31:0] AXICmdSplit_io_out_rresp_bits_rdata_13; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire [31:0] AXICmdSplit_io_out_rresp_bits_rdata_14; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire [31:0] AXICmdSplit_io_out_rresp_bits_rdata_15; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire [31:0] AXICmdSplit_io_out_rresp_bits_tag; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire  AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire [31:0] AXICmdSplit_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@17320.4]
  wire  AXICmdIssue_clock; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire  AXICmdIssue_reset; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire  AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire  AXICmdIssue_io_in_cmd_valid; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire [63:0] AXICmdIssue_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire  AXICmdIssue_io_in_rresp_ready; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire  AXICmdIssue_io_in_rresp_valid; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire [31:0] AXICmdIssue_io_in_rresp_bits_rdata_0; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire [31:0] AXICmdIssue_io_in_rresp_bits_rdata_1; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire [31:0] AXICmdIssue_io_in_rresp_bits_rdata_2; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire [31:0] AXICmdIssue_io_in_rresp_bits_rdata_3; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire [31:0] AXICmdIssue_io_in_rresp_bits_rdata_4; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire [31:0] AXICmdIssue_io_in_rresp_bits_rdata_5; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire [31:0] AXICmdIssue_io_in_rresp_bits_rdata_6; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire [31:0] AXICmdIssue_io_in_rresp_bits_rdata_7; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire [31:0] AXICmdIssue_io_in_rresp_bits_rdata_8; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire [31:0] AXICmdIssue_io_in_rresp_bits_rdata_9; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire [31:0] AXICmdIssue_io_in_rresp_bits_rdata_10; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire [31:0] AXICmdIssue_io_in_rresp_bits_rdata_11; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire [31:0] AXICmdIssue_io_in_rresp_bits_rdata_12; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire [31:0] AXICmdIssue_io_in_rresp_bits_rdata_13; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire [31:0] AXICmdIssue_io_in_rresp_bits_rdata_14; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire [31:0] AXICmdIssue_io_in_rresp_bits_rdata_15; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire [31:0] AXICmdIssue_io_in_rresp_bits_tag; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire  AXICmdIssue_io_in_wresp_ready; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire [31:0] AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire  AXICmdIssue_io_out_cmd_ready; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire  AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire [63:0] AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire  AXICmdIssue_io_out_wdata_ready; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire  AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire  AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire  AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire  AXICmdIssue_io_out_rresp_valid; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire [31:0] AXICmdIssue_io_out_rresp_bits_rdata_0; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire [31:0] AXICmdIssue_io_out_rresp_bits_rdata_1; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire [31:0] AXICmdIssue_io_out_rresp_bits_rdata_2; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire [31:0] AXICmdIssue_io_out_rresp_bits_rdata_3; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire [31:0] AXICmdIssue_io_out_rresp_bits_rdata_4; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire [31:0] AXICmdIssue_io_out_rresp_bits_rdata_5; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire [31:0] AXICmdIssue_io_out_rresp_bits_rdata_6; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire [31:0] AXICmdIssue_io_out_rresp_bits_rdata_7; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire [31:0] AXICmdIssue_io_out_rresp_bits_rdata_8; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire [31:0] AXICmdIssue_io_out_rresp_bits_rdata_9; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire [31:0] AXICmdIssue_io_out_rresp_bits_rdata_10; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire [31:0] AXICmdIssue_io_out_rresp_bits_rdata_11; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire [31:0] AXICmdIssue_io_out_rresp_bits_rdata_12; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire [31:0] AXICmdIssue_io_out_rresp_bits_rdata_13; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire [31:0] AXICmdIssue_io_out_rresp_bits_rdata_14; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire [31:0] AXICmdIssue_io_out_rresp_bits_rdata_15; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire [31:0] AXICmdIssue_io_out_rresp_bits_tag; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire  AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 97:26:@17435.4]
  wire [31:0] AXICmdIssue_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@17435.4]
  reg [63:0] _T_1835; // @[DRAMArbiter.scala 119:24:@17666.4]
  reg [63:0] _RAND_0;
  wire [64:0] _T_1837; // @[DRAMArbiter.scala 121:18:@17668.6]
  wire [63:0] _T_1838; // @[DRAMArbiter.scala 121:18:@17669.6]
  wire [63:0] _GEN_0; // @[DRAMArbiter.scala 120:19:@17667.4]
  wire  _T_1839; // @[DRAMArbiter.scala 137:60:@17673.4]
  wire  _T_1846; // @[DRAMArbiter.scala 138:57:@17680.4]
  reg [63:0] _T_1849; // @[DRAMArbiter.scala 119:24:@17681.4]
  reg [63:0] _RAND_1;
  wire [64:0] _T_1851; // @[DRAMArbiter.scala 121:18:@17683.6]
  wire [63:0] _T_1852; // @[DRAMArbiter.scala 121:18:@17684.6]
  wire [63:0] _GEN_2; // @[DRAMArbiter.scala 120:19:@17682.4]
  wire  _T_1853; // @[DRAMArbiter.scala 139:70:@17687.4]
  reg [63:0] _T_1856; // @[DRAMArbiter.scala 119:24:@17688.4]
  reg [63:0] _RAND_2;
  wire [64:0] _T_1858; // @[DRAMArbiter.scala 121:18:@17690.6]
  wire [63:0] _T_1859; // @[DRAMArbiter.scala 121:18:@17691.6]
  wire [63:0] _GEN_3; // @[DRAMArbiter.scala 120:19:@17689.4]
  wire  _T_1860; // @[DRAMArbiter.scala 142:52:@17695.4]
  reg [63:0] _T_1863; // @[DRAMArbiter.scala 119:24:@17696.4]
  reg [63:0] _RAND_3;
  wire [64:0] _T_1865; // @[DRAMArbiter.scala 121:18:@17698.6]
  wire [63:0] _T_1866; // @[DRAMArbiter.scala 121:18:@17699.6]
  wire [63:0] _GEN_4; // @[DRAMArbiter.scala 120:19:@17697.4]
  wire  _T_1869; // @[DRAMArbiter.scala 143:74:@17704.4]
  wire  _T_1870; // @[DRAMArbiter.scala 143:72:@17705.4]
  reg [63:0] _T_1873; // @[DRAMArbiter.scala 119:24:@17706.4]
  reg [63:0] _RAND_4;
  wire [64:0] _T_1875; // @[DRAMArbiter.scala 121:18:@17708.6]
  wire [63:0] _T_1876; // @[DRAMArbiter.scala 121:18:@17709.6]
  wire [63:0] _GEN_5; // @[DRAMArbiter.scala 120:19:@17707.4]
  wire  _T_1878; // @[DRAMArbiter.scala 144:72:@17714.4]
  reg [63:0] _T_1881; // @[DRAMArbiter.scala 119:24:@17715.4]
  reg [63:0] _RAND_5;
  wire [64:0] _T_1883; // @[DRAMArbiter.scala 121:18:@17717.6]
  wire [63:0] _T_1884; // @[DRAMArbiter.scala 121:18:@17718.6]
  wire [63:0] _GEN_6; // @[DRAMArbiter.scala 120:19:@17716.4]
  wire  _T_1885; // @[DRAMArbiter.scala 148:59:@17722.4]
  wire  _T_1886; // @[DRAMArbiter.scala 148:76:@17723.4]
  reg [63:0] _T_1889; // @[DRAMArbiter.scala 119:24:@17724.4]
  reg [63:0] _RAND_6;
  wire [64:0] _T_1891; // @[DRAMArbiter.scala 121:18:@17726.6]
  wire [63:0] _T_1892; // @[DRAMArbiter.scala 121:18:@17727.6]
  wire [63:0] _GEN_7; // @[DRAMArbiter.scala 120:19:@17725.4]
  wire  _T_1893; // @[DRAMArbiter.scala 154:60:@17731.4]
  wire  _T_1894; // @[DRAMArbiter.scala 154:78:@17732.4]
  reg [63:0] _T_1897; // @[DRAMArbiter.scala 119:24:@17733.4]
  reg [63:0] _RAND_7;
  wire [64:0] _T_1899; // @[DRAMArbiter.scala 121:18:@17735.6]
  wire [63:0] _T_1900; // @[DRAMArbiter.scala 121:18:@17736.6]
  wire [63:0] _GEN_8; // @[DRAMArbiter.scala 120:19:@17734.4]
  reg [63:0] _T_1904; // @[DRAMArbiter.scala 119:24:@17741.4]
  reg [63:0] _RAND_8;
  wire [64:0] _T_1906; // @[DRAMArbiter.scala 121:18:@17743.6]
  wire [63:0] _T_1907; // @[DRAMArbiter.scala 121:18:@17744.6]
  wire [63:0] _GEN_9; // @[DRAMArbiter.scala 120:19:@17742.4]
  wire  _T_1909; // @[DRAMArbiter.scala 159:56:@17748.4]
  wire  _T_1910; // @[DRAMArbiter.scala 159:54:@17749.4]
  reg [63:0] _T_1913; // @[DRAMArbiter.scala 119:24:@17750.4]
  reg [63:0] _RAND_9;
  wire [64:0] _T_1915; // @[DRAMArbiter.scala 121:18:@17752.6]
  wire [63:0] _T_1916; // @[DRAMArbiter.scala 121:18:@17753.6]
  wire [63:0] _GEN_10; // @[DRAMArbiter.scala 120:19:@17751.4]
  wire  _T_1918; // @[DRAMArbiter.scala 160:34:@17757.4]
  wire  _T_1919; // @[DRAMArbiter.scala 160:55:@17758.4]
  reg [63:0] _T_1922; // @[DRAMArbiter.scala 119:24:@17759.4]
  reg [63:0] _RAND_10;
  wire [64:0] _T_1924; // @[DRAMArbiter.scala 121:18:@17761.6]
  wire [63:0] _T_1925; // @[DRAMArbiter.scala 121:18:@17762.6]
  wire [63:0] _GEN_11; // @[DRAMArbiter.scala 120:19:@17760.4]
  wire [7:0] _T_1932; // @[FringeBundles.scala 132:28:@17770.4]
  wire  _T_1936; // @[DRAMArbiter.scala 163:116:@17776.4]
  wire  _T_1937; // @[DRAMArbiter.scala 163:78:@17777.4]
  reg [63:0] _T_1940; // @[DRAMArbiter.scala 119:24:@17778.4]
  reg [63:0] _RAND_11;
  wire [64:0] _T_1942; // @[DRAMArbiter.scala 121:18:@17780.6]
  wire [63:0] _T_1943; // @[DRAMArbiter.scala 121:18:@17781.6]
  wire [63:0] _GEN_12; // @[DRAMArbiter.scala 120:19:@17779.4]
  wire  _T_1944; // @[DRAMArbiter.scala 165:54:@17785.4]
  reg [63:0] _T_1947; // @[DRAMArbiter.scala 119:24:@17786.4]
  reg [63:0] _RAND_12;
  wire [64:0] _T_1949; // @[DRAMArbiter.scala 121:18:@17788.6]
  wire [63:0] _T_1950; // @[DRAMArbiter.scala 121:18:@17789.6]
  wire [63:0] _GEN_13; // @[DRAMArbiter.scala 120:19:@17787.4]
  wire  _T_1952; // @[DRAMArbiter.scala 166:56:@17793.4]
  wire  _T_1953; // @[DRAMArbiter.scala 166:54:@17794.4]
  reg [63:0] _T_1956; // @[DRAMArbiter.scala 119:24:@17795.4]
  reg [63:0] _RAND_13;
  wire [64:0] _T_1958; // @[DRAMArbiter.scala 121:18:@17797.6]
  wire [63:0] _T_1959; // @[DRAMArbiter.scala 121:18:@17798.6]
  wire [63:0] _GEN_14; // @[DRAMArbiter.scala 120:19:@17796.4]
  wire  _T_1961; // @[DRAMArbiter.scala 167:34:@17802.4]
  wire  _T_1962; // @[DRAMArbiter.scala 167:55:@17803.4]
  reg [63:0] _T_1965; // @[DRAMArbiter.scala 119:24:@17804.4]
  reg [63:0] _RAND_14;
  wire [64:0] _T_1967; // @[DRAMArbiter.scala 121:18:@17806.6]
  wire [63:0] _T_1968; // @[DRAMArbiter.scala 121:18:@17807.6]
  wire [63:0] _GEN_15; // @[DRAMArbiter.scala 120:19:@17805.4]
  wire  _T_1969; // @[DRAMArbiter.scala 174:70:@17811.4]
  reg [63:0] _T_1971; // @[DRAMArbiter.scala 127:25:@17812.4]
  reg [63:0] _RAND_15;
  wire [63:0] _GEN_16; // @[DRAMArbiter.scala 128:19:@17813.4]
  reg [31:0] _T_1974; // @[DRAMArbiter.scala 127:25:@17818.4]
  reg [31:0] _RAND_16;
  wire [31:0] _GEN_17; // @[DRAMArbiter.scala 128:19:@17819.4]
  reg [31:0] _T_1977; // @[DRAMArbiter.scala 127:25:@17824.4]
  reg [31:0] _RAND_17;
  wire [31:0] _GEN_18; // @[DRAMArbiter.scala 128:19:@17825.4]
  reg  _T_1980; // @[DRAMArbiter.scala 127:25:@17830.4]
  reg [31:0] _RAND_18;
  wire  _GEN_19; // @[DRAMArbiter.scala 128:19:@17831.4]
  wire  _T_1983; // @[DRAMArbiter.scala 178:115:@17836.4]
  wire  _T_1984; // @[DRAMArbiter.scala 178:102:@17837.4]
  reg [31:0] _T_1986; // @[DRAMArbiter.scala 127:25:@17838.4]
  reg [31:0] _RAND_19;
  wire [31:0] _GEN_20; // @[DRAMArbiter.scala 128:19:@17839.4]
  reg  _T_1992; // @[DRAMArbiter.scala 127:25:@17846.4]
  reg [31:0] _RAND_20;
  wire  _GEN_21; // @[DRAMArbiter.scala 128:19:@17847.4]
  wire  _T_1995; // @[DRAMArbiter.scala 180:115:@17852.4]
  wire  _T_1996; // @[DRAMArbiter.scala 180:102:@17853.4]
  reg [31:0] _T_1998; // @[DRAMArbiter.scala 127:25:@17854.4]
  reg [31:0] _RAND_21;
  wire [31:0] _GEN_22; // @[DRAMArbiter.scala 128:19:@17855.4]
  reg  _T_2004; // @[DRAMArbiter.scala 127:25:@17862.4]
  reg [31:0] _RAND_22;
  wire  _GEN_23; // @[DRAMArbiter.scala 128:19:@17863.4]
  wire  _T_2005; // @[DRAMArbiter.scala 182:92:@17867.4]
  reg [63:0] _T_2007; // @[DRAMArbiter.scala 127:25:@17868.4]
  reg [63:0] _RAND_23;
  wire [63:0] _GEN_24; // @[DRAMArbiter.scala 128:19:@17869.4]
  reg [31:0] _T_2010; // @[DRAMArbiter.scala 127:25:@17874.4]
  reg [31:0] _RAND_24;
  wire [31:0] _GEN_25; // @[DRAMArbiter.scala 128:19:@17875.4]
  reg [31:0] _T_2013; // @[DRAMArbiter.scala 127:25:@17880.4]
  reg [31:0] _RAND_25;
  wire [31:0] _GEN_26; // @[DRAMArbiter.scala 128:19:@17881.4]
  reg [15:0] _T_2016; // @[DRAMArbiter.scala 127:25:@17886.4]
  reg [31:0] _RAND_26;
  wire [15:0] _GEN_27; // @[DRAMArbiter.scala 128:19:@17887.4]
  wire  _T_2019; // @[DRAMArbiter.scala 186:148:@17892.4]
  wire  _T_2020; // @[DRAMArbiter.scala 186:132:@17893.4]
  reg [31:0] _T_2022; // @[DRAMArbiter.scala 127:25:@17894.4]
  reg [31:0] _RAND_27;
  wire [31:0] _GEN_28; // @[DRAMArbiter.scala 128:19:@17895.4]
  reg [15:0] _T_2028; // @[DRAMArbiter.scala 127:25:@17902.4]
  reg [31:0] _RAND_28;
  wire [15:0] _GEN_29; // @[DRAMArbiter.scala 128:19:@17903.4]
  wire  _T_2031; // @[DRAMArbiter.scala 188:148:@17908.4]
  wire  _T_2032; // @[DRAMArbiter.scala 188:132:@17909.4]
  reg [31:0] _T_2034; // @[DRAMArbiter.scala 127:25:@17910.4]
  reg [31:0] _RAND_29;
  wire [31:0] _GEN_30; // @[DRAMArbiter.scala 128:19:@17911.4]
  reg [15:0] _T_2040; // @[DRAMArbiter.scala 127:25:@17918.4]
  reg [31:0] _RAND_30;
  wire [15:0] _GEN_31; // @[DRAMArbiter.scala 128:19:@17919.4]
  reg [63:0] _T_2112; // @[DRAMArbiter.scala 119:24:@18000.4]
  reg [63:0] _RAND_31;
  wire [64:0] _T_2114; // @[DRAMArbiter.scala 121:18:@18002.6]
  wire [63:0] _T_2115; // @[DRAMArbiter.scala 121:18:@18003.6]
  StreamControllerLoad StreamControllerLoad ( // @[DRAMArbiter.scala 60:21:@17082.4]
    .clock(StreamControllerLoad_clock),
    .reset(StreamControllerLoad_reset),
    .io_dram_cmd_ready(StreamControllerLoad_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamControllerLoad_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamControllerLoad_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamControllerLoad_io_dram_cmd_bits_size),
    .io_dram_rresp_ready(StreamControllerLoad_io_dram_rresp_ready),
    .io_dram_rresp_valid(StreamControllerLoad_io_dram_rresp_valid),
    .io_dram_rresp_bits_rdata_0(StreamControllerLoad_io_dram_rresp_bits_rdata_0),
    .io_dram_rresp_bits_rdata_1(StreamControllerLoad_io_dram_rresp_bits_rdata_1),
    .io_dram_rresp_bits_rdata_2(StreamControllerLoad_io_dram_rresp_bits_rdata_2),
    .io_dram_rresp_bits_rdata_3(StreamControllerLoad_io_dram_rresp_bits_rdata_3),
    .io_dram_rresp_bits_rdata_4(StreamControllerLoad_io_dram_rresp_bits_rdata_4),
    .io_dram_rresp_bits_rdata_5(StreamControllerLoad_io_dram_rresp_bits_rdata_5),
    .io_dram_rresp_bits_rdata_6(StreamControllerLoad_io_dram_rresp_bits_rdata_6),
    .io_dram_rresp_bits_rdata_7(StreamControllerLoad_io_dram_rresp_bits_rdata_7),
    .io_dram_rresp_bits_rdata_8(StreamControllerLoad_io_dram_rresp_bits_rdata_8),
    .io_dram_rresp_bits_rdata_9(StreamControllerLoad_io_dram_rresp_bits_rdata_9),
    .io_dram_rresp_bits_rdata_10(StreamControllerLoad_io_dram_rresp_bits_rdata_10),
    .io_dram_rresp_bits_rdata_11(StreamControllerLoad_io_dram_rresp_bits_rdata_11),
    .io_dram_rresp_bits_rdata_12(StreamControllerLoad_io_dram_rresp_bits_rdata_12),
    .io_dram_rresp_bits_rdata_13(StreamControllerLoad_io_dram_rresp_bits_rdata_13),
    .io_dram_rresp_bits_rdata_14(StreamControllerLoad_io_dram_rresp_bits_rdata_14),
    .io_dram_rresp_bits_rdata_15(StreamControllerLoad_io_dram_rresp_bits_rdata_15),
    .io_load_cmd_ready(StreamControllerLoad_io_load_cmd_ready),
    .io_load_cmd_valid(StreamControllerLoad_io_load_cmd_valid),
    .io_load_cmd_bits_addr(StreamControllerLoad_io_load_cmd_bits_addr),
    .io_load_cmd_bits_size(StreamControllerLoad_io_load_cmd_bits_size),
    .io_load_data_ready(StreamControllerLoad_io_load_data_ready),
    .io_load_data_valid(StreamControllerLoad_io_load_data_valid),
    .io_load_data_bits_rdata_0(StreamControllerLoad_io_load_data_bits_rdata_0)
  );
  StreamArbiter StreamArbiter ( // @[DRAMArbiter.scala 86:27:@17092.4]
    .clock(StreamArbiter_clock),
    .reset(StreamArbiter_reset),
    .io_app_0_cmd_ready(StreamArbiter_io_app_0_cmd_ready),
    .io_app_0_cmd_valid(StreamArbiter_io_app_0_cmd_valid),
    .io_app_0_cmd_bits_addr(StreamArbiter_io_app_0_cmd_bits_addr),
    .io_app_0_cmd_bits_size(StreamArbiter_io_app_0_cmd_bits_size),
    .io_app_0_rresp_ready(StreamArbiter_io_app_0_rresp_ready),
    .io_app_0_rresp_valid(StreamArbiter_io_app_0_rresp_valid),
    .io_app_0_rresp_bits_rdata_0(StreamArbiter_io_app_0_rresp_bits_rdata_0),
    .io_app_0_rresp_bits_rdata_1(StreamArbiter_io_app_0_rresp_bits_rdata_1),
    .io_app_0_rresp_bits_rdata_2(StreamArbiter_io_app_0_rresp_bits_rdata_2),
    .io_app_0_rresp_bits_rdata_3(StreamArbiter_io_app_0_rresp_bits_rdata_3),
    .io_app_0_rresp_bits_rdata_4(StreamArbiter_io_app_0_rresp_bits_rdata_4),
    .io_app_0_rresp_bits_rdata_5(StreamArbiter_io_app_0_rresp_bits_rdata_5),
    .io_app_0_rresp_bits_rdata_6(StreamArbiter_io_app_0_rresp_bits_rdata_6),
    .io_app_0_rresp_bits_rdata_7(StreamArbiter_io_app_0_rresp_bits_rdata_7),
    .io_app_0_rresp_bits_rdata_8(StreamArbiter_io_app_0_rresp_bits_rdata_8),
    .io_app_0_rresp_bits_rdata_9(StreamArbiter_io_app_0_rresp_bits_rdata_9),
    .io_app_0_rresp_bits_rdata_10(StreamArbiter_io_app_0_rresp_bits_rdata_10),
    .io_app_0_rresp_bits_rdata_11(StreamArbiter_io_app_0_rresp_bits_rdata_11),
    .io_app_0_rresp_bits_rdata_12(StreamArbiter_io_app_0_rresp_bits_rdata_12),
    .io_app_0_rresp_bits_rdata_13(StreamArbiter_io_app_0_rresp_bits_rdata_13),
    .io_app_0_rresp_bits_rdata_14(StreamArbiter_io_app_0_rresp_bits_rdata_14),
    .io_app_0_rresp_bits_rdata_15(StreamArbiter_io_app_0_rresp_bits_rdata_15),
    .io_dram_cmd_ready(StreamArbiter_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamArbiter_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamArbiter_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamArbiter_io_dram_cmd_bits_size),
    .io_dram_rresp_ready(StreamArbiter_io_dram_rresp_ready),
    .io_dram_rresp_valid(StreamArbiter_io_dram_rresp_valid),
    .io_dram_rresp_bits_rdata_0(StreamArbiter_io_dram_rresp_bits_rdata_0),
    .io_dram_rresp_bits_rdata_1(StreamArbiter_io_dram_rresp_bits_rdata_1),
    .io_dram_rresp_bits_rdata_2(StreamArbiter_io_dram_rresp_bits_rdata_2),
    .io_dram_rresp_bits_rdata_3(StreamArbiter_io_dram_rresp_bits_rdata_3),
    .io_dram_rresp_bits_rdata_4(StreamArbiter_io_dram_rresp_bits_rdata_4),
    .io_dram_rresp_bits_rdata_5(StreamArbiter_io_dram_rresp_bits_rdata_5),
    .io_dram_rresp_bits_rdata_6(StreamArbiter_io_dram_rresp_bits_rdata_6),
    .io_dram_rresp_bits_rdata_7(StreamArbiter_io_dram_rresp_bits_rdata_7),
    .io_dram_rresp_bits_rdata_8(StreamArbiter_io_dram_rresp_bits_rdata_8),
    .io_dram_rresp_bits_rdata_9(StreamArbiter_io_dram_rresp_bits_rdata_9),
    .io_dram_rresp_bits_rdata_10(StreamArbiter_io_dram_rresp_bits_rdata_10),
    .io_dram_rresp_bits_rdata_11(StreamArbiter_io_dram_rresp_bits_rdata_11),
    .io_dram_rresp_bits_rdata_12(StreamArbiter_io_dram_rresp_bits_rdata_12),
    .io_dram_rresp_bits_rdata_13(StreamArbiter_io_dram_rresp_bits_rdata_13),
    .io_dram_rresp_bits_rdata_14(StreamArbiter_io_dram_rresp_bits_rdata_14),
    .io_dram_rresp_bits_rdata_15(StreamArbiter_io_dram_rresp_bits_rdata_15),
    .io_dram_rresp_bits_tag(StreamArbiter_io_dram_rresp_bits_tag)
  );
  AXICmdSplit AXICmdSplit ( // @[DRAMArbiter.scala 94:26:@17320.4]
    .clock(AXICmdSplit_clock),
    .reset(AXICmdSplit_reset),
    .io_in_cmd_ready(AXICmdSplit_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdSplit_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdSplit_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdSplit_io_in_cmd_bits_size),
    .io_in_rresp_ready(AXICmdSplit_io_in_rresp_ready),
    .io_in_rresp_valid(AXICmdSplit_io_in_rresp_valid),
    .io_in_rresp_bits_rdata_0(AXICmdSplit_io_in_rresp_bits_rdata_0),
    .io_in_rresp_bits_rdata_1(AXICmdSplit_io_in_rresp_bits_rdata_1),
    .io_in_rresp_bits_rdata_2(AXICmdSplit_io_in_rresp_bits_rdata_2),
    .io_in_rresp_bits_rdata_3(AXICmdSplit_io_in_rresp_bits_rdata_3),
    .io_in_rresp_bits_rdata_4(AXICmdSplit_io_in_rresp_bits_rdata_4),
    .io_in_rresp_bits_rdata_5(AXICmdSplit_io_in_rresp_bits_rdata_5),
    .io_in_rresp_bits_rdata_6(AXICmdSplit_io_in_rresp_bits_rdata_6),
    .io_in_rresp_bits_rdata_7(AXICmdSplit_io_in_rresp_bits_rdata_7),
    .io_in_rresp_bits_rdata_8(AXICmdSplit_io_in_rresp_bits_rdata_8),
    .io_in_rresp_bits_rdata_9(AXICmdSplit_io_in_rresp_bits_rdata_9),
    .io_in_rresp_bits_rdata_10(AXICmdSplit_io_in_rresp_bits_rdata_10),
    .io_in_rresp_bits_rdata_11(AXICmdSplit_io_in_rresp_bits_rdata_11),
    .io_in_rresp_bits_rdata_12(AXICmdSplit_io_in_rresp_bits_rdata_12),
    .io_in_rresp_bits_rdata_13(AXICmdSplit_io_in_rresp_bits_rdata_13),
    .io_in_rresp_bits_rdata_14(AXICmdSplit_io_in_rresp_bits_rdata_14),
    .io_in_rresp_bits_rdata_15(AXICmdSplit_io_in_rresp_bits_rdata_15),
    .io_in_rresp_bits_tag(AXICmdSplit_io_in_rresp_bits_tag),
    .io_out_cmd_ready(AXICmdSplit_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdSplit_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdSplit_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdSplit_io_out_cmd_bits_size),
    .io_out_cmd_bits_tag(AXICmdSplit_io_out_cmd_bits_tag),
    .io_out_rresp_ready(AXICmdSplit_io_out_rresp_ready),
    .io_out_rresp_valid(AXICmdSplit_io_out_rresp_valid),
    .io_out_rresp_bits_rdata_0(AXICmdSplit_io_out_rresp_bits_rdata_0),
    .io_out_rresp_bits_rdata_1(AXICmdSplit_io_out_rresp_bits_rdata_1),
    .io_out_rresp_bits_rdata_2(AXICmdSplit_io_out_rresp_bits_rdata_2),
    .io_out_rresp_bits_rdata_3(AXICmdSplit_io_out_rresp_bits_rdata_3),
    .io_out_rresp_bits_rdata_4(AXICmdSplit_io_out_rresp_bits_rdata_4),
    .io_out_rresp_bits_rdata_5(AXICmdSplit_io_out_rresp_bits_rdata_5),
    .io_out_rresp_bits_rdata_6(AXICmdSplit_io_out_rresp_bits_rdata_6),
    .io_out_rresp_bits_rdata_7(AXICmdSplit_io_out_rresp_bits_rdata_7),
    .io_out_rresp_bits_rdata_8(AXICmdSplit_io_out_rresp_bits_rdata_8),
    .io_out_rresp_bits_rdata_9(AXICmdSplit_io_out_rresp_bits_rdata_9),
    .io_out_rresp_bits_rdata_10(AXICmdSplit_io_out_rresp_bits_rdata_10),
    .io_out_rresp_bits_rdata_11(AXICmdSplit_io_out_rresp_bits_rdata_11),
    .io_out_rresp_bits_rdata_12(AXICmdSplit_io_out_rresp_bits_rdata_12),
    .io_out_rresp_bits_rdata_13(AXICmdSplit_io_out_rresp_bits_rdata_13),
    .io_out_rresp_bits_rdata_14(AXICmdSplit_io_out_rresp_bits_rdata_14),
    .io_out_rresp_bits_rdata_15(AXICmdSplit_io_out_rresp_bits_rdata_15),
    .io_out_rresp_bits_tag(AXICmdSplit_io_out_rresp_bits_tag),
    .io_out_wresp_ready(AXICmdSplit_io_out_wresp_ready),
    .io_out_wresp_bits_tag(AXICmdSplit_io_out_wresp_bits_tag)
  );
  AXICmdIssue AXICmdIssue ( // @[DRAMArbiter.scala 97:26:@17435.4]
    .clock(AXICmdIssue_clock),
    .reset(AXICmdIssue_reset),
    .io_in_cmd_ready(AXICmdIssue_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdIssue_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdIssue_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdIssue_io_in_cmd_bits_size),
    .io_in_cmd_bits_tag(AXICmdIssue_io_in_cmd_bits_tag),
    .io_in_rresp_ready(AXICmdIssue_io_in_rresp_ready),
    .io_in_rresp_valid(AXICmdIssue_io_in_rresp_valid),
    .io_in_rresp_bits_rdata_0(AXICmdIssue_io_in_rresp_bits_rdata_0),
    .io_in_rresp_bits_rdata_1(AXICmdIssue_io_in_rresp_bits_rdata_1),
    .io_in_rresp_bits_rdata_2(AXICmdIssue_io_in_rresp_bits_rdata_2),
    .io_in_rresp_bits_rdata_3(AXICmdIssue_io_in_rresp_bits_rdata_3),
    .io_in_rresp_bits_rdata_4(AXICmdIssue_io_in_rresp_bits_rdata_4),
    .io_in_rresp_bits_rdata_5(AXICmdIssue_io_in_rresp_bits_rdata_5),
    .io_in_rresp_bits_rdata_6(AXICmdIssue_io_in_rresp_bits_rdata_6),
    .io_in_rresp_bits_rdata_7(AXICmdIssue_io_in_rresp_bits_rdata_7),
    .io_in_rresp_bits_rdata_8(AXICmdIssue_io_in_rresp_bits_rdata_8),
    .io_in_rresp_bits_rdata_9(AXICmdIssue_io_in_rresp_bits_rdata_9),
    .io_in_rresp_bits_rdata_10(AXICmdIssue_io_in_rresp_bits_rdata_10),
    .io_in_rresp_bits_rdata_11(AXICmdIssue_io_in_rresp_bits_rdata_11),
    .io_in_rresp_bits_rdata_12(AXICmdIssue_io_in_rresp_bits_rdata_12),
    .io_in_rresp_bits_rdata_13(AXICmdIssue_io_in_rresp_bits_rdata_13),
    .io_in_rresp_bits_rdata_14(AXICmdIssue_io_in_rresp_bits_rdata_14),
    .io_in_rresp_bits_rdata_15(AXICmdIssue_io_in_rresp_bits_rdata_15),
    .io_in_rresp_bits_tag(AXICmdIssue_io_in_rresp_bits_tag),
    .io_in_wresp_ready(AXICmdIssue_io_in_wresp_ready),
    .io_in_wresp_bits_tag(AXICmdIssue_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdIssue_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdIssue_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdIssue_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdIssue_io_out_cmd_bits_size),
    .io_out_cmd_bits_tag(AXICmdIssue_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdIssue_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdIssue_io_out_wdata_valid),
    .io_out_wdata_bits_wlast(AXICmdIssue_io_out_wdata_bits_wlast),
    .io_out_rresp_ready(AXICmdIssue_io_out_rresp_ready),
    .io_out_rresp_valid(AXICmdIssue_io_out_rresp_valid),
    .io_out_rresp_bits_rdata_0(AXICmdIssue_io_out_rresp_bits_rdata_0),
    .io_out_rresp_bits_rdata_1(AXICmdIssue_io_out_rresp_bits_rdata_1),
    .io_out_rresp_bits_rdata_2(AXICmdIssue_io_out_rresp_bits_rdata_2),
    .io_out_rresp_bits_rdata_3(AXICmdIssue_io_out_rresp_bits_rdata_3),
    .io_out_rresp_bits_rdata_4(AXICmdIssue_io_out_rresp_bits_rdata_4),
    .io_out_rresp_bits_rdata_5(AXICmdIssue_io_out_rresp_bits_rdata_5),
    .io_out_rresp_bits_rdata_6(AXICmdIssue_io_out_rresp_bits_rdata_6),
    .io_out_rresp_bits_rdata_7(AXICmdIssue_io_out_rresp_bits_rdata_7),
    .io_out_rresp_bits_rdata_8(AXICmdIssue_io_out_rresp_bits_rdata_8),
    .io_out_rresp_bits_rdata_9(AXICmdIssue_io_out_rresp_bits_rdata_9),
    .io_out_rresp_bits_rdata_10(AXICmdIssue_io_out_rresp_bits_rdata_10),
    .io_out_rresp_bits_rdata_11(AXICmdIssue_io_out_rresp_bits_rdata_11),
    .io_out_rresp_bits_rdata_12(AXICmdIssue_io_out_rresp_bits_rdata_12),
    .io_out_rresp_bits_rdata_13(AXICmdIssue_io_out_rresp_bits_rdata_13),
    .io_out_rresp_bits_rdata_14(AXICmdIssue_io_out_rresp_bits_rdata_14),
    .io_out_rresp_bits_rdata_15(AXICmdIssue_io_out_rresp_bits_rdata_15),
    .io_out_rresp_bits_tag(AXICmdIssue_io_out_rresp_bits_tag),
    .io_out_wresp_ready(AXICmdIssue_io_out_wresp_ready),
    .io_out_wresp_bits_tag(AXICmdIssue_io_out_wresp_bits_tag)
  );
  assign _T_1837 = _T_1835 + 64'h1; // @[DRAMArbiter.scala 121:18:@17668.6]
  assign _T_1838 = _T_1835 + 64'h1; // @[DRAMArbiter.scala 121:18:@17669.6]
  assign _GEN_0 = io_enable ? _T_1838 : _T_1835; // @[DRAMArbiter.scala 120:19:@17667.4]
  assign _T_1839 = io_dram_rresp_valid & io_dram_rresp_ready; // @[DRAMArbiter.scala 137:60:@17673.4]
  assign _T_1846 = io_dram_wdata_valid & io_dram_wdata_ready; // @[DRAMArbiter.scala 138:57:@17680.4]
  assign _T_1851 = _T_1849 + 64'h1; // @[DRAMArbiter.scala 121:18:@17683.6]
  assign _T_1852 = _T_1849 + 64'h1; // @[DRAMArbiter.scala 121:18:@17684.6]
  assign _GEN_2 = _T_1846 ? _T_1852 : _T_1849; // @[DRAMArbiter.scala 120:19:@17682.4]
  assign _T_1853 = io_app_stores_0_data_valid & io_app_stores_0_data_ready; // @[DRAMArbiter.scala 139:70:@17687.4]
  assign _T_1858 = _T_1856 + 64'h1; // @[DRAMArbiter.scala 121:18:@17690.6]
  assign _T_1859 = _T_1856 + 64'h1; // @[DRAMArbiter.scala 121:18:@17691.6]
  assign _GEN_3 = _T_1853 ? _T_1859 : _T_1856; // @[DRAMArbiter.scala 120:19:@17689.4]
  assign _T_1860 = io_dram_cmd_ready & io_dram_cmd_valid; // @[DRAMArbiter.scala 142:52:@17695.4]
  assign _T_1865 = _T_1863 + 64'h1; // @[DRAMArbiter.scala 121:18:@17698.6]
  assign _T_1866 = _T_1863 + 64'h1; // @[DRAMArbiter.scala 121:18:@17699.6]
  assign _GEN_4 = _T_1860 ? _T_1866 : _T_1863; // @[DRAMArbiter.scala 120:19:@17697.4]
  assign _T_1869 = io_dram_cmd_bits_isWr == 1'h0; // @[DRAMArbiter.scala 143:74:@17704.4]
  assign _T_1870 = _T_1860 & _T_1869; // @[DRAMArbiter.scala 143:72:@17705.4]
  assign _T_1875 = _T_1873 + 64'h1; // @[DRAMArbiter.scala 121:18:@17708.6]
  assign _T_1876 = _T_1873 + 64'h1; // @[DRAMArbiter.scala 121:18:@17709.6]
  assign _GEN_5 = _T_1870 ? _T_1876 : _T_1873; // @[DRAMArbiter.scala 120:19:@17707.4]
  assign _T_1878 = _T_1860 & io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 144:72:@17714.4]
  assign _T_1883 = _T_1881 + 64'h1; // @[DRAMArbiter.scala 121:18:@17717.6]
  assign _T_1884 = _T_1881 + 64'h1; // @[DRAMArbiter.scala 121:18:@17718.6]
  assign _GEN_6 = _T_1878 ? _T_1884 : _T_1881; // @[DRAMArbiter.scala 120:19:@17716.4]
  assign _T_1885 = io_enable & io_app_loads_0_cmd_valid; // @[DRAMArbiter.scala 148:59:@17722.4]
  assign _T_1886 = _T_1885 & io_app_loads_0_cmd_ready; // @[DRAMArbiter.scala 148:76:@17723.4]
  assign _T_1891 = _T_1889 + 64'h1; // @[DRAMArbiter.scala 121:18:@17726.6]
  assign _T_1892 = _T_1889 + 64'h1; // @[DRAMArbiter.scala 121:18:@17727.6]
  assign _GEN_7 = _T_1886 ? _T_1892 : _T_1889; // @[DRAMArbiter.scala 120:19:@17725.4]
  assign _T_1893 = io_enable & io_app_stores_0_cmd_valid; // @[DRAMArbiter.scala 154:60:@17731.4]
  assign _T_1894 = _T_1893 & io_app_stores_0_cmd_ready; // @[DRAMArbiter.scala 154:78:@17732.4]
  assign _T_1899 = _T_1897 + 64'h1; // @[DRAMArbiter.scala 121:18:@17735.6]
  assign _T_1900 = _T_1897 + 64'h1; // @[DRAMArbiter.scala 121:18:@17736.6]
  assign _GEN_8 = _T_1894 ? _T_1900 : _T_1897; // @[DRAMArbiter.scala 120:19:@17734.4]
  assign _T_1906 = _T_1904 + 64'h1; // @[DRAMArbiter.scala 121:18:@17743.6]
  assign _T_1907 = _T_1904 + 64'h1; // @[DRAMArbiter.scala 121:18:@17744.6]
  assign _GEN_9 = _T_1839 ? _T_1907 : _T_1904; // @[DRAMArbiter.scala 120:19:@17742.4]
  assign _T_1909 = io_dram_rresp_ready == 1'h0; // @[DRAMArbiter.scala 159:56:@17748.4]
  assign _T_1910 = io_dram_rresp_valid & _T_1909; // @[DRAMArbiter.scala 159:54:@17749.4]
  assign _T_1915 = _T_1913 + 64'h1; // @[DRAMArbiter.scala 121:18:@17752.6]
  assign _T_1916 = _T_1913 + 64'h1; // @[DRAMArbiter.scala 121:18:@17753.6]
  assign _GEN_10 = _T_1910 ? _T_1916 : _T_1913; // @[DRAMArbiter.scala 120:19:@17751.4]
  assign _T_1918 = io_dram_rresp_valid == 1'h0; // @[DRAMArbiter.scala 160:34:@17757.4]
  assign _T_1919 = _T_1918 & io_dram_rresp_ready; // @[DRAMArbiter.scala 160:55:@17758.4]
  assign _T_1924 = _T_1922 + 64'h1; // @[DRAMArbiter.scala 121:18:@17761.6]
  assign _T_1925 = _T_1922 + 64'h1; // @[DRAMArbiter.scala 121:18:@17762.6]
  assign _GEN_11 = _T_1919 ? _T_1925 : _T_1922; // @[DRAMArbiter.scala 120:19:@17760.4]
  assign _T_1932 = io_dram_rresp_bits_tag[7:0]; // @[FringeBundles.scala 132:28:@17770.4]
  assign _T_1936 = _T_1932 == 8'h0; // @[DRAMArbiter.scala 163:116:@17776.4]
  assign _T_1937 = _T_1839 & _T_1936; // @[DRAMArbiter.scala 163:78:@17777.4]
  assign _T_1942 = _T_1940 + 64'h1; // @[DRAMArbiter.scala 121:18:@17780.6]
  assign _T_1943 = _T_1940 + 64'h1; // @[DRAMArbiter.scala 121:18:@17781.6]
  assign _GEN_12 = _T_1937 ? _T_1943 : _T_1940; // @[DRAMArbiter.scala 120:19:@17779.4]
  assign _T_1944 = io_dram_wresp_valid & io_dram_wresp_ready; // @[DRAMArbiter.scala 165:54:@17785.4]
  assign _T_1949 = _T_1947 + 64'h1; // @[DRAMArbiter.scala 121:18:@17788.6]
  assign _T_1950 = _T_1947 + 64'h1; // @[DRAMArbiter.scala 121:18:@17789.6]
  assign _GEN_13 = _T_1944 ? _T_1950 : _T_1947; // @[DRAMArbiter.scala 120:19:@17787.4]
  assign _T_1952 = io_dram_wresp_ready == 1'h0; // @[DRAMArbiter.scala 166:56:@17793.4]
  assign _T_1953 = io_dram_wresp_valid & _T_1952; // @[DRAMArbiter.scala 166:54:@17794.4]
  assign _T_1958 = _T_1956 + 64'h1; // @[DRAMArbiter.scala 121:18:@17797.6]
  assign _T_1959 = _T_1956 + 64'h1; // @[DRAMArbiter.scala 121:18:@17798.6]
  assign _GEN_14 = _T_1953 ? _T_1959 : _T_1956; // @[DRAMArbiter.scala 120:19:@17796.4]
  assign _T_1961 = io_dram_wresp_valid == 1'h0; // @[DRAMArbiter.scala 167:34:@17802.4]
  assign _T_1962 = _T_1961 & io_dram_wresp_ready; // @[DRAMArbiter.scala 167:55:@17803.4]
  assign _T_1967 = _T_1965 + 64'h1; // @[DRAMArbiter.scala 121:18:@17806.6]
  assign _T_1968 = _T_1965 + 64'h1; // @[DRAMArbiter.scala 121:18:@17807.6]
  assign _GEN_15 = _T_1962 ? _T_1968 : _T_1965; // @[DRAMArbiter.scala 120:19:@17805.4]
  assign _T_1969 = io_dram_cmd_valid & io_dram_cmd_ready; // @[DRAMArbiter.scala 174:70:@17811.4]
  assign _GEN_16 = _T_1969 ? io_dram_cmd_bits_addr : _T_1971; // @[DRAMArbiter.scala 128:19:@17813.4]
  assign _GEN_17 = _T_1969 ? io_dram_cmd_bits_size : _T_1974; // @[DRAMArbiter.scala 128:19:@17819.4]
  assign _GEN_18 = _T_1846 ? io_dram_wdata_bits_wdata_0 : _T_1977; // @[DRAMArbiter.scala 128:19:@17825.4]
  assign _GEN_19 = _T_1846 ? io_dram_wdata_bits_wstrb_0 : _T_1980; // @[DRAMArbiter.scala 128:19:@17831.4]
  assign _T_1983 = _T_1849 == 64'h0; // @[DRAMArbiter.scala 178:115:@17836.4]
  assign _T_1984 = _T_1846 & _T_1983; // @[DRAMArbiter.scala 178:102:@17837.4]
  assign _GEN_20 = _T_1984 ? io_dram_wdata_bits_wdata_0 : _T_1986; // @[DRAMArbiter.scala 128:19:@17839.4]
  assign _GEN_21 = _T_1984 ? io_dram_wdata_bits_wstrb_0 : _T_1992; // @[DRAMArbiter.scala 128:19:@17847.4]
  assign _T_1995 = _T_1849 == 64'h1; // @[DRAMArbiter.scala 180:115:@17852.4]
  assign _T_1996 = _T_1846 & _T_1995; // @[DRAMArbiter.scala 180:102:@17853.4]
  assign _GEN_22 = _T_1996 ? io_dram_wdata_bits_wdata_0 : _T_1998; // @[DRAMArbiter.scala 128:19:@17855.4]
  assign _GEN_23 = _T_1996 ? io_dram_wdata_bits_wstrb_0 : _T_2004; // @[DRAMArbiter.scala 128:19:@17863.4]
  assign _T_2005 = io_app_stores_0_cmd_valid & io_app_stores_0_cmd_ready; // @[DRAMArbiter.scala 182:92:@17867.4]
  assign _GEN_24 = _T_2005 ? io_app_stores_0_cmd_bits_addr : _T_2007; // @[DRAMArbiter.scala 128:19:@17869.4]
  assign _GEN_25 = _T_2005 ? io_app_stores_0_cmd_bits_size : _T_2010; // @[DRAMArbiter.scala 128:19:@17875.4]
  assign _GEN_26 = _T_1853 ? io_app_stores_0_data_bits_wdata_0 : _T_2013; // @[DRAMArbiter.scala 128:19:@17881.4]
  assign _GEN_27 = _T_1853 ? io_app_stores_0_data_bits_wstrb : _T_2016; // @[DRAMArbiter.scala 128:19:@17887.4]
  assign _T_2019 = _T_1856 == 64'h0; // @[DRAMArbiter.scala 186:148:@17892.4]
  assign _T_2020 = _T_1853 & _T_2019; // @[DRAMArbiter.scala 186:132:@17893.4]
  assign _GEN_28 = _T_2020 ? io_app_stores_0_data_bits_wdata_0 : _T_2022; // @[DRAMArbiter.scala 128:19:@17895.4]
  assign _GEN_29 = _T_2020 ? io_app_stores_0_data_bits_wstrb : _T_2028; // @[DRAMArbiter.scala 128:19:@17903.4]
  assign _T_2031 = _T_1856 == 64'h1; // @[DRAMArbiter.scala 188:148:@17908.4]
  assign _T_2032 = _T_1853 & _T_2031; // @[DRAMArbiter.scala 188:132:@17909.4]
  assign _GEN_30 = _T_2032 ? io_app_stores_0_data_bits_wdata_0 : _T_2034; // @[DRAMArbiter.scala 128:19:@17911.4]
  assign _GEN_31 = _T_2032 ? io_app_stores_0_data_bits_wstrb : _T_2040; // @[DRAMArbiter.scala 128:19:@17919.4]
  assign _T_2114 = _T_2112 + 64'h1; // @[DRAMArbiter.scala 121:18:@18002.6]
  assign _T_2115 = _T_2112 + 64'h1; // @[DRAMArbiter.scala 121:18:@18003.6]
  assign io_app_loads_0_cmd_ready = StreamControllerLoad_io_load_cmd_ready; // @[DRAMArbiter.scala 61:17:@17091.4]
  assign io_app_loads_0_data_valid = StreamControllerLoad_io_load_data_valid; // @[DRAMArbiter.scala 61:17:@17086.4]
  assign io_app_loads_0_data_bits_rdata_0 = StreamControllerLoad_io_load_data_bits_rdata_0; // @[DRAMArbiter.scala 61:17:@17085.4]
  assign io_app_stores_0_cmd_ready = 1'h0;
  assign io_app_stores_0_data_ready = 1'h0;
  assign io_dram_cmd_valid = io_enable & AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 99:13:@17660.4 DRAMArbiter.scala 100:23:@17663.4]
  assign io_dram_cmd_bits_addr = AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 99:13:@17659.4]
  assign io_dram_cmd_bits_size = AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 99:13:@17658.4]
  assign io_dram_cmd_bits_isWr = 1'h0; // @[DRAMArbiter.scala 99:13:@17656.4]
  assign io_dram_cmd_bits_tag = AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 99:13:@17655.4]
  assign io_dram_wdata_valid = 1'h0; // @[DRAMArbiter.scala 99:13:@17653.4 DRAMArbiter.scala 101:25:@17665.4]
  assign io_dram_wdata_bits_wdata_0 = 32'h0; // @[DRAMArbiter.scala 99:13:@17637.4]
  assign io_dram_wdata_bits_wstrb_0 = 1'h0; // @[DRAMArbiter.scala 99:13:@17573.4]
  assign io_dram_wdata_bits_wlast = AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 99:13:@17572.4]
  assign io_dram_rresp_ready = AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 99:13:@17571.4]
  assign io_dram_wresp_ready = AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 99:13:@17552.4]
  assign io_debugSignals_0 = _T_1835[31:0]; // @[DRAMArbiter.scala 110:39:@17672.4]
  assign io_debugSignals_1 = _T_1849[31:0]; // @[DRAMArbiter.scala 110:39:@17694.4]
  assign io_debugSignals_2 = _T_1863[31:0]; // @[DRAMArbiter.scala 110:39:@17702.4]
  assign io_debugSignals_3 = _T_1873[31:0]; // @[DRAMArbiter.scala 110:39:@17712.4]
  assign io_debugSignals_4 = _T_1881[31:0]; // @[DRAMArbiter.scala 110:39:@17721.4]
  assign io_debugSignals_5 = _T_1889[31:0]; // @[DRAMArbiter.scala 110:39:@17730.4]
  assign io_debugSignals_6 = _T_1897[31:0]; // @[DRAMArbiter.scala 110:39:@17739.4]
  assign io_debugSignals_7 = _T_1904[31:0]; // @[DRAMArbiter.scala 110:39:@17747.4]
  assign io_debugSignals_8 = _T_1913[31:0]; // @[DRAMArbiter.scala 110:39:@17756.4]
  assign io_debugSignals_9 = _T_1922[31:0]; // @[DRAMArbiter.scala 110:39:@17765.4]
  assign io_debugSignals_10 = _T_1940[31:0]; // @[DRAMArbiter.scala 110:39:@17784.4]
  assign io_debugSignals_11 = _T_1947[31:0]; // @[DRAMArbiter.scala 110:39:@17792.4]
  assign io_debugSignals_12 = _T_1956[31:0]; // @[DRAMArbiter.scala 110:39:@17801.4]
  assign io_debugSignals_13 = _T_1965[31:0]; // @[DRAMArbiter.scala 110:39:@17810.4]
  assign io_debugSignals_14 = _T_1971[31:0]; // @[DRAMArbiter.scala 110:39:@17816.4]
  assign io_debugSignals_15 = _T_1974; // @[DRAMArbiter.scala 110:39:@17822.4]
  assign io_debugSignals_16 = _T_1977; // @[DRAMArbiter.scala 110:39:@17828.4]
  assign io_debugSignals_17 = {{31'd0}, _T_1980}; // @[DRAMArbiter.scala 110:39:@17834.4]
  assign io_debugSignals_18 = _T_1986; // @[DRAMArbiter.scala 110:39:@17842.4]
  assign io_debugSignals_19 = {{31'd0}, _T_1992}; // @[DRAMArbiter.scala 110:39:@17850.4]
  assign io_debugSignals_20 = _T_1998; // @[DRAMArbiter.scala 110:39:@17858.4]
  assign io_debugSignals_21 = {{31'd0}, _T_2004}; // @[DRAMArbiter.scala 110:39:@17866.4]
  assign io_debugSignals_22 = _T_2007[31:0]; // @[DRAMArbiter.scala 110:39:@17872.4]
  assign io_debugSignals_23 = _T_2010; // @[DRAMArbiter.scala 110:39:@17878.4]
  assign io_debugSignals_24 = _T_2013; // @[DRAMArbiter.scala 110:39:@17884.4]
  assign io_debugSignals_25 = {{16'd0}, _T_2016}; // @[DRAMArbiter.scala 110:39:@17890.4]
  assign io_debugSignals_26 = _T_2022; // @[DRAMArbiter.scala 110:39:@17898.4]
  assign io_debugSignals_27 = {{16'd0}, _T_2028}; // @[DRAMArbiter.scala 110:39:@17906.4]
  assign io_debugSignals_28 = _T_2034; // @[DRAMArbiter.scala 110:39:@17914.4]
  assign io_debugSignals_29 = {{16'd0}, _T_2040}; // @[DRAMArbiter.scala 110:39:@17922.4]
  assign io_debugSignals_40 = _T_2112[31:0]; // @[DRAMArbiter.scala 110:39:@18006.4]
  assign StreamControllerLoad_clock = clock; // @[:@17083.4]
  assign StreamControllerLoad_reset = reset; // @[:@17084.4]
  assign StreamControllerLoad_io_dram_cmd_ready = StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 87:32:@17207.4]
  assign StreamControllerLoad_io_dram_rresp_valid = StreamArbiter_io_app_0_rresp_valid; // @[DRAMArbiter.scala 87:32:@17116.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_0 = StreamArbiter_io_app_0_rresp_bits_rdata_0; // @[DRAMArbiter.scala 87:32:@17100.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_1 = StreamArbiter_io_app_0_rresp_bits_rdata_1; // @[DRAMArbiter.scala 87:32:@17101.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_2 = StreamArbiter_io_app_0_rresp_bits_rdata_2; // @[DRAMArbiter.scala 87:32:@17102.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_3 = StreamArbiter_io_app_0_rresp_bits_rdata_3; // @[DRAMArbiter.scala 87:32:@17103.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_4 = StreamArbiter_io_app_0_rresp_bits_rdata_4; // @[DRAMArbiter.scala 87:32:@17104.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_5 = StreamArbiter_io_app_0_rresp_bits_rdata_5; // @[DRAMArbiter.scala 87:32:@17105.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_6 = StreamArbiter_io_app_0_rresp_bits_rdata_6; // @[DRAMArbiter.scala 87:32:@17106.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_7 = StreamArbiter_io_app_0_rresp_bits_rdata_7; // @[DRAMArbiter.scala 87:32:@17107.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_8 = StreamArbiter_io_app_0_rresp_bits_rdata_8; // @[DRAMArbiter.scala 87:32:@17108.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_9 = StreamArbiter_io_app_0_rresp_bits_rdata_9; // @[DRAMArbiter.scala 87:32:@17109.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_10 = StreamArbiter_io_app_0_rresp_bits_rdata_10; // @[DRAMArbiter.scala 87:32:@17110.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_11 = StreamArbiter_io_app_0_rresp_bits_rdata_11; // @[DRAMArbiter.scala 87:32:@17111.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_12 = StreamArbiter_io_app_0_rresp_bits_rdata_12; // @[DRAMArbiter.scala 87:32:@17112.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_13 = StreamArbiter_io_app_0_rresp_bits_rdata_13; // @[DRAMArbiter.scala 87:32:@17113.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_14 = StreamArbiter_io_app_0_rresp_bits_rdata_14; // @[DRAMArbiter.scala 87:32:@17114.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_15 = StreamArbiter_io_app_0_rresp_bits_rdata_15; // @[DRAMArbiter.scala 87:32:@17115.4]
  assign StreamControllerLoad_io_load_cmd_valid = io_app_loads_0_cmd_valid; // @[DRAMArbiter.scala 61:17:@17090.4]
  assign StreamControllerLoad_io_load_cmd_bits_addr = io_app_loads_0_cmd_bits_addr; // @[DRAMArbiter.scala 61:17:@17089.4]
  assign StreamControllerLoad_io_load_cmd_bits_size = io_app_loads_0_cmd_bits_size; // @[DRAMArbiter.scala 61:17:@17088.4]
  assign StreamControllerLoad_io_load_data_ready = io_app_loads_0_data_ready; // @[DRAMArbiter.scala 61:17:@17087.4]
  assign StreamArbiter_clock = clock; // @[:@17093.4]
  assign StreamArbiter_reset = reset; // @[:@17094.4]
  assign StreamArbiter_io_app_0_cmd_valid = StreamControllerLoad_io_dram_cmd_valid; // @[DRAMArbiter.scala 87:22:@17318.4]
  assign StreamArbiter_io_app_0_cmd_bits_addr = StreamControllerLoad_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 87:22:@17317.4]
  assign StreamArbiter_io_app_0_cmd_bits_size = StreamControllerLoad_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 87:22:@17316.4]
  assign StreamArbiter_io_app_0_rresp_ready = StreamControllerLoad_io_dram_rresp_ready; // @[DRAMArbiter.scala 87:22:@17229.4]
  assign StreamArbiter_io_dram_cmd_ready = AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 95:20:@17434.4]
  assign StreamArbiter_io_dram_rresp_valid = AXICmdSplit_io_in_rresp_valid; // @[DRAMArbiter.scala 95:20:@17343.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_0 = AXICmdSplit_io_in_rresp_bits_rdata_0; // @[DRAMArbiter.scala 95:20:@17327.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_1 = AXICmdSplit_io_in_rresp_bits_rdata_1; // @[DRAMArbiter.scala 95:20:@17328.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_2 = AXICmdSplit_io_in_rresp_bits_rdata_2; // @[DRAMArbiter.scala 95:20:@17329.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_3 = AXICmdSplit_io_in_rresp_bits_rdata_3; // @[DRAMArbiter.scala 95:20:@17330.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_4 = AXICmdSplit_io_in_rresp_bits_rdata_4; // @[DRAMArbiter.scala 95:20:@17331.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_5 = AXICmdSplit_io_in_rresp_bits_rdata_5; // @[DRAMArbiter.scala 95:20:@17332.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_6 = AXICmdSplit_io_in_rresp_bits_rdata_6; // @[DRAMArbiter.scala 95:20:@17333.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_7 = AXICmdSplit_io_in_rresp_bits_rdata_7; // @[DRAMArbiter.scala 95:20:@17334.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_8 = AXICmdSplit_io_in_rresp_bits_rdata_8; // @[DRAMArbiter.scala 95:20:@17335.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_9 = AXICmdSplit_io_in_rresp_bits_rdata_9; // @[DRAMArbiter.scala 95:20:@17336.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_10 = AXICmdSplit_io_in_rresp_bits_rdata_10; // @[DRAMArbiter.scala 95:20:@17337.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_11 = AXICmdSplit_io_in_rresp_bits_rdata_11; // @[DRAMArbiter.scala 95:20:@17338.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_12 = AXICmdSplit_io_in_rresp_bits_rdata_12; // @[DRAMArbiter.scala 95:20:@17339.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_13 = AXICmdSplit_io_in_rresp_bits_rdata_13; // @[DRAMArbiter.scala 95:20:@17340.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_14 = AXICmdSplit_io_in_rresp_bits_rdata_14; // @[DRAMArbiter.scala 95:20:@17341.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_15 = AXICmdSplit_io_in_rresp_bits_rdata_15; // @[DRAMArbiter.scala 95:20:@17342.4]
  assign StreamArbiter_io_dram_rresp_bits_tag = AXICmdSplit_io_in_rresp_bits_tag; // @[DRAMArbiter.scala 95:20:@17326.4]
  assign AXICmdSplit_clock = clock; // @[:@17321.4]
  assign AXICmdSplit_reset = reset; // @[:@17322.4]
  assign AXICmdSplit_io_in_cmd_valid = StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 95:20:@17433.4]
  assign AXICmdSplit_io_in_cmd_bits_addr = StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 95:20:@17432.4]
  assign AXICmdSplit_io_in_cmd_bits_size = StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 95:20:@17431.4]
  assign AXICmdSplit_io_in_rresp_ready = StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 95:20:@17344.4]
  assign AXICmdSplit_io_out_cmd_ready = AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 98:20:@17549.4]
  assign AXICmdSplit_io_out_rresp_valid = AXICmdIssue_io_in_rresp_valid; // @[DRAMArbiter.scala 98:20:@17458.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_0 = AXICmdIssue_io_in_rresp_bits_rdata_0; // @[DRAMArbiter.scala 98:20:@17442.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_1 = AXICmdIssue_io_in_rresp_bits_rdata_1; // @[DRAMArbiter.scala 98:20:@17443.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_2 = AXICmdIssue_io_in_rresp_bits_rdata_2; // @[DRAMArbiter.scala 98:20:@17444.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_3 = AXICmdIssue_io_in_rresp_bits_rdata_3; // @[DRAMArbiter.scala 98:20:@17445.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_4 = AXICmdIssue_io_in_rresp_bits_rdata_4; // @[DRAMArbiter.scala 98:20:@17446.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_5 = AXICmdIssue_io_in_rresp_bits_rdata_5; // @[DRAMArbiter.scala 98:20:@17447.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_6 = AXICmdIssue_io_in_rresp_bits_rdata_6; // @[DRAMArbiter.scala 98:20:@17448.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_7 = AXICmdIssue_io_in_rresp_bits_rdata_7; // @[DRAMArbiter.scala 98:20:@17449.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_8 = AXICmdIssue_io_in_rresp_bits_rdata_8; // @[DRAMArbiter.scala 98:20:@17450.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_9 = AXICmdIssue_io_in_rresp_bits_rdata_9; // @[DRAMArbiter.scala 98:20:@17451.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_10 = AXICmdIssue_io_in_rresp_bits_rdata_10; // @[DRAMArbiter.scala 98:20:@17452.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_11 = AXICmdIssue_io_in_rresp_bits_rdata_11; // @[DRAMArbiter.scala 98:20:@17453.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_12 = AXICmdIssue_io_in_rresp_bits_rdata_12; // @[DRAMArbiter.scala 98:20:@17454.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_13 = AXICmdIssue_io_in_rresp_bits_rdata_13; // @[DRAMArbiter.scala 98:20:@17455.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_14 = AXICmdIssue_io_in_rresp_bits_rdata_14; // @[DRAMArbiter.scala 98:20:@17456.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_15 = AXICmdIssue_io_in_rresp_bits_rdata_15; // @[DRAMArbiter.scala 98:20:@17457.4]
  assign AXICmdSplit_io_out_rresp_bits_tag = AXICmdIssue_io_in_rresp_bits_tag; // @[DRAMArbiter.scala 98:20:@17441.4]
  assign AXICmdSplit_io_out_wresp_bits_tag = AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 98:20:@17438.4]
  assign AXICmdIssue_clock = clock; // @[:@17436.4]
  assign AXICmdIssue_reset = reset; // @[:@17437.4]
  assign AXICmdIssue_io_in_cmd_valid = AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 98:20:@17548.4]
  assign AXICmdIssue_io_in_cmd_bits_addr = AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 98:20:@17547.4]
  assign AXICmdIssue_io_in_cmd_bits_size = AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 98:20:@17546.4]
  assign AXICmdIssue_io_in_cmd_bits_tag = AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 98:20:@17543.4]
  assign AXICmdIssue_io_in_rresp_ready = AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 98:20:@17459.4]
  assign AXICmdIssue_io_in_wresp_ready = AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 98:20:@17440.4]
  assign AXICmdIssue_io_out_cmd_ready = io_dram_cmd_ready; // @[DRAMArbiter.scala 99:13:@17661.4]
  assign AXICmdIssue_io_out_wdata_ready = io_dram_wdata_ready; // @[DRAMArbiter.scala 99:13:@17654.4]
  assign AXICmdIssue_io_out_rresp_valid = io_dram_rresp_valid; // @[DRAMArbiter.scala 99:13:@17570.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_0 = io_dram_rresp_bits_rdata_0; // @[DRAMArbiter.scala 99:13:@17554.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_1 = io_dram_rresp_bits_rdata_1; // @[DRAMArbiter.scala 99:13:@17555.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_2 = io_dram_rresp_bits_rdata_2; // @[DRAMArbiter.scala 99:13:@17556.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_3 = io_dram_rresp_bits_rdata_3; // @[DRAMArbiter.scala 99:13:@17557.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_4 = io_dram_rresp_bits_rdata_4; // @[DRAMArbiter.scala 99:13:@17558.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_5 = io_dram_rresp_bits_rdata_5; // @[DRAMArbiter.scala 99:13:@17559.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_6 = io_dram_rresp_bits_rdata_6; // @[DRAMArbiter.scala 99:13:@17560.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_7 = io_dram_rresp_bits_rdata_7; // @[DRAMArbiter.scala 99:13:@17561.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_8 = io_dram_rresp_bits_rdata_8; // @[DRAMArbiter.scala 99:13:@17562.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_9 = io_dram_rresp_bits_rdata_9; // @[DRAMArbiter.scala 99:13:@17563.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_10 = io_dram_rresp_bits_rdata_10; // @[DRAMArbiter.scala 99:13:@17564.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_11 = io_dram_rresp_bits_rdata_11; // @[DRAMArbiter.scala 99:13:@17565.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_12 = io_dram_rresp_bits_rdata_12; // @[DRAMArbiter.scala 99:13:@17566.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_13 = io_dram_rresp_bits_rdata_13; // @[DRAMArbiter.scala 99:13:@17567.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_14 = io_dram_rresp_bits_rdata_14; // @[DRAMArbiter.scala 99:13:@17568.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_15 = io_dram_rresp_bits_rdata_15; // @[DRAMArbiter.scala 99:13:@17569.4]
  assign AXICmdIssue_io_out_rresp_bits_tag = io_dram_rresp_bits_tag; // @[DRAMArbiter.scala 99:13:@17553.4]
  assign AXICmdIssue_io_out_wresp_bits_tag = io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 99:13:@17550.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  _T_1835 = _RAND_0[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {2{`RANDOM}};
  _T_1849 = _RAND_1[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {2{`RANDOM}};
  _T_1856 = _RAND_2[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {2{`RANDOM}};
  _T_1863 = _RAND_3[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {2{`RANDOM}};
  _T_1873 = _RAND_4[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {2{`RANDOM}};
  _T_1881 = _RAND_5[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {2{`RANDOM}};
  _T_1889 = _RAND_6[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {2{`RANDOM}};
  _T_1897 = _RAND_7[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {2{`RANDOM}};
  _T_1904 = _RAND_8[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {2{`RANDOM}};
  _T_1913 = _RAND_9[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {2{`RANDOM}};
  _T_1922 = _RAND_10[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {2{`RANDOM}};
  _T_1940 = _RAND_11[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {2{`RANDOM}};
  _T_1947 = _RAND_12[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {2{`RANDOM}};
  _T_1956 = _RAND_13[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {2{`RANDOM}};
  _T_1965 = _RAND_14[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {2{`RANDOM}};
  _T_1971 = _RAND_15[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_1974 = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_1977 = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_1980 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_1986 = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_1992 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_1998 = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_2004 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {2{`RANDOM}};
  _T_2007 = _RAND_23[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_2010 = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_2013 = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_2016 = _RAND_26[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_2022 = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_2028 = _RAND_28[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_2034 = _RAND_29[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_2040 = _RAND_30[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {2{`RANDOM}};
  _T_2112 = _RAND_31[63:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_1835 <= 64'h0;
    end else begin
      if (io_enable) begin
        _T_1835 <= _T_1838;
      end
    end
    if (reset) begin
      _T_1849 <= 64'h0;
    end else begin
      if (_T_1846) begin
        _T_1849 <= _T_1852;
      end
    end
    if (reset) begin
      _T_1856 <= 64'h0;
    end else begin
      if (_T_1853) begin
        _T_1856 <= _T_1859;
      end
    end
    if (reset) begin
      _T_1863 <= 64'h0;
    end else begin
      if (_T_1860) begin
        _T_1863 <= _T_1866;
      end
    end
    if (reset) begin
      _T_1873 <= 64'h0;
    end else begin
      if (_T_1870) begin
        _T_1873 <= _T_1876;
      end
    end
    if (reset) begin
      _T_1881 <= 64'h0;
    end else begin
      if (_T_1878) begin
        _T_1881 <= _T_1884;
      end
    end
    if (reset) begin
      _T_1889 <= 64'h0;
    end else begin
      if (_T_1886) begin
        _T_1889 <= _T_1892;
      end
    end
    if (reset) begin
      _T_1897 <= 64'h0;
    end else begin
      if (_T_1894) begin
        _T_1897 <= _T_1900;
      end
    end
    if (reset) begin
      _T_1904 <= 64'h0;
    end else begin
      if (_T_1839) begin
        _T_1904 <= _T_1907;
      end
    end
    if (reset) begin
      _T_1913 <= 64'h0;
    end else begin
      if (_T_1910) begin
        _T_1913 <= _T_1916;
      end
    end
    if (reset) begin
      _T_1922 <= 64'h0;
    end else begin
      if (_T_1919) begin
        _T_1922 <= _T_1925;
      end
    end
    if (reset) begin
      _T_1940 <= 64'h0;
    end else begin
      if (_T_1937) begin
        _T_1940 <= _T_1943;
      end
    end
    if (reset) begin
      _T_1947 <= 64'h0;
    end else begin
      if (_T_1944) begin
        _T_1947 <= _T_1950;
      end
    end
    if (reset) begin
      _T_1956 <= 64'h0;
    end else begin
      if (_T_1953) begin
        _T_1956 <= _T_1959;
      end
    end
    if (reset) begin
      _T_1965 <= 64'h0;
    end else begin
      if (_T_1962) begin
        _T_1965 <= _T_1968;
      end
    end
    if (reset) begin
      _T_1971 <= io_dram_cmd_bits_addr;
    end else begin
      if (_T_1969) begin
        _T_1971 <= io_dram_cmd_bits_addr;
      end
    end
    if (reset) begin
      _T_1974 <= io_dram_cmd_bits_size;
    end else begin
      if (_T_1969) begin
        _T_1974 <= io_dram_cmd_bits_size;
      end
    end
    if (reset) begin
      _T_1977 <= io_dram_wdata_bits_wdata_0;
    end else begin
      if (_T_1846) begin
        _T_1977 <= io_dram_wdata_bits_wdata_0;
      end
    end
    if (reset) begin
      _T_1980 <= io_dram_wdata_bits_wstrb_0;
    end else begin
      if (_T_1846) begin
        _T_1980 <= io_dram_wdata_bits_wstrb_0;
      end
    end
    if (reset) begin
      _T_1986 <= io_dram_wdata_bits_wdata_0;
    end else begin
      if (_T_1984) begin
        _T_1986 <= io_dram_wdata_bits_wdata_0;
      end
    end
    if (reset) begin
      _T_1992 <= io_dram_wdata_bits_wstrb_0;
    end else begin
      if (_T_1984) begin
        _T_1992 <= io_dram_wdata_bits_wstrb_0;
      end
    end
    if (reset) begin
      _T_1998 <= io_dram_wdata_bits_wdata_0;
    end else begin
      if (_T_1996) begin
        _T_1998 <= io_dram_wdata_bits_wdata_0;
      end
    end
    if (reset) begin
      _T_2004 <= io_dram_wdata_bits_wstrb_0;
    end else begin
      if (_T_1996) begin
        _T_2004 <= io_dram_wdata_bits_wstrb_0;
      end
    end
    if (reset) begin
      _T_2007 <= io_app_stores_0_cmd_bits_addr;
    end else begin
      if (_T_2005) begin
        _T_2007 <= io_app_stores_0_cmd_bits_addr;
      end
    end
    if (reset) begin
      _T_2010 <= io_app_stores_0_cmd_bits_size;
    end else begin
      if (_T_2005) begin
        _T_2010 <= io_app_stores_0_cmd_bits_size;
      end
    end
    if (reset) begin
      _T_2013 <= io_app_stores_0_data_bits_wdata_0;
    end else begin
      if (_T_1853) begin
        _T_2013 <= io_app_stores_0_data_bits_wdata_0;
      end
    end
    if (reset) begin
      _T_2016 <= io_app_stores_0_data_bits_wstrb;
    end else begin
      if (_T_1853) begin
        _T_2016 <= io_app_stores_0_data_bits_wstrb;
      end
    end
    if (reset) begin
      _T_2022 <= io_app_stores_0_data_bits_wdata_0;
    end else begin
      if (_T_2020) begin
        _T_2022 <= io_app_stores_0_data_bits_wdata_0;
      end
    end
    if (reset) begin
      _T_2028 <= io_app_stores_0_data_bits_wstrb;
    end else begin
      if (_T_2020) begin
        _T_2028 <= io_app_stores_0_data_bits_wstrb;
      end
    end
    if (reset) begin
      _T_2034 <= io_app_stores_0_data_bits_wdata_0;
    end else begin
      if (_T_2032) begin
        _T_2034 <= io_app_stores_0_data_bits_wdata_0;
      end
    end
    if (reset) begin
      _T_2040 <= io_app_stores_0_data_bits_wstrb;
    end else begin
      if (_T_2032) begin
        _T_2040 <= io_app_stores_0_data_bits_wstrb;
      end
    end
    if (reset) begin
      _T_2112 <= 64'h0;
    end else begin
      _T_2112 <= _T_2115;
    end
  end
endmodule
module DRAMHeap( // @[:@18109.2]
  input         io_accel_0_req_valid, // @[:@18112.4]
  input         io_accel_0_req_bits_allocDealloc, // @[:@18112.4]
  input  [63:0] io_accel_0_req_bits_sizeAddr, // @[:@18112.4]
  output        io_accel_0_resp_valid, // @[:@18112.4]
  output        io_accel_0_resp_bits_allocDealloc, // @[:@18112.4]
  output [63:0] io_accel_0_resp_bits_sizeAddr, // @[:@18112.4]
  output        io_host_0_req_valid, // @[:@18112.4]
  output        io_host_0_req_bits_allocDealloc, // @[:@18112.4]
  output [63:0] io_host_0_req_bits_sizeAddr, // @[:@18112.4]
  input         io_host_0_resp_valid, // @[:@18112.4]
  input         io_host_0_resp_bits_allocDealloc, // @[:@18112.4]
  input  [63:0] io_host_0_resp_bits_sizeAddr // @[:@18112.4]
);
  assign io_accel_0_resp_valid = io_host_0_resp_valid; // @[DRAMHeap.scala 24:18:@18119.4]
  assign io_accel_0_resp_bits_allocDealloc = io_host_0_resp_bits_allocDealloc; // @[DRAMHeap.scala 25:17:@18121.4]
  assign io_accel_0_resp_bits_sizeAddr = io_host_0_resp_bits_sizeAddr; // @[DRAMHeap.scala 25:17:@18120.4]
  assign io_host_0_req_valid = io_accel_0_req_valid; // @[DRAMHeap.scala 21:18:@18116.4]
  assign io_host_0_req_bits_allocDealloc = io_accel_0_req_bits_allocDealloc; // @[DRAMHeap.scala 21:18:@18115.4]
  assign io_host_0_req_bits_sizeAddr = io_accel_0_req_bits_sizeAddr; // @[DRAMHeap.scala 21:18:@18114.4]
endmodule
module RetimeWrapper_105( // @[:@18135.2]
  input         clock, // @[:@18136.4]
  input         reset, // @[:@18137.4]
  input         io_flow, // @[:@18138.4]
  input  [63:0] io_in, // @[:@18138.4]
  output [63:0] io_out // @[:@18138.4]
);
  wire [63:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@18140.4]
  wire [63:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@18140.4]
  wire [63:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@18140.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@18140.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@18140.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@18140.4]
  RetimeShiftRegister #(.WIDTH(64), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@18140.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@18153.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@18152.4]
  assign sr_init = 64'h0; // @[RetimeShiftRegister.scala 19:16:@18151.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@18150.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@18149.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@18147.4]
endmodule
module FringeFF( // @[:@18155.2]
  input         clock, // @[:@18156.4]
  input         reset, // @[:@18157.4]
  input  [63:0] io_in, // @[:@18158.4]
  input         io_reset, // @[:@18158.4]
  output [63:0] io_out, // @[:@18158.4]
  input         io_enable // @[:@18158.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@18161.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@18161.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@18161.4]
  wire [63:0] RetimeWrapper_io_in; // @[package.scala 93:22:@18161.4]
  wire [63:0] RetimeWrapper_io_out; // @[package.scala 93:22:@18161.4]
  wire [63:0] _T_18; // @[package.scala 96:25:@18166.4 package.scala 96:25:@18167.4]
  wire [63:0] _GEN_0; // @[FringeFF.scala 21:27:@18172.6]
  RetimeWrapper_105 RetimeWrapper ( // @[package.scala 93:22:@18161.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@18166.4 package.scala 96:25:@18167.4]
  assign _GEN_0 = io_reset ? 64'h0 : _T_18; // @[FringeFF.scala 21:27:@18172.6]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@18178.4]
  assign RetimeWrapper_clock = clock; // @[:@18162.4]
  assign RetimeWrapper_reset = reset; // @[:@18163.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@18165.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _GEN_0; // @[package.scala 94:16:@18164.4]
endmodule
module MuxN( // @[:@47649.2]
  input  [63:0] io_ins_0, // @[:@47652.4]
  input  [63:0] io_ins_1, // @[:@47652.4]
  input  [63:0] io_ins_2, // @[:@47652.4]
  input  [63:0] io_ins_3, // @[:@47652.4]
  input  [63:0] io_ins_4, // @[:@47652.4]
  input  [63:0] io_ins_5, // @[:@47652.4]
  input  [63:0] io_ins_6, // @[:@47652.4]
  input  [63:0] io_ins_7, // @[:@47652.4]
  input  [63:0] io_ins_8, // @[:@47652.4]
  input  [63:0] io_ins_9, // @[:@47652.4]
  input  [63:0] io_ins_10, // @[:@47652.4]
  input  [63:0] io_ins_11, // @[:@47652.4]
  input  [63:0] io_ins_12, // @[:@47652.4]
  input  [63:0] io_ins_13, // @[:@47652.4]
  input  [63:0] io_ins_14, // @[:@47652.4]
  input  [63:0] io_ins_15, // @[:@47652.4]
  input  [63:0] io_ins_16, // @[:@47652.4]
  input  [63:0] io_ins_17, // @[:@47652.4]
  input  [63:0] io_ins_18, // @[:@47652.4]
  input  [63:0] io_ins_19, // @[:@47652.4]
  input  [63:0] io_ins_20, // @[:@47652.4]
  input  [63:0] io_ins_21, // @[:@47652.4]
  input  [63:0] io_ins_22, // @[:@47652.4]
  input  [63:0] io_ins_23, // @[:@47652.4]
  input  [63:0] io_ins_24, // @[:@47652.4]
  input  [63:0] io_ins_25, // @[:@47652.4]
  input  [63:0] io_ins_26, // @[:@47652.4]
  input  [63:0] io_ins_27, // @[:@47652.4]
  input  [63:0] io_ins_28, // @[:@47652.4]
  input  [63:0] io_ins_29, // @[:@47652.4]
  input  [63:0] io_ins_30, // @[:@47652.4]
  input  [63:0] io_ins_31, // @[:@47652.4]
  input  [63:0] io_ins_32, // @[:@47652.4]
  input  [63:0] io_ins_33, // @[:@47652.4]
  input  [63:0] io_ins_34, // @[:@47652.4]
  input  [63:0] io_ins_35, // @[:@47652.4]
  input  [63:0] io_ins_36, // @[:@47652.4]
  input  [63:0] io_ins_37, // @[:@47652.4]
  input  [63:0] io_ins_38, // @[:@47652.4]
  input  [63:0] io_ins_39, // @[:@47652.4]
  input  [63:0] io_ins_40, // @[:@47652.4]
  input  [63:0] io_ins_41, // @[:@47652.4]
  input  [63:0] io_ins_42, // @[:@47652.4]
  input  [63:0] io_ins_43, // @[:@47652.4]
  input  [63:0] io_ins_44, // @[:@47652.4]
  input  [63:0] io_ins_45, // @[:@47652.4]
  input  [63:0] io_ins_46, // @[:@47652.4]
  input  [63:0] io_ins_47, // @[:@47652.4]
  input  [63:0] io_ins_48, // @[:@47652.4]
  input  [63:0] io_ins_49, // @[:@47652.4]
  input  [63:0] io_ins_50, // @[:@47652.4]
  input  [63:0] io_ins_51, // @[:@47652.4]
  input  [63:0] io_ins_52, // @[:@47652.4]
  input  [63:0] io_ins_53, // @[:@47652.4]
  input  [63:0] io_ins_54, // @[:@47652.4]
  input  [63:0] io_ins_55, // @[:@47652.4]
  input  [63:0] io_ins_56, // @[:@47652.4]
  input  [63:0] io_ins_57, // @[:@47652.4]
  input  [63:0] io_ins_58, // @[:@47652.4]
  input  [63:0] io_ins_59, // @[:@47652.4]
  input  [63:0] io_ins_60, // @[:@47652.4]
  input  [63:0] io_ins_61, // @[:@47652.4]
  input  [63:0] io_ins_62, // @[:@47652.4]
  input  [63:0] io_ins_63, // @[:@47652.4]
  input  [63:0] io_ins_64, // @[:@47652.4]
  input  [63:0] io_ins_65, // @[:@47652.4]
  input  [63:0] io_ins_66, // @[:@47652.4]
  input  [63:0] io_ins_67, // @[:@47652.4]
  input  [63:0] io_ins_68, // @[:@47652.4]
  input  [63:0] io_ins_69, // @[:@47652.4]
  input  [63:0] io_ins_70, // @[:@47652.4]
  input  [63:0] io_ins_71, // @[:@47652.4]
  input  [63:0] io_ins_72, // @[:@47652.4]
  input  [63:0] io_ins_73, // @[:@47652.4]
  input  [63:0] io_ins_74, // @[:@47652.4]
  input  [63:0] io_ins_75, // @[:@47652.4]
  input  [63:0] io_ins_76, // @[:@47652.4]
  input  [63:0] io_ins_77, // @[:@47652.4]
  input  [63:0] io_ins_78, // @[:@47652.4]
  input  [63:0] io_ins_79, // @[:@47652.4]
  input  [63:0] io_ins_80, // @[:@47652.4]
  input  [63:0] io_ins_81, // @[:@47652.4]
  input  [63:0] io_ins_82, // @[:@47652.4]
  input  [63:0] io_ins_83, // @[:@47652.4]
  input  [63:0] io_ins_84, // @[:@47652.4]
  input  [63:0] io_ins_85, // @[:@47652.4]
  input  [63:0] io_ins_86, // @[:@47652.4]
  input  [63:0] io_ins_87, // @[:@47652.4]
  input  [63:0] io_ins_88, // @[:@47652.4]
  input  [63:0] io_ins_89, // @[:@47652.4]
  input  [63:0] io_ins_90, // @[:@47652.4]
  input  [63:0] io_ins_91, // @[:@47652.4]
  input  [63:0] io_ins_92, // @[:@47652.4]
  input  [63:0] io_ins_93, // @[:@47652.4]
  input  [63:0] io_ins_94, // @[:@47652.4]
  input  [63:0] io_ins_95, // @[:@47652.4]
  input  [63:0] io_ins_96, // @[:@47652.4]
  input  [63:0] io_ins_97, // @[:@47652.4]
  input  [63:0] io_ins_98, // @[:@47652.4]
  input  [63:0] io_ins_99, // @[:@47652.4]
  input  [63:0] io_ins_100, // @[:@47652.4]
  input  [63:0] io_ins_101, // @[:@47652.4]
  input  [63:0] io_ins_102, // @[:@47652.4]
  input  [63:0] io_ins_103, // @[:@47652.4]
  input  [63:0] io_ins_104, // @[:@47652.4]
  input  [63:0] io_ins_105, // @[:@47652.4]
  input  [63:0] io_ins_106, // @[:@47652.4]
  input  [63:0] io_ins_107, // @[:@47652.4]
  input  [63:0] io_ins_108, // @[:@47652.4]
  input  [63:0] io_ins_109, // @[:@47652.4]
  input  [63:0] io_ins_110, // @[:@47652.4]
  input  [63:0] io_ins_111, // @[:@47652.4]
  input  [63:0] io_ins_112, // @[:@47652.4]
  input  [63:0] io_ins_113, // @[:@47652.4]
  input  [63:0] io_ins_114, // @[:@47652.4]
  input  [63:0] io_ins_115, // @[:@47652.4]
  input  [63:0] io_ins_116, // @[:@47652.4]
  input  [63:0] io_ins_117, // @[:@47652.4]
  input  [63:0] io_ins_118, // @[:@47652.4]
  input  [63:0] io_ins_119, // @[:@47652.4]
  input  [63:0] io_ins_120, // @[:@47652.4]
  input  [63:0] io_ins_121, // @[:@47652.4]
  input  [63:0] io_ins_122, // @[:@47652.4]
  input  [63:0] io_ins_123, // @[:@47652.4]
  input  [63:0] io_ins_124, // @[:@47652.4]
  input  [63:0] io_ins_125, // @[:@47652.4]
  input  [63:0] io_ins_126, // @[:@47652.4]
  input  [63:0] io_ins_127, // @[:@47652.4]
  input  [63:0] io_ins_128, // @[:@47652.4]
  input  [63:0] io_ins_129, // @[:@47652.4]
  input  [63:0] io_ins_130, // @[:@47652.4]
  input  [63:0] io_ins_131, // @[:@47652.4]
  input  [63:0] io_ins_132, // @[:@47652.4]
  input  [63:0] io_ins_133, // @[:@47652.4]
  input  [63:0] io_ins_134, // @[:@47652.4]
  input  [63:0] io_ins_135, // @[:@47652.4]
  input  [63:0] io_ins_136, // @[:@47652.4]
  input  [63:0] io_ins_137, // @[:@47652.4]
  input  [63:0] io_ins_138, // @[:@47652.4]
  input  [63:0] io_ins_139, // @[:@47652.4]
  input  [63:0] io_ins_140, // @[:@47652.4]
  input  [63:0] io_ins_141, // @[:@47652.4]
  input  [63:0] io_ins_142, // @[:@47652.4]
  input  [63:0] io_ins_143, // @[:@47652.4]
  input  [63:0] io_ins_144, // @[:@47652.4]
  input  [63:0] io_ins_145, // @[:@47652.4]
  input  [63:0] io_ins_146, // @[:@47652.4]
  input  [63:0] io_ins_147, // @[:@47652.4]
  input  [63:0] io_ins_148, // @[:@47652.4]
  input  [63:0] io_ins_149, // @[:@47652.4]
  input  [63:0] io_ins_150, // @[:@47652.4]
  input  [63:0] io_ins_151, // @[:@47652.4]
  input  [63:0] io_ins_152, // @[:@47652.4]
  input  [63:0] io_ins_153, // @[:@47652.4]
  input  [63:0] io_ins_154, // @[:@47652.4]
  input  [63:0] io_ins_155, // @[:@47652.4]
  input  [63:0] io_ins_156, // @[:@47652.4]
  input  [63:0] io_ins_157, // @[:@47652.4]
  input  [63:0] io_ins_158, // @[:@47652.4]
  input  [63:0] io_ins_159, // @[:@47652.4]
  input  [63:0] io_ins_160, // @[:@47652.4]
  input  [63:0] io_ins_161, // @[:@47652.4]
  input  [63:0] io_ins_162, // @[:@47652.4]
  input  [63:0] io_ins_163, // @[:@47652.4]
  input  [63:0] io_ins_164, // @[:@47652.4]
  input  [63:0] io_ins_165, // @[:@47652.4]
  input  [63:0] io_ins_166, // @[:@47652.4]
  input  [63:0] io_ins_167, // @[:@47652.4]
  input  [63:0] io_ins_168, // @[:@47652.4]
  input  [63:0] io_ins_169, // @[:@47652.4]
  input  [63:0] io_ins_170, // @[:@47652.4]
  input  [63:0] io_ins_171, // @[:@47652.4]
  input  [63:0] io_ins_172, // @[:@47652.4]
  input  [63:0] io_ins_173, // @[:@47652.4]
  input  [63:0] io_ins_174, // @[:@47652.4]
  input  [63:0] io_ins_175, // @[:@47652.4]
  input  [63:0] io_ins_176, // @[:@47652.4]
  input  [63:0] io_ins_177, // @[:@47652.4]
  input  [63:0] io_ins_178, // @[:@47652.4]
  input  [63:0] io_ins_179, // @[:@47652.4]
  input  [63:0] io_ins_180, // @[:@47652.4]
  input  [63:0] io_ins_181, // @[:@47652.4]
  input  [63:0] io_ins_182, // @[:@47652.4]
  input  [63:0] io_ins_183, // @[:@47652.4]
  input  [63:0] io_ins_184, // @[:@47652.4]
  input  [63:0] io_ins_185, // @[:@47652.4]
  input  [63:0] io_ins_186, // @[:@47652.4]
  input  [63:0] io_ins_187, // @[:@47652.4]
  input  [63:0] io_ins_188, // @[:@47652.4]
  input  [63:0] io_ins_189, // @[:@47652.4]
  input  [63:0] io_ins_190, // @[:@47652.4]
  input  [63:0] io_ins_191, // @[:@47652.4]
  input  [63:0] io_ins_192, // @[:@47652.4]
  input  [63:0] io_ins_193, // @[:@47652.4]
  input  [63:0] io_ins_194, // @[:@47652.4]
  input  [63:0] io_ins_195, // @[:@47652.4]
  input  [63:0] io_ins_196, // @[:@47652.4]
  input  [63:0] io_ins_197, // @[:@47652.4]
  input  [63:0] io_ins_198, // @[:@47652.4]
  input  [63:0] io_ins_199, // @[:@47652.4]
  input  [63:0] io_ins_200, // @[:@47652.4]
  input  [63:0] io_ins_201, // @[:@47652.4]
  input  [63:0] io_ins_202, // @[:@47652.4]
  input  [63:0] io_ins_203, // @[:@47652.4]
  input  [63:0] io_ins_204, // @[:@47652.4]
  input  [63:0] io_ins_205, // @[:@47652.4]
  input  [63:0] io_ins_206, // @[:@47652.4]
  input  [63:0] io_ins_207, // @[:@47652.4]
  input  [63:0] io_ins_208, // @[:@47652.4]
  input  [63:0] io_ins_209, // @[:@47652.4]
  input  [63:0] io_ins_210, // @[:@47652.4]
  input  [63:0] io_ins_211, // @[:@47652.4]
  input  [63:0] io_ins_212, // @[:@47652.4]
  input  [63:0] io_ins_213, // @[:@47652.4]
  input  [63:0] io_ins_214, // @[:@47652.4]
  input  [63:0] io_ins_215, // @[:@47652.4]
  input  [63:0] io_ins_216, // @[:@47652.4]
  input  [63:0] io_ins_217, // @[:@47652.4]
  input  [63:0] io_ins_218, // @[:@47652.4]
  input  [63:0] io_ins_219, // @[:@47652.4]
  input  [63:0] io_ins_220, // @[:@47652.4]
  input  [63:0] io_ins_221, // @[:@47652.4]
  input  [63:0] io_ins_222, // @[:@47652.4]
  input  [63:0] io_ins_223, // @[:@47652.4]
  input  [63:0] io_ins_224, // @[:@47652.4]
  input  [63:0] io_ins_225, // @[:@47652.4]
  input  [63:0] io_ins_226, // @[:@47652.4]
  input  [63:0] io_ins_227, // @[:@47652.4]
  input  [63:0] io_ins_228, // @[:@47652.4]
  input  [63:0] io_ins_229, // @[:@47652.4]
  input  [63:0] io_ins_230, // @[:@47652.4]
  input  [63:0] io_ins_231, // @[:@47652.4]
  input  [63:0] io_ins_232, // @[:@47652.4]
  input  [63:0] io_ins_233, // @[:@47652.4]
  input  [63:0] io_ins_234, // @[:@47652.4]
  input  [63:0] io_ins_235, // @[:@47652.4]
  input  [63:0] io_ins_236, // @[:@47652.4]
  input  [63:0] io_ins_237, // @[:@47652.4]
  input  [63:0] io_ins_238, // @[:@47652.4]
  input  [63:0] io_ins_239, // @[:@47652.4]
  input  [63:0] io_ins_240, // @[:@47652.4]
  input  [63:0] io_ins_241, // @[:@47652.4]
  input  [63:0] io_ins_242, // @[:@47652.4]
  input  [63:0] io_ins_243, // @[:@47652.4]
  input  [63:0] io_ins_244, // @[:@47652.4]
  input  [63:0] io_ins_245, // @[:@47652.4]
  input  [63:0] io_ins_246, // @[:@47652.4]
  input  [63:0] io_ins_247, // @[:@47652.4]
  input  [63:0] io_ins_248, // @[:@47652.4]
  input  [63:0] io_ins_249, // @[:@47652.4]
  input  [63:0] io_ins_250, // @[:@47652.4]
  input  [63:0] io_ins_251, // @[:@47652.4]
  input  [63:0] io_ins_252, // @[:@47652.4]
  input  [63:0] io_ins_253, // @[:@47652.4]
  input  [63:0] io_ins_254, // @[:@47652.4]
  input  [63:0] io_ins_255, // @[:@47652.4]
  input  [63:0] io_ins_256, // @[:@47652.4]
  input  [63:0] io_ins_257, // @[:@47652.4]
  input  [63:0] io_ins_258, // @[:@47652.4]
  input  [63:0] io_ins_259, // @[:@47652.4]
  input  [63:0] io_ins_260, // @[:@47652.4]
  input  [63:0] io_ins_261, // @[:@47652.4]
  input  [63:0] io_ins_262, // @[:@47652.4]
  input  [63:0] io_ins_263, // @[:@47652.4]
  input  [63:0] io_ins_264, // @[:@47652.4]
  input  [63:0] io_ins_265, // @[:@47652.4]
  input  [63:0] io_ins_266, // @[:@47652.4]
  input  [63:0] io_ins_267, // @[:@47652.4]
  input  [63:0] io_ins_268, // @[:@47652.4]
  input  [63:0] io_ins_269, // @[:@47652.4]
  input  [63:0] io_ins_270, // @[:@47652.4]
  input  [63:0] io_ins_271, // @[:@47652.4]
  input  [63:0] io_ins_272, // @[:@47652.4]
  input  [63:0] io_ins_273, // @[:@47652.4]
  input  [63:0] io_ins_274, // @[:@47652.4]
  input  [63:0] io_ins_275, // @[:@47652.4]
  input  [63:0] io_ins_276, // @[:@47652.4]
  input  [63:0] io_ins_277, // @[:@47652.4]
  input  [63:0] io_ins_278, // @[:@47652.4]
  input  [63:0] io_ins_279, // @[:@47652.4]
  input  [63:0] io_ins_280, // @[:@47652.4]
  input  [63:0] io_ins_281, // @[:@47652.4]
  input  [63:0] io_ins_282, // @[:@47652.4]
  input  [63:0] io_ins_283, // @[:@47652.4]
  input  [63:0] io_ins_284, // @[:@47652.4]
  input  [63:0] io_ins_285, // @[:@47652.4]
  input  [63:0] io_ins_286, // @[:@47652.4]
  input  [63:0] io_ins_287, // @[:@47652.4]
  input  [63:0] io_ins_288, // @[:@47652.4]
  input  [63:0] io_ins_289, // @[:@47652.4]
  input  [63:0] io_ins_290, // @[:@47652.4]
  input  [63:0] io_ins_291, // @[:@47652.4]
  input  [63:0] io_ins_292, // @[:@47652.4]
  input  [63:0] io_ins_293, // @[:@47652.4]
  input  [63:0] io_ins_294, // @[:@47652.4]
  input  [63:0] io_ins_295, // @[:@47652.4]
  input  [63:0] io_ins_296, // @[:@47652.4]
  input  [63:0] io_ins_297, // @[:@47652.4]
  input  [63:0] io_ins_298, // @[:@47652.4]
  input  [63:0] io_ins_299, // @[:@47652.4]
  input  [63:0] io_ins_300, // @[:@47652.4]
  input  [63:0] io_ins_301, // @[:@47652.4]
  input  [63:0] io_ins_302, // @[:@47652.4]
  input  [63:0] io_ins_303, // @[:@47652.4]
  input  [63:0] io_ins_304, // @[:@47652.4]
  input  [63:0] io_ins_305, // @[:@47652.4]
  input  [63:0] io_ins_306, // @[:@47652.4]
  input  [63:0] io_ins_307, // @[:@47652.4]
  input  [63:0] io_ins_308, // @[:@47652.4]
  input  [63:0] io_ins_309, // @[:@47652.4]
  input  [63:0] io_ins_310, // @[:@47652.4]
  input  [63:0] io_ins_311, // @[:@47652.4]
  input  [63:0] io_ins_312, // @[:@47652.4]
  input  [63:0] io_ins_313, // @[:@47652.4]
  input  [63:0] io_ins_314, // @[:@47652.4]
  input  [63:0] io_ins_315, // @[:@47652.4]
  input  [63:0] io_ins_316, // @[:@47652.4]
  input  [63:0] io_ins_317, // @[:@47652.4]
  input  [63:0] io_ins_318, // @[:@47652.4]
  input  [63:0] io_ins_319, // @[:@47652.4]
  input  [63:0] io_ins_320, // @[:@47652.4]
  input  [63:0] io_ins_321, // @[:@47652.4]
  input  [63:0] io_ins_322, // @[:@47652.4]
  input  [63:0] io_ins_323, // @[:@47652.4]
  input  [63:0] io_ins_324, // @[:@47652.4]
  input  [63:0] io_ins_325, // @[:@47652.4]
  input  [63:0] io_ins_326, // @[:@47652.4]
  input  [63:0] io_ins_327, // @[:@47652.4]
  input  [63:0] io_ins_328, // @[:@47652.4]
  input  [63:0] io_ins_329, // @[:@47652.4]
  input  [63:0] io_ins_330, // @[:@47652.4]
  input  [63:0] io_ins_331, // @[:@47652.4]
  input  [63:0] io_ins_332, // @[:@47652.4]
  input  [63:0] io_ins_333, // @[:@47652.4]
  input  [63:0] io_ins_334, // @[:@47652.4]
  input  [63:0] io_ins_335, // @[:@47652.4]
  input  [63:0] io_ins_336, // @[:@47652.4]
  input  [63:0] io_ins_337, // @[:@47652.4]
  input  [63:0] io_ins_338, // @[:@47652.4]
  input  [63:0] io_ins_339, // @[:@47652.4]
  input  [63:0] io_ins_340, // @[:@47652.4]
  input  [63:0] io_ins_341, // @[:@47652.4]
  input  [63:0] io_ins_342, // @[:@47652.4]
  input  [63:0] io_ins_343, // @[:@47652.4]
  input  [63:0] io_ins_344, // @[:@47652.4]
  input  [63:0] io_ins_345, // @[:@47652.4]
  input  [63:0] io_ins_346, // @[:@47652.4]
  input  [63:0] io_ins_347, // @[:@47652.4]
  input  [63:0] io_ins_348, // @[:@47652.4]
  input  [63:0] io_ins_349, // @[:@47652.4]
  input  [63:0] io_ins_350, // @[:@47652.4]
  input  [63:0] io_ins_351, // @[:@47652.4]
  input  [63:0] io_ins_352, // @[:@47652.4]
  input  [63:0] io_ins_353, // @[:@47652.4]
  input  [63:0] io_ins_354, // @[:@47652.4]
  input  [63:0] io_ins_355, // @[:@47652.4]
  input  [63:0] io_ins_356, // @[:@47652.4]
  input  [63:0] io_ins_357, // @[:@47652.4]
  input  [63:0] io_ins_358, // @[:@47652.4]
  input  [63:0] io_ins_359, // @[:@47652.4]
  input  [63:0] io_ins_360, // @[:@47652.4]
  input  [63:0] io_ins_361, // @[:@47652.4]
  input  [63:0] io_ins_362, // @[:@47652.4]
  input  [63:0] io_ins_363, // @[:@47652.4]
  input  [63:0] io_ins_364, // @[:@47652.4]
  input  [63:0] io_ins_365, // @[:@47652.4]
  input  [63:0] io_ins_366, // @[:@47652.4]
  input  [63:0] io_ins_367, // @[:@47652.4]
  input  [63:0] io_ins_368, // @[:@47652.4]
  input  [63:0] io_ins_369, // @[:@47652.4]
  input  [63:0] io_ins_370, // @[:@47652.4]
  input  [63:0] io_ins_371, // @[:@47652.4]
  input  [63:0] io_ins_372, // @[:@47652.4]
  input  [63:0] io_ins_373, // @[:@47652.4]
  input  [63:0] io_ins_374, // @[:@47652.4]
  input  [63:0] io_ins_375, // @[:@47652.4]
  input  [63:0] io_ins_376, // @[:@47652.4]
  input  [63:0] io_ins_377, // @[:@47652.4]
  input  [63:0] io_ins_378, // @[:@47652.4]
  input  [63:0] io_ins_379, // @[:@47652.4]
  input  [63:0] io_ins_380, // @[:@47652.4]
  input  [63:0] io_ins_381, // @[:@47652.4]
  input  [63:0] io_ins_382, // @[:@47652.4]
  input  [63:0] io_ins_383, // @[:@47652.4]
  input  [63:0] io_ins_384, // @[:@47652.4]
  input  [63:0] io_ins_385, // @[:@47652.4]
  input  [63:0] io_ins_386, // @[:@47652.4]
  input  [63:0] io_ins_387, // @[:@47652.4]
  input  [63:0] io_ins_388, // @[:@47652.4]
  input  [63:0] io_ins_389, // @[:@47652.4]
  input  [63:0] io_ins_390, // @[:@47652.4]
  input  [63:0] io_ins_391, // @[:@47652.4]
  input  [63:0] io_ins_392, // @[:@47652.4]
  input  [63:0] io_ins_393, // @[:@47652.4]
  input  [63:0] io_ins_394, // @[:@47652.4]
  input  [63:0] io_ins_395, // @[:@47652.4]
  input  [63:0] io_ins_396, // @[:@47652.4]
  input  [63:0] io_ins_397, // @[:@47652.4]
  input  [63:0] io_ins_398, // @[:@47652.4]
  input  [63:0] io_ins_399, // @[:@47652.4]
  input  [63:0] io_ins_400, // @[:@47652.4]
  input  [63:0] io_ins_401, // @[:@47652.4]
  input  [63:0] io_ins_402, // @[:@47652.4]
  input  [63:0] io_ins_403, // @[:@47652.4]
  input  [63:0] io_ins_404, // @[:@47652.4]
  input  [63:0] io_ins_405, // @[:@47652.4]
  input  [63:0] io_ins_406, // @[:@47652.4]
  input  [63:0] io_ins_407, // @[:@47652.4]
  input  [63:0] io_ins_408, // @[:@47652.4]
  input  [63:0] io_ins_409, // @[:@47652.4]
  input  [63:0] io_ins_410, // @[:@47652.4]
  input  [63:0] io_ins_411, // @[:@47652.4]
  input  [63:0] io_ins_412, // @[:@47652.4]
  input  [63:0] io_ins_413, // @[:@47652.4]
  input  [63:0] io_ins_414, // @[:@47652.4]
  input  [63:0] io_ins_415, // @[:@47652.4]
  input  [63:0] io_ins_416, // @[:@47652.4]
  input  [63:0] io_ins_417, // @[:@47652.4]
  input  [63:0] io_ins_418, // @[:@47652.4]
  input  [63:0] io_ins_419, // @[:@47652.4]
  input  [63:0] io_ins_420, // @[:@47652.4]
  input  [63:0] io_ins_421, // @[:@47652.4]
  input  [63:0] io_ins_422, // @[:@47652.4]
  input  [63:0] io_ins_423, // @[:@47652.4]
  input  [63:0] io_ins_424, // @[:@47652.4]
  input  [63:0] io_ins_425, // @[:@47652.4]
  input  [63:0] io_ins_426, // @[:@47652.4]
  input  [63:0] io_ins_427, // @[:@47652.4]
  input  [63:0] io_ins_428, // @[:@47652.4]
  input  [63:0] io_ins_429, // @[:@47652.4]
  input  [63:0] io_ins_430, // @[:@47652.4]
  input  [63:0] io_ins_431, // @[:@47652.4]
  input  [63:0] io_ins_432, // @[:@47652.4]
  input  [63:0] io_ins_433, // @[:@47652.4]
  input  [63:0] io_ins_434, // @[:@47652.4]
  input  [63:0] io_ins_435, // @[:@47652.4]
  input  [63:0] io_ins_436, // @[:@47652.4]
  input  [63:0] io_ins_437, // @[:@47652.4]
  input  [63:0] io_ins_438, // @[:@47652.4]
  input  [63:0] io_ins_439, // @[:@47652.4]
  input  [63:0] io_ins_440, // @[:@47652.4]
  input  [63:0] io_ins_441, // @[:@47652.4]
  input  [63:0] io_ins_442, // @[:@47652.4]
  input  [63:0] io_ins_443, // @[:@47652.4]
  input  [63:0] io_ins_444, // @[:@47652.4]
  input  [63:0] io_ins_445, // @[:@47652.4]
  input  [63:0] io_ins_446, // @[:@47652.4]
  input  [63:0] io_ins_447, // @[:@47652.4]
  input  [63:0] io_ins_448, // @[:@47652.4]
  input  [63:0] io_ins_449, // @[:@47652.4]
  input  [63:0] io_ins_450, // @[:@47652.4]
  input  [63:0] io_ins_451, // @[:@47652.4]
  input  [63:0] io_ins_452, // @[:@47652.4]
  input  [63:0] io_ins_453, // @[:@47652.4]
  input  [63:0] io_ins_454, // @[:@47652.4]
  input  [63:0] io_ins_455, // @[:@47652.4]
  input  [63:0] io_ins_456, // @[:@47652.4]
  input  [63:0] io_ins_457, // @[:@47652.4]
  input  [63:0] io_ins_458, // @[:@47652.4]
  input  [63:0] io_ins_459, // @[:@47652.4]
  input  [63:0] io_ins_460, // @[:@47652.4]
  input  [63:0] io_ins_461, // @[:@47652.4]
  input  [63:0] io_ins_462, // @[:@47652.4]
  input  [63:0] io_ins_463, // @[:@47652.4]
  input  [63:0] io_ins_464, // @[:@47652.4]
  input  [63:0] io_ins_465, // @[:@47652.4]
  input  [63:0] io_ins_466, // @[:@47652.4]
  input  [63:0] io_ins_467, // @[:@47652.4]
  input  [63:0] io_ins_468, // @[:@47652.4]
  input  [63:0] io_ins_469, // @[:@47652.4]
  input  [63:0] io_ins_470, // @[:@47652.4]
  input  [63:0] io_ins_471, // @[:@47652.4]
  input  [63:0] io_ins_472, // @[:@47652.4]
  input  [63:0] io_ins_473, // @[:@47652.4]
  input  [63:0] io_ins_474, // @[:@47652.4]
  input  [63:0] io_ins_475, // @[:@47652.4]
  input  [63:0] io_ins_476, // @[:@47652.4]
  input  [63:0] io_ins_477, // @[:@47652.4]
  input  [63:0] io_ins_478, // @[:@47652.4]
  input  [63:0] io_ins_479, // @[:@47652.4]
  input  [63:0] io_ins_480, // @[:@47652.4]
  input  [63:0] io_ins_481, // @[:@47652.4]
  input  [63:0] io_ins_482, // @[:@47652.4]
  input  [63:0] io_ins_483, // @[:@47652.4]
  input  [63:0] io_ins_484, // @[:@47652.4]
  input  [63:0] io_ins_485, // @[:@47652.4]
  input  [63:0] io_ins_486, // @[:@47652.4]
  input  [63:0] io_ins_487, // @[:@47652.4]
  input  [63:0] io_ins_488, // @[:@47652.4]
  input  [63:0] io_ins_489, // @[:@47652.4]
  input  [63:0] io_ins_490, // @[:@47652.4]
  input  [63:0] io_ins_491, // @[:@47652.4]
  input  [63:0] io_ins_492, // @[:@47652.4]
  input  [63:0] io_ins_493, // @[:@47652.4]
  input  [63:0] io_ins_494, // @[:@47652.4]
  input  [63:0] io_ins_495, // @[:@47652.4]
  input  [63:0] io_ins_496, // @[:@47652.4]
  input  [63:0] io_ins_497, // @[:@47652.4]
  input  [63:0] io_ins_498, // @[:@47652.4]
  input  [63:0] io_ins_499, // @[:@47652.4]
  input  [63:0] io_ins_500, // @[:@47652.4]
  input  [63:0] io_ins_501, // @[:@47652.4]
  input  [63:0] io_ins_502, // @[:@47652.4]
  input  [63:0] io_ins_503, // @[:@47652.4]
  input  [63:0] io_ins_504, // @[:@47652.4]
  input  [63:0] io_ins_505, // @[:@47652.4]
  input  [63:0] io_ins_506, // @[:@47652.4]
  input  [63:0] io_ins_507, // @[:@47652.4]
  input  [63:0] io_ins_508, // @[:@47652.4]
  input  [63:0] io_ins_509, // @[:@47652.4]
  input  [63:0] io_ins_510, // @[:@47652.4]
  input  [63:0] io_ins_511, // @[:@47652.4]
  input  [63:0] io_ins_512, // @[:@47652.4]
  input  [63:0] io_ins_513, // @[:@47652.4]
  input  [63:0] io_ins_514, // @[:@47652.4]
  input  [63:0] io_ins_515, // @[:@47652.4]
  input  [63:0] io_ins_516, // @[:@47652.4]
  input  [63:0] io_ins_517, // @[:@47652.4]
  input  [9:0]  io_sel, // @[:@47652.4]
  output [63:0] io_out // @[:@47652.4]
);
  wire [63:0] _GEN_1; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_2; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_3; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_4; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_5; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_6; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_7; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_8; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_9; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_10; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_11; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_12; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_13; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_14; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_15; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_16; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_17; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_18; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_19; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_20; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_21; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_22; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_23; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_24; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_25; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_26; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_27; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_28; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_29; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_30; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_31; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_32; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_33; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_34; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_35; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_36; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_37; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_38; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_39; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_40; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_41; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_42; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_43; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_44; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_45; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_46; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_47; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_48; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_49; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_50; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_51; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_52; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_53; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_54; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_55; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_56; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_57; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_58; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_59; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_60; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_61; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_62; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_63; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_64; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_65; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_66; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_67; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_68; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_69; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_70; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_71; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_72; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_73; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_74; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_75; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_76; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_77; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_78; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_79; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_80; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_81; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_82; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_83; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_84; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_85; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_86; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_87; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_88; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_89; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_90; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_91; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_92; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_93; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_94; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_95; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_96; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_97; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_98; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_99; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_100; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_101; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_102; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_103; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_104; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_105; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_106; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_107; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_108; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_109; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_110; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_111; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_112; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_113; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_114; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_115; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_116; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_117; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_118; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_119; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_120; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_121; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_122; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_123; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_124; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_125; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_126; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_127; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_128; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_129; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_130; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_131; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_132; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_133; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_134; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_135; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_136; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_137; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_138; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_139; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_140; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_141; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_142; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_143; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_144; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_145; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_146; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_147; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_148; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_149; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_150; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_151; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_152; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_153; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_154; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_155; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_156; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_157; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_158; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_159; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_160; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_161; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_162; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_163; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_164; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_165; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_166; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_167; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_168; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_169; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_170; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_171; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_172; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_173; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_174; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_175; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_176; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_177; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_178; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_179; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_180; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_181; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_182; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_183; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_184; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_185; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_186; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_187; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_188; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_189; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_190; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_191; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_192; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_193; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_194; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_195; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_196; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_197; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_198; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_199; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_200; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_201; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_202; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_203; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_204; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_205; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_206; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_207; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_208; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_209; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_210; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_211; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_212; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_213; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_214; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_215; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_216; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_217; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_218; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_219; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_220; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_221; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_222; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_223; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_224; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_225; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_226; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_227; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_228; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_229; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_230; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_231; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_232; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_233; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_234; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_235; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_236; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_237; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_238; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_239; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_240; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_241; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_242; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_243; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_244; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_245; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_246; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_247; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_248; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_249; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_250; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_251; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_252; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_253; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_254; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_255; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_256; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_257; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_258; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_259; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_260; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_261; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_262; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_263; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_264; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_265; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_266; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_267; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_268; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_269; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_270; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_271; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_272; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_273; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_274; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_275; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_276; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_277; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_278; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_279; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_280; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_281; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_282; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_283; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_284; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_285; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_286; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_287; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_288; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_289; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_290; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_291; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_292; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_293; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_294; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_295; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_296; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_297; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_298; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_299; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_300; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_301; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_302; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_303; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_304; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_305; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_306; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_307; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_308; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_309; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_310; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_311; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_312; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_313; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_314; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_315; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_316; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_317; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_318; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_319; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_320; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_321; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_322; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_323; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_324; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_325; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_326; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_327; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_328; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_329; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_330; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_331; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_332; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_333; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_334; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_335; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_336; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_337; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_338; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_339; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_340; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_341; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_342; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_343; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_344; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_345; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_346; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_347; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_348; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_349; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_350; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_351; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_352; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_353; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_354; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_355; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_356; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_357; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_358; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_359; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_360; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_361; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_362; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_363; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_364; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_365; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_366; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_367; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_368; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_369; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_370; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_371; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_372; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_373; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_374; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_375; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_376; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_377; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_378; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_379; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_380; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_381; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_382; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_383; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_384; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_385; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_386; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_387; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_388; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_389; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_390; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_391; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_392; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_393; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_394; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_395; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_396; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_397; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_398; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_399; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_400; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_401; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_402; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_403; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_404; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_405; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_406; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_407; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_408; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_409; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_410; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_411; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_412; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_413; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_414; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_415; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_416; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_417; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_418; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_419; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_420; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_421; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_422; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_423; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_424; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_425; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_426; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_427; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_428; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_429; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_430; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_431; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_432; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_433; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_434; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_435; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_436; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_437; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_438; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_439; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_440; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_441; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_442; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_443; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_444; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_445; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_446; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_447; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_448; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_449; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_450; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_451; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_452; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_453; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_454; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_455; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_456; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_457; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_458; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_459; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_460; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_461; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_462; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_463; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_464; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_465; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_466; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_467; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_468; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_469; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_470; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_471; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_472; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_473; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_474; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_475; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_476; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_477; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_478; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_479; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_480; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_481; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_482; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_483; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_484; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_485; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_486; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_487; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_488; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_489; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_490; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_491; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_492; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_493; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_494; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_495; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_496; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_497; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_498; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_499; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_500; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_501; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_502; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_503; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_504; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_505; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_506; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_507; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_508; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_509; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_510; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_511; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_512; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_513; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_514; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_515; // @[MuxN.scala 16:10:@47654.4]
  wire [63:0] _GEN_516; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_1 = 10'h1 == io_sel ? io_ins_1 : io_ins_0; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_2 = 10'h2 == io_sel ? io_ins_2 : _GEN_1; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_3 = 10'h3 == io_sel ? io_ins_3 : _GEN_2; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_4 = 10'h4 == io_sel ? io_ins_4 : _GEN_3; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_5 = 10'h5 == io_sel ? io_ins_5 : _GEN_4; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_6 = 10'h6 == io_sel ? io_ins_6 : _GEN_5; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_7 = 10'h7 == io_sel ? io_ins_7 : _GEN_6; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_8 = 10'h8 == io_sel ? io_ins_8 : _GEN_7; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_9 = 10'h9 == io_sel ? io_ins_9 : _GEN_8; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_10 = 10'ha == io_sel ? io_ins_10 : _GEN_9; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_11 = 10'hb == io_sel ? io_ins_11 : _GEN_10; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_12 = 10'hc == io_sel ? io_ins_12 : _GEN_11; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_13 = 10'hd == io_sel ? io_ins_13 : _GEN_12; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_14 = 10'he == io_sel ? io_ins_14 : _GEN_13; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_15 = 10'hf == io_sel ? io_ins_15 : _GEN_14; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_16 = 10'h10 == io_sel ? io_ins_16 : _GEN_15; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_17 = 10'h11 == io_sel ? io_ins_17 : _GEN_16; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_18 = 10'h12 == io_sel ? io_ins_18 : _GEN_17; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_19 = 10'h13 == io_sel ? io_ins_19 : _GEN_18; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_20 = 10'h14 == io_sel ? io_ins_20 : _GEN_19; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_21 = 10'h15 == io_sel ? io_ins_21 : _GEN_20; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_22 = 10'h16 == io_sel ? io_ins_22 : _GEN_21; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_23 = 10'h17 == io_sel ? io_ins_23 : _GEN_22; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_24 = 10'h18 == io_sel ? io_ins_24 : _GEN_23; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_25 = 10'h19 == io_sel ? io_ins_25 : _GEN_24; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_26 = 10'h1a == io_sel ? io_ins_26 : _GEN_25; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_27 = 10'h1b == io_sel ? io_ins_27 : _GEN_26; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_28 = 10'h1c == io_sel ? io_ins_28 : _GEN_27; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_29 = 10'h1d == io_sel ? io_ins_29 : _GEN_28; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_30 = 10'h1e == io_sel ? io_ins_30 : _GEN_29; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_31 = 10'h1f == io_sel ? io_ins_31 : _GEN_30; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_32 = 10'h20 == io_sel ? io_ins_32 : _GEN_31; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_33 = 10'h21 == io_sel ? io_ins_33 : _GEN_32; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_34 = 10'h22 == io_sel ? io_ins_34 : _GEN_33; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_35 = 10'h23 == io_sel ? io_ins_35 : _GEN_34; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_36 = 10'h24 == io_sel ? io_ins_36 : _GEN_35; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_37 = 10'h25 == io_sel ? io_ins_37 : _GEN_36; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_38 = 10'h26 == io_sel ? io_ins_38 : _GEN_37; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_39 = 10'h27 == io_sel ? io_ins_39 : _GEN_38; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_40 = 10'h28 == io_sel ? io_ins_40 : _GEN_39; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_41 = 10'h29 == io_sel ? io_ins_41 : _GEN_40; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_42 = 10'h2a == io_sel ? io_ins_42 : _GEN_41; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_43 = 10'h2b == io_sel ? io_ins_43 : _GEN_42; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_44 = 10'h2c == io_sel ? io_ins_44 : _GEN_43; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_45 = 10'h2d == io_sel ? io_ins_45 : _GEN_44; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_46 = 10'h2e == io_sel ? io_ins_46 : _GEN_45; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_47 = 10'h2f == io_sel ? io_ins_47 : _GEN_46; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_48 = 10'h30 == io_sel ? io_ins_48 : _GEN_47; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_49 = 10'h31 == io_sel ? io_ins_49 : _GEN_48; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_50 = 10'h32 == io_sel ? io_ins_50 : _GEN_49; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_51 = 10'h33 == io_sel ? io_ins_51 : _GEN_50; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_52 = 10'h34 == io_sel ? io_ins_52 : _GEN_51; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_53 = 10'h35 == io_sel ? io_ins_53 : _GEN_52; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_54 = 10'h36 == io_sel ? io_ins_54 : _GEN_53; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_55 = 10'h37 == io_sel ? io_ins_55 : _GEN_54; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_56 = 10'h38 == io_sel ? io_ins_56 : _GEN_55; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_57 = 10'h39 == io_sel ? io_ins_57 : _GEN_56; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_58 = 10'h3a == io_sel ? io_ins_58 : _GEN_57; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_59 = 10'h3b == io_sel ? io_ins_59 : _GEN_58; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_60 = 10'h3c == io_sel ? io_ins_60 : _GEN_59; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_61 = 10'h3d == io_sel ? io_ins_61 : _GEN_60; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_62 = 10'h3e == io_sel ? io_ins_62 : _GEN_61; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_63 = 10'h3f == io_sel ? io_ins_63 : _GEN_62; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_64 = 10'h40 == io_sel ? io_ins_64 : _GEN_63; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_65 = 10'h41 == io_sel ? io_ins_65 : _GEN_64; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_66 = 10'h42 == io_sel ? io_ins_66 : _GEN_65; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_67 = 10'h43 == io_sel ? io_ins_67 : _GEN_66; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_68 = 10'h44 == io_sel ? io_ins_68 : _GEN_67; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_69 = 10'h45 == io_sel ? io_ins_69 : _GEN_68; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_70 = 10'h46 == io_sel ? io_ins_70 : _GEN_69; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_71 = 10'h47 == io_sel ? io_ins_71 : _GEN_70; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_72 = 10'h48 == io_sel ? io_ins_72 : _GEN_71; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_73 = 10'h49 == io_sel ? io_ins_73 : _GEN_72; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_74 = 10'h4a == io_sel ? io_ins_74 : _GEN_73; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_75 = 10'h4b == io_sel ? io_ins_75 : _GEN_74; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_76 = 10'h4c == io_sel ? io_ins_76 : _GEN_75; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_77 = 10'h4d == io_sel ? io_ins_77 : _GEN_76; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_78 = 10'h4e == io_sel ? io_ins_78 : _GEN_77; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_79 = 10'h4f == io_sel ? io_ins_79 : _GEN_78; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_80 = 10'h50 == io_sel ? io_ins_80 : _GEN_79; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_81 = 10'h51 == io_sel ? io_ins_81 : _GEN_80; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_82 = 10'h52 == io_sel ? io_ins_82 : _GEN_81; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_83 = 10'h53 == io_sel ? io_ins_83 : _GEN_82; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_84 = 10'h54 == io_sel ? io_ins_84 : _GEN_83; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_85 = 10'h55 == io_sel ? io_ins_85 : _GEN_84; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_86 = 10'h56 == io_sel ? io_ins_86 : _GEN_85; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_87 = 10'h57 == io_sel ? io_ins_87 : _GEN_86; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_88 = 10'h58 == io_sel ? io_ins_88 : _GEN_87; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_89 = 10'h59 == io_sel ? io_ins_89 : _GEN_88; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_90 = 10'h5a == io_sel ? io_ins_90 : _GEN_89; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_91 = 10'h5b == io_sel ? io_ins_91 : _GEN_90; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_92 = 10'h5c == io_sel ? io_ins_92 : _GEN_91; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_93 = 10'h5d == io_sel ? io_ins_93 : _GEN_92; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_94 = 10'h5e == io_sel ? io_ins_94 : _GEN_93; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_95 = 10'h5f == io_sel ? io_ins_95 : _GEN_94; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_96 = 10'h60 == io_sel ? io_ins_96 : _GEN_95; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_97 = 10'h61 == io_sel ? io_ins_97 : _GEN_96; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_98 = 10'h62 == io_sel ? io_ins_98 : _GEN_97; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_99 = 10'h63 == io_sel ? io_ins_99 : _GEN_98; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_100 = 10'h64 == io_sel ? io_ins_100 : _GEN_99; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_101 = 10'h65 == io_sel ? io_ins_101 : _GEN_100; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_102 = 10'h66 == io_sel ? io_ins_102 : _GEN_101; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_103 = 10'h67 == io_sel ? io_ins_103 : _GEN_102; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_104 = 10'h68 == io_sel ? io_ins_104 : _GEN_103; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_105 = 10'h69 == io_sel ? io_ins_105 : _GEN_104; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_106 = 10'h6a == io_sel ? io_ins_106 : _GEN_105; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_107 = 10'h6b == io_sel ? io_ins_107 : _GEN_106; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_108 = 10'h6c == io_sel ? io_ins_108 : _GEN_107; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_109 = 10'h6d == io_sel ? io_ins_109 : _GEN_108; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_110 = 10'h6e == io_sel ? io_ins_110 : _GEN_109; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_111 = 10'h6f == io_sel ? io_ins_111 : _GEN_110; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_112 = 10'h70 == io_sel ? io_ins_112 : _GEN_111; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_113 = 10'h71 == io_sel ? io_ins_113 : _GEN_112; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_114 = 10'h72 == io_sel ? io_ins_114 : _GEN_113; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_115 = 10'h73 == io_sel ? io_ins_115 : _GEN_114; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_116 = 10'h74 == io_sel ? io_ins_116 : _GEN_115; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_117 = 10'h75 == io_sel ? io_ins_117 : _GEN_116; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_118 = 10'h76 == io_sel ? io_ins_118 : _GEN_117; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_119 = 10'h77 == io_sel ? io_ins_119 : _GEN_118; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_120 = 10'h78 == io_sel ? io_ins_120 : _GEN_119; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_121 = 10'h79 == io_sel ? io_ins_121 : _GEN_120; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_122 = 10'h7a == io_sel ? io_ins_122 : _GEN_121; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_123 = 10'h7b == io_sel ? io_ins_123 : _GEN_122; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_124 = 10'h7c == io_sel ? io_ins_124 : _GEN_123; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_125 = 10'h7d == io_sel ? io_ins_125 : _GEN_124; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_126 = 10'h7e == io_sel ? io_ins_126 : _GEN_125; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_127 = 10'h7f == io_sel ? io_ins_127 : _GEN_126; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_128 = 10'h80 == io_sel ? io_ins_128 : _GEN_127; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_129 = 10'h81 == io_sel ? io_ins_129 : _GEN_128; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_130 = 10'h82 == io_sel ? io_ins_130 : _GEN_129; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_131 = 10'h83 == io_sel ? io_ins_131 : _GEN_130; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_132 = 10'h84 == io_sel ? io_ins_132 : _GEN_131; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_133 = 10'h85 == io_sel ? io_ins_133 : _GEN_132; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_134 = 10'h86 == io_sel ? io_ins_134 : _GEN_133; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_135 = 10'h87 == io_sel ? io_ins_135 : _GEN_134; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_136 = 10'h88 == io_sel ? io_ins_136 : _GEN_135; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_137 = 10'h89 == io_sel ? io_ins_137 : _GEN_136; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_138 = 10'h8a == io_sel ? io_ins_138 : _GEN_137; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_139 = 10'h8b == io_sel ? io_ins_139 : _GEN_138; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_140 = 10'h8c == io_sel ? io_ins_140 : _GEN_139; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_141 = 10'h8d == io_sel ? io_ins_141 : _GEN_140; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_142 = 10'h8e == io_sel ? io_ins_142 : _GEN_141; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_143 = 10'h8f == io_sel ? io_ins_143 : _GEN_142; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_144 = 10'h90 == io_sel ? io_ins_144 : _GEN_143; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_145 = 10'h91 == io_sel ? io_ins_145 : _GEN_144; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_146 = 10'h92 == io_sel ? io_ins_146 : _GEN_145; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_147 = 10'h93 == io_sel ? io_ins_147 : _GEN_146; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_148 = 10'h94 == io_sel ? io_ins_148 : _GEN_147; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_149 = 10'h95 == io_sel ? io_ins_149 : _GEN_148; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_150 = 10'h96 == io_sel ? io_ins_150 : _GEN_149; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_151 = 10'h97 == io_sel ? io_ins_151 : _GEN_150; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_152 = 10'h98 == io_sel ? io_ins_152 : _GEN_151; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_153 = 10'h99 == io_sel ? io_ins_153 : _GEN_152; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_154 = 10'h9a == io_sel ? io_ins_154 : _GEN_153; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_155 = 10'h9b == io_sel ? io_ins_155 : _GEN_154; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_156 = 10'h9c == io_sel ? io_ins_156 : _GEN_155; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_157 = 10'h9d == io_sel ? io_ins_157 : _GEN_156; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_158 = 10'h9e == io_sel ? io_ins_158 : _GEN_157; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_159 = 10'h9f == io_sel ? io_ins_159 : _GEN_158; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_160 = 10'ha0 == io_sel ? io_ins_160 : _GEN_159; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_161 = 10'ha1 == io_sel ? io_ins_161 : _GEN_160; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_162 = 10'ha2 == io_sel ? io_ins_162 : _GEN_161; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_163 = 10'ha3 == io_sel ? io_ins_163 : _GEN_162; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_164 = 10'ha4 == io_sel ? io_ins_164 : _GEN_163; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_165 = 10'ha5 == io_sel ? io_ins_165 : _GEN_164; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_166 = 10'ha6 == io_sel ? io_ins_166 : _GEN_165; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_167 = 10'ha7 == io_sel ? io_ins_167 : _GEN_166; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_168 = 10'ha8 == io_sel ? io_ins_168 : _GEN_167; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_169 = 10'ha9 == io_sel ? io_ins_169 : _GEN_168; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_170 = 10'haa == io_sel ? io_ins_170 : _GEN_169; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_171 = 10'hab == io_sel ? io_ins_171 : _GEN_170; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_172 = 10'hac == io_sel ? io_ins_172 : _GEN_171; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_173 = 10'had == io_sel ? io_ins_173 : _GEN_172; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_174 = 10'hae == io_sel ? io_ins_174 : _GEN_173; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_175 = 10'haf == io_sel ? io_ins_175 : _GEN_174; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_176 = 10'hb0 == io_sel ? io_ins_176 : _GEN_175; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_177 = 10'hb1 == io_sel ? io_ins_177 : _GEN_176; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_178 = 10'hb2 == io_sel ? io_ins_178 : _GEN_177; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_179 = 10'hb3 == io_sel ? io_ins_179 : _GEN_178; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_180 = 10'hb4 == io_sel ? io_ins_180 : _GEN_179; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_181 = 10'hb5 == io_sel ? io_ins_181 : _GEN_180; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_182 = 10'hb6 == io_sel ? io_ins_182 : _GEN_181; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_183 = 10'hb7 == io_sel ? io_ins_183 : _GEN_182; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_184 = 10'hb8 == io_sel ? io_ins_184 : _GEN_183; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_185 = 10'hb9 == io_sel ? io_ins_185 : _GEN_184; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_186 = 10'hba == io_sel ? io_ins_186 : _GEN_185; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_187 = 10'hbb == io_sel ? io_ins_187 : _GEN_186; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_188 = 10'hbc == io_sel ? io_ins_188 : _GEN_187; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_189 = 10'hbd == io_sel ? io_ins_189 : _GEN_188; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_190 = 10'hbe == io_sel ? io_ins_190 : _GEN_189; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_191 = 10'hbf == io_sel ? io_ins_191 : _GEN_190; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_192 = 10'hc0 == io_sel ? io_ins_192 : _GEN_191; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_193 = 10'hc1 == io_sel ? io_ins_193 : _GEN_192; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_194 = 10'hc2 == io_sel ? io_ins_194 : _GEN_193; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_195 = 10'hc3 == io_sel ? io_ins_195 : _GEN_194; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_196 = 10'hc4 == io_sel ? io_ins_196 : _GEN_195; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_197 = 10'hc5 == io_sel ? io_ins_197 : _GEN_196; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_198 = 10'hc6 == io_sel ? io_ins_198 : _GEN_197; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_199 = 10'hc7 == io_sel ? io_ins_199 : _GEN_198; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_200 = 10'hc8 == io_sel ? io_ins_200 : _GEN_199; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_201 = 10'hc9 == io_sel ? io_ins_201 : _GEN_200; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_202 = 10'hca == io_sel ? io_ins_202 : _GEN_201; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_203 = 10'hcb == io_sel ? io_ins_203 : _GEN_202; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_204 = 10'hcc == io_sel ? io_ins_204 : _GEN_203; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_205 = 10'hcd == io_sel ? io_ins_205 : _GEN_204; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_206 = 10'hce == io_sel ? io_ins_206 : _GEN_205; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_207 = 10'hcf == io_sel ? io_ins_207 : _GEN_206; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_208 = 10'hd0 == io_sel ? io_ins_208 : _GEN_207; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_209 = 10'hd1 == io_sel ? io_ins_209 : _GEN_208; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_210 = 10'hd2 == io_sel ? io_ins_210 : _GEN_209; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_211 = 10'hd3 == io_sel ? io_ins_211 : _GEN_210; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_212 = 10'hd4 == io_sel ? io_ins_212 : _GEN_211; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_213 = 10'hd5 == io_sel ? io_ins_213 : _GEN_212; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_214 = 10'hd6 == io_sel ? io_ins_214 : _GEN_213; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_215 = 10'hd7 == io_sel ? io_ins_215 : _GEN_214; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_216 = 10'hd8 == io_sel ? io_ins_216 : _GEN_215; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_217 = 10'hd9 == io_sel ? io_ins_217 : _GEN_216; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_218 = 10'hda == io_sel ? io_ins_218 : _GEN_217; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_219 = 10'hdb == io_sel ? io_ins_219 : _GEN_218; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_220 = 10'hdc == io_sel ? io_ins_220 : _GEN_219; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_221 = 10'hdd == io_sel ? io_ins_221 : _GEN_220; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_222 = 10'hde == io_sel ? io_ins_222 : _GEN_221; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_223 = 10'hdf == io_sel ? io_ins_223 : _GEN_222; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_224 = 10'he0 == io_sel ? io_ins_224 : _GEN_223; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_225 = 10'he1 == io_sel ? io_ins_225 : _GEN_224; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_226 = 10'he2 == io_sel ? io_ins_226 : _GEN_225; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_227 = 10'he3 == io_sel ? io_ins_227 : _GEN_226; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_228 = 10'he4 == io_sel ? io_ins_228 : _GEN_227; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_229 = 10'he5 == io_sel ? io_ins_229 : _GEN_228; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_230 = 10'he6 == io_sel ? io_ins_230 : _GEN_229; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_231 = 10'he7 == io_sel ? io_ins_231 : _GEN_230; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_232 = 10'he8 == io_sel ? io_ins_232 : _GEN_231; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_233 = 10'he9 == io_sel ? io_ins_233 : _GEN_232; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_234 = 10'hea == io_sel ? io_ins_234 : _GEN_233; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_235 = 10'heb == io_sel ? io_ins_235 : _GEN_234; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_236 = 10'hec == io_sel ? io_ins_236 : _GEN_235; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_237 = 10'hed == io_sel ? io_ins_237 : _GEN_236; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_238 = 10'hee == io_sel ? io_ins_238 : _GEN_237; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_239 = 10'hef == io_sel ? io_ins_239 : _GEN_238; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_240 = 10'hf0 == io_sel ? io_ins_240 : _GEN_239; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_241 = 10'hf1 == io_sel ? io_ins_241 : _GEN_240; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_242 = 10'hf2 == io_sel ? io_ins_242 : _GEN_241; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_243 = 10'hf3 == io_sel ? io_ins_243 : _GEN_242; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_244 = 10'hf4 == io_sel ? io_ins_244 : _GEN_243; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_245 = 10'hf5 == io_sel ? io_ins_245 : _GEN_244; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_246 = 10'hf6 == io_sel ? io_ins_246 : _GEN_245; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_247 = 10'hf7 == io_sel ? io_ins_247 : _GEN_246; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_248 = 10'hf8 == io_sel ? io_ins_248 : _GEN_247; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_249 = 10'hf9 == io_sel ? io_ins_249 : _GEN_248; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_250 = 10'hfa == io_sel ? io_ins_250 : _GEN_249; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_251 = 10'hfb == io_sel ? io_ins_251 : _GEN_250; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_252 = 10'hfc == io_sel ? io_ins_252 : _GEN_251; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_253 = 10'hfd == io_sel ? io_ins_253 : _GEN_252; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_254 = 10'hfe == io_sel ? io_ins_254 : _GEN_253; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_255 = 10'hff == io_sel ? io_ins_255 : _GEN_254; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_256 = 10'h100 == io_sel ? io_ins_256 : _GEN_255; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_257 = 10'h101 == io_sel ? io_ins_257 : _GEN_256; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_258 = 10'h102 == io_sel ? io_ins_258 : _GEN_257; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_259 = 10'h103 == io_sel ? io_ins_259 : _GEN_258; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_260 = 10'h104 == io_sel ? io_ins_260 : _GEN_259; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_261 = 10'h105 == io_sel ? io_ins_261 : _GEN_260; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_262 = 10'h106 == io_sel ? io_ins_262 : _GEN_261; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_263 = 10'h107 == io_sel ? io_ins_263 : _GEN_262; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_264 = 10'h108 == io_sel ? io_ins_264 : _GEN_263; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_265 = 10'h109 == io_sel ? io_ins_265 : _GEN_264; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_266 = 10'h10a == io_sel ? io_ins_266 : _GEN_265; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_267 = 10'h10b == io_sel ? io_ins_267 : _GEN_266; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_268 = 10'h10c == io_sel ? io_ins_268 : _GEN_267; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_269 = 10'h10d == io_sel ? io_ins_269 : _GEN_268; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_270 = 10'h10e == io_sel ? io_ins_270 : _GEN_269; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_271 = 10'h10f == io_sel ? io_ins_271 : _GEN_270; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_272 = 10'h110 == io_sel ? io_ins_272 : _GEN_271; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_273 = 10'h111 == io_sel ? io_ins_273 : _GEN_272; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_274 = 10'h112 == io_sel ? io_ins_274 : _GEN_273; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_275 = 10'h113 == io_sel ? io_ins_275 : _GEN_274; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_276 = 10'h114 == io_sel ? io_ins_276 : _GEN_275; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_277 = 10'h115 == io_sel ? io_ins_277 : _GEN_276; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_278 = 10'h116 == io_sel ? io_ins_278 : _GEN_277; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_279 = 10'h117 == io_sel ? io_ins_279 : _GEN_278; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_280 = 10'h118 == io_sel ? io_ins_280 : _GEN_279; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_281 = 10'h119 == io_sel ? io_ins_281 : _GEN_280; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_282 = 10'h11a == io_sel ? io_ins_282 : _GEN_281; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_283 = 10'h11b == io_sel ? io_ins_283 : _GEN_282; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_284 = 10'h11c == io_sel ? io_ins_284 : _GEN_283; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_285 = 10'h11d == io_sel ? io_ins_285 : _GEN_284; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_286 = 10'h11e == io_sel ? io_ins_286 : _GEN_285; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_287 = 10'h11f == io_sel ? io_ins_287 : _GEN_286; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_288 = 10'h120 == io_sel ? io_ins_288 : _GEN_287; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_289 = 10'h121 == io_sel ? io_ins_289 : _GEN_288; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_290 = 10'h122 == io_sel ? io_ins_290 : _GEN_289; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_291 = 10'h123 == io_sel ? io_ins_291 : _GEN_290; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_292 = 10'h124 == io_sel ? io_ins_292 : _GEN_291; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_293 = 10'h125 == io_sel ? io_ins_293 : _GEN_292; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_294 = 10'h126 == io_sel ? io_ins_294 : _GEN_293; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_295 = 10'h127 == io_sel ? io_ins_295 : _GEN_294; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_296 = 10'h128 == io_sel ? io_ins_296 : _GEN_295; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_297 = 10'h129 == io_sel ? io_ins_297 : _GEN_296; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_298 = 10'h12a == io_sel ? io_ins_298 : _GEN_297; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_299 = 10'h12b == io_sel ? io_ins_299 : _GEN_298; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_300 = 10'h12c == io_sel ? io_ins_300 : _GEN_299; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_301 = 10'h12d == io_sel ? io_ins_301 : _GEN_300; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_302 = 10'h12e == io_sel ? io_ins_302 : _GEN_301; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_303 = 10'h12f == io_sel ? io_ins_303 : _GEN_302; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_304 = 10'h130 == io_sel ? io_ins_304 : _GEN_303; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_305 = 10'h131 == io_sel ? io_ins_305 : _GEN_304; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_306 = 10'h132 == io_sel ? io_ins_306 : _GEN_305; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_307 = 10'h133 == io_sel ? io_ins_307 : _GEN_306; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_308 = 10'h134 == io_sel ? io_ins_308 : _GEN_307; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_309 = 10'h135 == io_sel ? io_ins_309 : _GEN_308; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_310 = 10'h136 == io_sel ? io_ins_310 : _GEN_309; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_311 = 10'h137 == io_sel ? io_ins_311 : _GEN_310; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_312 = 10'h138 == io_sel ? io_ins_312 : _GEN_311; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_313 = 10'h139 == io_sel ? io_ins_313 : _GEN_312; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_314 = 10'h13a == io_sel ? io_ins_314 : _GEN_313; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_315 = 10'h13b == io_sel ? io_ins_315 : _GEN_314; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_316 = 10'h13c == io_sel ? io_ins_316 : _GEN_315; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_317 = 10'h13d == io_sel ? io_ins_317 : _GEN_316; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_318 = 10'h13e == io_sel ? io_ins_318 : _GEN_317; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_319 = 10'h13f == io_sel ? io_ins_319 : _GEN_318; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_320 = 10'h140 == io_sel ? io_ins_320 : _GEN_319; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_321 = 10'h141 == io_sel ? io_ins_321 : _GEN_320; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_322 = 10'h142 == io_sel ? io_ins_322 : _GEN_321; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_323 = 10'h143 == io_sel ? io_ins_323 : _GEN_322; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_324 = 10'h144 == io_sel ? io_ins_324 : _GEN_323; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_325 = 10'h145 == io_sel ? io_ins_325 : _GEN_324; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_326 = 10'h146 == io_sel ? io_ins_326 : _GEN_325; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_327 = 10'h147 == io_sel ? io_ins_327 : _GEN_326; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_328 = 10'h148 == io_sel ? io_ins_328 : _GEN_327; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_329 = 10'h149 == io_sel ? io_ins_329 : _GEN_328; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_330 = 10'h14a == io_sel ? io_ins_330 : _GEN_329; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_331 = 10'h14b == io_sel ? io_ins_331 : _GEN_330; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_332 = 10'h14c == io_sel ? io_ins_332 : _GEN_331; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_333 = 10'h14d == io_sel ? io_ins_333 : _GEN_332; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_334 = 10'h14e == io_sel ? io_ins_334 : _GEN_333; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_335 = 10'h14f == io_sel ? io_ins_335 : _GEN_334; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_336 = 10'h150 == io_sel ? io_ins_336 : _GEN_335; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_337 = 10'h151 == io_sel ? io_ins_337 : _GEN_336; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_338 = 10'h152 == io_sel ? io_ins_338 : _GEN_337; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_339 = 10'h153 == io_sel ? io_ins_339 : _GEN_338; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_340 = 10'h154 == io_sel ? io_ins_340 : _GEN_339; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_341 = 10'h155 == io_sel ? io_ins_341 : _GEN_340; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_342 = 10'h156 == io_sel ? io_ins_342 : _GEN_341; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_343 = 10'h157 == io_sel ? io_ins_343 : _GEN_342; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_344 = 10'h158 == io_sel ? io_ins_344 : _GEN_343; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_345 = 10'h159 == io_sel ? io_ins_345 : _GEN_344; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_346 = 10'h15a == io_sel ? io_ins_346 : _GEN_345; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_347 = 10'h15b == io_sel ? io_ins_347 : _GEN_346; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_348 = 10'h15c == io_sel ? io_ins_348 : _GEN_347; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_349 = 10'h15d == io_sel ? io_ins_349 : _GEN_348; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_350 = 10'h15e == io_sel ? io_ins_350 : _GEN_349; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_351 = 10'h15f == io_sel ? io_ins_351 : _GEN_350; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_352 = 10'h160 == io_sel ? io_ins_352 : _GEN_351; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_353 = 10'h161 == io_sel ? io_ins_353 : _GEN_352; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_354 = 10'h162 == io_sel ? io_ins_354 : _GEN_353; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_355 = 10'h163 == io_sel ? io_ins_355 : _GEN_354; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_356 = 10'h164 == io_sel ? io_ins_356 : _GEN_355; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_357 = 10'h165 == io_sel ? io_ins_357 : _GEN_356; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_358 = 10'h166 == io_sel ? io_ins_358 : _GEN_357; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_359 = 10'h167 == io_sel ? io_ins_359 : _GEN_358; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_360 = 10'h168 == io_sel ? io_ins_360 : _GEN_359; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_361 = 10'h169 == io_sel ? io_ins_361 : _GEN_360; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_362 = 10'h16a == io_sel ? io_ins_362 : _GEN_361; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_363 = 10'h16b == io_sel ? io_ins_363 : _GEN_362; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_364 = 10'h16c == io_sel ? io_ins_364 : _GEN_363; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_365 = 10'h16d == io_sel ? io_ins_365 : _GEN_364; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_366 = 10'h16e == io_sel ? io_ins_366 : _GEN_365; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_367 = 10'h16f == io_sel ? io_ins_367 : _GEN_366; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_368 = 10'h170 == io_sel ? io_ins_368 : _GEN_367; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_369 = 10'h171 == io_sel ? io_ins_369 : _GEN_368; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_370 = 10'h172 == io_sel ? io_ins_370 : _GEN_369; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_371 = 10'h173 == io_sel ? io_ins_371 : _GEN_370; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_372 = 10'h174 == io_sel ? io_ins_372 : _GEN_371; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_373 = 10'h175 == io_sel ? io_ins_373 : _GEN_372; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_374 = 10'h176 == io_sel ? io_ins_374 : _GEN_373; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_375 = 10'h177 == io_sel ? io_ins_375 : _GEN_374; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_376 = 10'h178 == io_sel ? io_ins_376 : _GEN_375; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_377 = 10'h179 == io_sel ? io_ins_377 : _GEN_376; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_378 = 10'h17a == io_sel ? io_ins_378 : _GEN_377; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_379 = 10'h17b == io_sel ? io_ins_379 : _GEN_378; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_380 = 10'h17c == io_sel ? io_ins_380 : _GEN_379; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_381 = 10'h17d == io_sel ? io_ins_381 : _GEN_380; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_382 = 10'h17e == io_sel ? io_ins_382 : _GEN_381; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_383 = 10'h17f == io_sel ? io_ins_383 : _GEN_382; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_384 = 10'h180 == io_sel ? io_ins_384 : _GEN_383; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_385 = 10'h181 == io_sel ? io_ins_385 : _GEN_384; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_386 = 10'h182 == io_sel ? io_ins_386 : _GEN_385; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_387 = 10'h183 == io_sel ? io_ins_387 : _GEN_386; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_388 = 10'h184 == io_sel ? io_ins_388 : _GEN_387; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_389 = 10'h185 == io_sel ? io_ins_389 : _GEN_388; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_390 = 10'h186 == io_sel ? io_ins_390 : _GEN_389; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_391 = 10'h187 == io_sel ? io_ins_391 : _GEN_390; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_392 = 10'h188 == io_sel ? io_ins_392 : _GEN_391; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_393 = 10'h189 == io_sel ? io_ins_393 : _GEN_392; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_394 = 10'h18a == io_sel ? io_ins_394 : _GEN_393; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_395 = 10'h18b == io_sel ? io_ins_395 : _GEN_394; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_396 = 10'h18c == io_sel ? io_ins_396 : _GEN_395; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_397 = 10'h18d == io_sel ? io_ins_397 : _GEN_396; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_398 = 10'h18e == io_sel ? io_ins_398 : _GEN_397; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_399 = 10'h18f == io_sel ? io_ins_399 : _GEN_398; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_400 = 10'h190 == io_sel ? io_ins_400 : _GEN_399; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_401 = 10'h191 == io_sel ? io_ins_401 : _GEN_400; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_402 = 10'h192 == io_sel ? io_ins_402 : _GEN_401; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_403 = 10'h193 == io_sel ? io_ins_403 : _GEN_402; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_404 = 10'h194 == io_sel ? io_ins_404 : _GEN_403; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_405 = 10'h195 == io_sel ? io_ins_405 : _GEN_404; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_406 = 10'h196 == io_sel ? io_ins_406 : _GEN_405; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_407 = 10'h197 == io_sel ? io_ins_407 : _GEN_406; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_408 = 10'h198 == io_sel ? io_ins_408 : _GEN_407; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_409 = 10'h199 == io_sel ? io_ins_409 : _GEN_408; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_410 = 10'h19a == io_sel ? io_ins_410 : _GEN_409; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_411 = 10'h19b == io_sel ? io_ins_411 : _GEN_410; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_412 = 10'h19c == io_sel ? io_ins_412 : _GEN_411; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_413 = 10'h19d == io_sel ? io_ins_413 : _GEN_412; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_414 = 10'h19e == io_sel ? io_ins_414 : _GEN_413; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_415 = 10'h19f == io_sel ? io_ins_415 : _GEN_414; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_416 = 10'h1a0 == io_sel ? io_ins_416 : _GEN_415; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_417 = 10'h1a1 == io_sel ? io_ins_417 : _GEN_416; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_418 = 10'h1a2 == io_sel ? io_ins_418 : _GEN_417; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_419 = 10'h1a3 == io_sel ? io_ins_419 : _GEN_418; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_420 = 10'h1a4 == io_sel ? io_ins_420 : _GEN_419; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_421 = 10'h1a5 == io_sel ? io_ins_421 : _GEN_420; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_422 = 10'h1a6 == io_sel ? io_ins_422 : _GEN_421; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_423 = 10'h1a7 == io_sel ? io_ins_423 : _GEN_422; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_424 = 10'h1a8 == io_sel ? io_ins_424 : _GEN_423; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_425 = 10'h1a9 == io_sel ? io_ins_425 : _GEN_424; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_426 = 10'h1aa == io_sel ? io_ins_426 : _GEN_425; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_427 = 10'h1ab == io_sel ? io_ins_427 : _GEN_426; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_428 = 10'h1ac == io_sel ? io_ins_428 : _GEN_427; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_429 = 10'h1ad == io_sel ? io_ins_429 : _GEN_428; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_430 = 10'h1ae == io_sel ? io_ins_430 : _GEN_429; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_431 = 10'h1af == io_sel ? io_ins_431 : _GEN_430; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_432 = 10'h1b0 == io_sel ? io_ins_432 : _GEN_431; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_433 = 10'h1b1 == io_sel ? io_ins_433 : _GEN_432; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_434 = 10'h1b2 == io_sel ? io_ins_434 : _GEN_433; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_435 = 10'h1b3 == io_sel ? io_ins_435 : _GEN_434; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_436 = 10'h1b4 == io_sel ? io_ins_436 : _GEN_435; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_437 = 10'h1b5 == io_sel ? io_ins_437 : _GEN_436; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_438 = 10'h1b6 == io_sel ? io_ins_438 : _GEN_437; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_439 = 10'h1b7 == io_sel ? io_ins_439 : _GEN_438; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_440 = 10'h1b8 == io_sel ? io_ins_440 : _GEN_439; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_441 = 10'h1b9 == io_sel ? io_ins_441 : _GEN_440; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_442 = 10'h1ba == io_sel ? io_ins_442 : _GEN_441; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_443 = 10'h1bb == io_sel ? io_ins_443 : _GEN_442; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_444 = 10'h1bc == io_sel ? io_ins_444 : _GEN_443; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_445 = 10'h1bd == io_sel ? io_ins_445 : _GEN_444; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_446 = 10'h1be == io_sel ? io_ins_446 : _GEN_445; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_447 = 10'h1bf == io_sel ? io_ins_447 : _GEN_446; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_448 = 10'h1c0 == io_sel ? io_ins_448 : _GEN_447; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_449 = 10'h1c1 == io_sel ? io_ins_449 : _GEN_448; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_450 = 10'h1c2 == io_sel ? io_ins_450 : _GEN_449; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_451 = 10'h1c3 == io_sel ? io_ins_451 : _GEN_450; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_452 = 10'h1c4 == io_sel ? io_ins_452 : _GEN_451; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_453 = 10'h1c5 == io_sel ? io_ins_453 : _GEN_452; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_454 = 10'h1c6 == io_sel ? io_ins_454 : _GEN_453; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_455 = 10'h1c7 == io_sel ? io_ins_455 : _GEN_454; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_456 = 10'h1c8 == io_sel ? io_ins_456 : _GEN_455; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_457 = 10'h1c9 == io_sel ? io_ins_457 : _GEN_456; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_458 = 10'h1ca == io_sel ? io_ins_458 : _GEN_457; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_459 = 10'h1cb == io_sel ? io_ins_459 : _GEN_458; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_460 = 10'h1cc == io_sel ? io_ins_460 : _GEN_459; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_461 = 10'h1cd == io_sel ? io_ins_461 : _GEN_460; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_462 = 10'h1ce == io_sel ? io_ins_462 : _GEN_461; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_463 = 10'h1cf == io_sel ? io_ins_463 : _GEN_462; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_464 = 10'h1d0 == io_sel ? io_ins_464 : _GEN_463; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_465 = 10'h1d1 == io_sel ? io_ins_465 : _GEN_464; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_466 = 10'h1d2 == io_sel ? io_ins_466 : _GEN_465; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_467 = 10'h1d3 == io_sel ? io_ins_467 : _GEN_466; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_468 = 10'h1d4 == io_sel ? io_ins_468 : _GEN_467; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_469 = 10'h1d5 == io_sel ? io_ins_469 : _GEN_468; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_470 = 10'h1d6 == io_sel ? io_ins_470 : _GEN_469; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_471 = 10'h1d7 == io_sel ? io_ins_471 : _GEN_470; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_472 = 10'h1d8 == io_sel ? io_ins_472 : _GEN_471; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_473 = 10'h1d9 == io_sel ? io_ins_473 : _GEN_472; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_474 = 10'h1da == io_sel ? io_ins_474 : _GEN_473; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_475 = 10'h1db == io_sel ? io_ins_475 : _GEN_474; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_476 = 10'h1dc == io_sel ? io_ins_476 : _GEN_475; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_477 = 10'h1dd == io_sel ? io_ins_477 : _GEN_476; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_478 = 10'h1de == io_sel ? io_ins_478 : _GEN_477; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_479 = 10'h1df == io_sel ? io_ins_479 : _GEN_478; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_480 = 10'h1e0 == io_sel ? io_ins_480 : _GEN_479; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_481 = 10'h1e1 == io_sel ? io_ins_481 : _GEN_480; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_482 = 10'h1e2 == io_sel ? io_ins_482 : _GEN_481; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_483 = 10'h1e3 == io_sel ? io_ins_483 : _GEN_482; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_484 = 10'h1e4 == io_sel ? io_ins_484 : _GEN_483; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_485 = 10'h1e5 == io_sel ? io_ins_485 : _GEN_484; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_486 = 10'h1e6 == io_sel ? io_ins_486 : _GEN_485; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_487 = 10'h1e7 == io_sel ? io_ins_487 : _GEN_486; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_488 = 10'h1e8 == io_sel ? io_ins_488 : _GEN_487; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_489 = 10'h1e9 == io_sel ? io_ins_489 : _GEN_488; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_490 = 10'h1ea == io_sel ? io_ins_490 : _GEN_489; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_491 = 10'h1eb == io_sel ? io_ins_491 : _GEN_490; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_492 = 10'h1ec == io_sel ? io_ins_492 : _GEN_491; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_493 = 10'h1ed == io_sel ? io_ins_493 : _GEN_492; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_494 = 10'h1ee == io_sel ? io_ins_494 : _GEN_493; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_495 = 10'h1ef == io_sel ? io_ins_495 : _GEN_494; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_496 = 10'h1f0 == io_sel ? io_ins_496 : _GEN_495; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_497 = 10'h1f1 == io_sel ? io_ins_497 : _GEN_496; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_498 = 10'h1f2 == io_sel ? io_ins_498 : _GEN_497; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_499 = 10'h1f3 == io_sel ? io_ins_499 : _GEN_498; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_500 = 10'h1f4 == io_sel ? io_ins_500 : _GEN_499; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_501 = 10'h1f5 == io_sel ? io_ins_501 : _GEN_500; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_502 = 10'h1f6 == io_sel ? io_ins_502 : _GEN_501; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_503 = 10'h1f7 == io_sel ? io_ins_503 : _GEN_502; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_504 = 10'h1f8 == io_sel ? io_ins_504 : _GEN_503; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_505 = 10'h1f9 == io_sel ? io_ins_505 : _GEN_504; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_506 = 10'h1fa == io_sel ? io_ins_506 : _GEN_505; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_507 = 10'h1fb == io_sel ? io_ins_507 : _GEN_506; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_508 = 10'h1fc == io_sel ? io_ins_508 : _GEN_507; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_509 = 10'h1fd == io_sel ? io_ins_509 : _GEN_508; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_510 = 10'h1fe == io_sel ? io_ins_510 : _GEN_509; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_511 = 10'h1ff == io_sel ? io_ins_511 : _GEN_510; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_512 = 10'h200 == io_sel ? io_ins_512 : _GEN_511; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_513 = 10'h201 == io_sel ? io_ins_513 : _GEN_512; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_514 = 10'h202 == io_sel ? io_ins_514 : _GEN_513; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_515 = 10'h203 == io_sel ? io_ins_515 : _GEN_514; // @[MuxN.scala 16:10:@47654.4]
  assign _GEN_516 = 10'h204 == io_sel ? io_ins_516 : _GEN_515; // @[MuxN.scala 16:10:@47654.4]
  assign io_out = 10'h205 == io_sel ? io_ins_517 : _GEN_516; // @[MuxN.scala 16:10:@47654.4]
endmodule
module RegFile( // @[:@47656.2]
  input         clock, // @[:@47657.4]
  input         reset, // @[:@47658.4]
  input  [31:0] io_raddr, // @[:@47659.4]
  input         io_wen, // @[:@47659.4]
  input  [31:0] io_waddr, // @[:@47659.4]
  input  [63:0] io_wdata, // @[:@47659.4]
  output [63:0] io_rdata, // @[:@47659.4]
  input         io_reset, // @[:@47659.4]
  output [63:0] io_argIns_0, // @[:@47659.4]
  output [63:0] io_argIns_1, // @[:@47659.4]
  output [63:0] io_argIns_2, // @[:@47659.4]
  input         io_argOuts_0_valid, // @[:@47659.4]
  input  [63:0] io_argOuts_0_bits, // @[:@47659.4]
  input         io_argOuts_1_valid, // @[:@47659.4]
  input  [63:0] io_argOuts_1_bits, // @[:@47659.4]
  input         io_argOuts_2_valid, // @[:@47659.4]
  input  [63:0] io_argOuts_2_bits, // @[:@47659.4]
  input         io_argOuts_3_valid, // @[:@47659.4]
  input  [63:0] io_argOuts_3_bits, // @[:@47659.4]
  input         io_argOuts_4_valid, // @[:@47659.4]
  input  [63:0] io_argOuts_4_bits, // @[:@47659.4]
  input         io_argOuts_5_valid, // @[:@47659.4]
  input  [63:0] io_argOuts_5_bits, // @[:@47659.4]
  input         io_argOuts_6_valid, // @[:@47659.4]
  input  [63:0] io_argOuts_6_bits, // @[:@47659.4]
  input         io_argOuts_7_valid, // @[:@47659.4]
  input  [63:0] io_argOuts_7_bits, // @[:@47659.4]
  input         io_argOuts_8_valid, // @[:@47659.4]
  input  [63:0] io_argOuts_8_bits, // @[:@47659.4]
  input         io_argOuts_9_valid, // @[:@47659.4]
  input  [63:0] io_argOuts_9_bits, // @[:@47659.4]
  input         io_argOuts_10_valid, // @[:@47659.4]
  input  [63:0] io_argOuts_10_bits, // @[:@47659.4]
  input         io_argOuts_11_valid, // @[:@47659.4]
  input  [63:0] io_argOuts_11_bits, // @[:@47659.4]
  input         io_argOuts_12_valid, // @[:@47659.4]
  input  [63:0] io_argOuts_12_bits, // @[:@47659.4]
  input         io_argOuts_13_valid, // @[:@47659.4]
  input  [63:0] io_argOuts_13_bits, // @[:@47659.4]
  input         io_argOuts_14_valid, // @[:@47659.4]
  input  [63:0] io_argOuts_14_bits, // @[:@47659.4]
  input         io_argOuts_15_valid, // @[:@47659.4]
  input  [63:0] io_argOuts_15_bits, // @[:@47659.4]
  input         io_argOuts_16_valid, // @[:@47659.4]
  input  [63:0] io_argOuts_16_bits, // @[:@47659.4]
  input  [63:0] io_argOuts_17_bits, // @[:@47659.4]
  input  [63:0] io_argOuts_18_bits, // @[:@47659.4]
  input  [63:0] io_argOuts_19_bits, // @[:@47659.4]
  input  [63:0] io_argOuts_20_bits, // @[:@47659.4]
  input  [63:0] io_argOuts_21_bits, // @[:@47659.4]
  input  [63:0] io_argOuts_22_bits, // @[:@47659.4]
  input  [63:0] io_argOuts_23_bits, // @[:@47659.4]
  input  [63:0] io_argOuts_24_bits, // @[:@47659.4]
  input  [63:0] io_argOuts_25_bits, // @[:@47659.4]
  input  [63:0] io_argOuts_26_bits, // @[:@47659.4]
  input  [63:0] io_argOuts_27_bits, // @[:@47659.4]
  input  [63:0] io_argOuts_28_bits, // @[:@47659.4]
  input  [63:0] io_argOuts_29_bits, // @[:@47659.4]
  input  [63:0] io_argOuts_30_bits, // @[:@47659.4]
  input  [63:0] io_argOuts_31_bits, // @[:@47659.4]
  input  [63:0] io_argOuts_32_bits, // @[:@47659.4]
  input  [63:0] io_argOuts_33_bits, // @[:@47659.4]
  input  [63:0] io_argOuts_34_bits, // @[:@47659.4]
  input  [63:0] io_argOuts_35_bits, // @[:@47659.4]
  input  [63:0] io_argOuts_36_bits, // @[:@47659.4]
  input  [63:0] io_argOuts_37_bits, // @[:@47659.4]
  input  [63:0] io_argOuts_38_bits, // @[:@47659.4]
  input  [63:0] io_argOuts_39_bits, // @[:@47659.4]
  input  [63:0] io_argOuts_40_bits, // @[:@47659.4]
  input  [63:0] io_argOuts_41_bits, // @[:@47659.4]
  input  [63:0] io_argOuts_42_bits, // @[:@47659.4]
  input  [63:0] io_argOuts_43_bits, // @[:@47659.4]
  input  [63:0] io_argOuts_44_bits, // @[:@47659.4]
  input  [63:0] io_argOuts_45_bits, // @[:@47659.4]
  input  [63:0] io_argOuts_46_bits, // @[:@47659.4]
  input  [63:0] io_argOuts_57_bits // @[:@47659.4]
);
  wire  regs_0_clock; // @[RegFile.scala 66:20:@49729.4]
  wire  regs_0_reset; // @[RegFile.scala 66:20:@49729.4]
  wire [63:0] regs_0_io_in; // @[RegFile.scala 66:20:@49729.4]
  wire  regs_0_io_reset; // @[RegFile.scala 66:20:@49729.4]
  wire [63:0] regs_0_io_out; // @[RegFile.scala 66:20:@49729.4]
  wire  regs_0_io_enable; // @[RegFile.scala 66:20:@49729.4]
  wire  regs_1_clock; // @[RegFile.scala 66:20:@49741.4]
  wire  regs_1_reset; // @[RegFile.scala 66:20:@49741.4]
  wire [63:0] regs_1_io_in; // @[RegFile.scala 66:20:@49741.4]
  wire  regs_1_io_reset; // @[RegFile.scala 66:20:@49741.4]
  wire [63:0] regs_1_io_out; // @[RegFile.scala 66:20:@49741.4]
  wire  regs_1_io_enable; // @[RegFile.scala 66:20:@49741.4]
  wire  regs_2_clock; // @[RegFile.scala 66:20:@49760.4]
  wire  regs_2_reset; // @[RegFile.scala 66:20:@49760.4]
  wire [63:0] regs_2_io_in; // @[RegFile.scala 66:20:@49760.4]
  wire  regs_2_io_reset; // @[RegFile.scala 66:20:@49760.4]
  wire [63:0] regs_2_io_out; // @[RegFile.scala 66:20:@49760.4]
  wire  regs_2_io_enable; // @[RegFile.scala 66:20:@49760.4]
  wire  regs_3_clock; // @[RegFile.scala 66:20:@49772.4]
  wire  regs_3_reset; // @[RegFile.scala 66:20:@49772.4]
  wire [63:0] regs_3_io_in; // @[RegFile.scala 66:20:@49772.4]
  wire  regs_3_io_reset; // @[RegFile.scala 66:20:@49772.4]
  wire [63:0] regs_3_io_out; // @[RegFile.scala 66:20:@49772.4]
  wire  regs_3_io_enable; // @[RegFile.scala 66:20:@49772.4]
  wire  regs_4_clock; // @[RegFile.scala 66:20:@49786.4]
  wire  regs_4_reset; // @[RegFile.scala 66:20:@49786.4]
  wire [63:0] regs_4_io_in; // @[RegFile.scala 66:20:@49786.4]
  wire  regs_4_io_reset; // @[RegFile.scala 66:20:@49786.4]
  wire [63:0] regs_4_io_out; // @[RegFile.scala 66:20:@49786.4]
  wire  regs_4_io_enable; // @[RegFile.scala 66:20:@49786.4]
  wire  regs_5_clock; // @[RegFile.scala 66:20:@49800.4]
  wire  regs_5_reset; // @[RegFile.scala 66:20:@49800.4]
  wire [63:0] regs_5_io_in; // @[RegFile.scala 66:20:@49800.4]
  wire  regs_5_io_reset; // @[RegFile.scala 66:20:@49800.4]
  wire [63:0] regs_5_io_out; // @[RegFile.scala 66:20:@49800.4]
  wire  regs_5_io_enable; // @[RegFile.scala 66:20:@49800.4]
  wire  regs_6_clock; // @[RegFile.scala 66:20:@49814.4]
  wire  regs_6_reset; // @[RegFile.scala 66:20:@49814.4]
  wire [63:0] regs_6_io_in; // @[RegFile.scala 66:20:@49814.4]
  wire  regs_6_io_reset; // @[RegFile.scala 66:20:@49814.4]
  wire [63:0] regs_6_io_out; // @[RegFile.scala 66:20:@49814.4]
  wire  regs_6_io_enable; // @[RegFile.scala 66:20:@49814.4]
  wire  regs_7_clock; // @[RegFile.scala 66:20:@49828.4]
  wire  regs_7_reset; // @[RegFile.scala 66:20:@49828.4]
  wire [63:0] regs_7_io_in; // @[RegFile.scala 66:20:@49828.4]
  wire  regs_7_io_reset; // @[RegFile.scala 66:20:@49828.4]
  wire [63:0] regs_7_io_out; // @[RegFile.scala 66:20:@49828.4]
  wire  regs_7_io_enable; // @[RegFile.scala 66:20:@49828.4]
  wire  regs_8_clock; // @[RegFile.scala 66:20:@49842.4]
  wire  regs_8_reset; // @[RegFile.scala 66:20:@49842.4]
  wire [63:0] regs_8_io_in; // @[RegFile.scala 66:20:@49842.4]
  wire  regs_8_io_reset; // @[RegFile.scala 66:20:@49842.4]
  wire [63:0] regs_8_io_out; // @[RegFile.scala 66:20:@49842.4]
  wire  regs_8_io_enable; // @[RegFile.scala 66:20:@49842.4]
  wire  regs_9_clock; // @[RegFile.scala 66:20:@49856.4]
  wire  regs_9_reset; // @[RegFile.scala 66:20:@49856.4]
  wire [63:0] regs_9_io_in; // @[RegFile.scala 66:20:@49856.4]
  wire  regs_9_io_reset; // @[RegFile.scala 66:20:@49856.4]
  wire [63:0] regs_9_io_out; // @[RegFile.scala 66:20:@49856.4]
  wire  regs_9_io_enable; // @[RegFile.scala 66:20:@49856.4]
  wire  regs_10_clock; // @[RegFile.scala 66:20:@49870.4]
  wire  regs_10_reset; // @[RegFile.scala 66:20:@49870.4]
  wire [63:0] regs_10_io_in; // @[RegFile.scala 66:20:@49870.4]
  wire  regs_10_io_reset; // @[RegFile.scala 66:20:@49870.4]
  wire [63:0] regs_10_io_out; // @[RegFile.scala 66:20:@49870.4]
  wire  regs_10_io_enable; // @[RegFile.scala 66:20:@49870.4]
  wire  regs_11_clock; // @[RegFile.scala 66:20:@49884.4]
  wire  regs_11_reset; // @[RegFile.scala 66:20:@49884.4]
  wire [63:0] regs_11_io_in; // @[RegFile.scala 66:20:@49884.4]
  wire  regs_11_io_reset; // @[RegFile.scala 66:20:@49884.4]
  wire [63:0] regs_11_io_out; // @[RegFile.scala 66:20:@49884.4]
  wire  regs_11_io_enable; // @[RegFile.scala 66:20:@49884.4]
  wire  regs_12_clock; // @[RegFile.scala 66:20:@49898.4]
  wire  regs_12_reset; // @[RegFile.scala 66:20:@49898.4]
  wire [63:0] regs_12_io_in; // @[RegFile.scala 66:20:@49898.4]
  wire  regs_12_io_reset; // @[RegFile.scala 66:20:@49898.4]
  wire [63:0] regs_12_io_out; // @[RegFile.scala 66:20:@49898.4]
  wire  regs_12_io_enable; // @[RegFile.scala 66:20:@49898.4]
  wire  regs_13_clock; // @[RegFile.scala 66:20:@49912.4]
  wire  regs_13_reset; // @[RegFile.scala 66:20:@49912.4]
  wire [63:0] regs_13_io_in; // @[RegFile.scala 66:20:@49912.4]
  wire  regs_13_io_reset; // @[RegFile.scala 66:20:@49912.4]
  wire [63:0] regs_13_io_out; // @[RegFile.scala 66:20:@49912.4]
  wire  regs_13_io_enable; // @[RegFile.scala 66:20:@49912.4]
  wire  regs_14_clock; // @[RegFile.scala 66:20:@49926.4]
  wire  regs_14_reset; // @[RegFile.scala 66:20:@49926.4]
  wire [63:0] regs_14_io_in; // @[RegFile.scala 66:20:@49926.4]
  wire  regs_14_io_reset; // @[RegFile.scala 66:20:@49926.4]
  wire [63:0] regs_14_io_out; // @[RegFile.scala 66:20:@49926.4]
  wire  regs_14_io_enable; // @[RegFile.scala 66:20:@49926.4]
  wire  regs_15_clock; // @[RegFile.scala 66:20:@49940.4]
  wire  regs_15_reset; // @[RegFile.scala 66:20:@49940.4]
  wire [63:0] regs_15_io_in; // @[RegFile.scala 66:20:@49940.4]
  wire  regs_15_io_reset; // @[RegFile.scala 66:20:@49940.4]
  wire [63:0] regs_15_io_out; // @[RegFile.scala 66:20:@49940.4]
  wire  regs_15_io_enable; // @[RegFile.scala 66:20:@49940.4]
  wire  regs_16_clock; // @[RegFile.scala 66:20:@49954.4]
  wire  regs_16_reset; // @[RegFile.scala 66:20:@49954.4]
  wire [63:0] regs_16_io_in; // @[RegFile.scala 66:20:@49954.4]
  wire  regs_16_io_reset; // @[RegFile.scala 66:20:@49954.4]
  wire [63:0] regs_16_io_out; // @[RegFile.scala 66:20:@49954.4]
  wire  regs_16_io_enable; // @[RegFile.scala 66:20:@49954.4]
  wire  regs_17_clock; // @[RegFile.scala 66:20:@49968.4]
  wire  regs_17_reset; // @[RegFile.scala 66:20:@49968.4]
  wire [63:0] regs_17_io_in; // @[RegFile.scala 66:20:@49968.4]
  wire  regs_17_io_reset; // @[RegFile.scala 66:20:@49968.4]
  wire [63:0] regs_17_io_out; // @[RegFile.scala 66:20:@49968.4]
  wire  regs_17_io_enable; // @[RegFile.scala 66:20:@49968.4]
  wire  regs_18_clock; // @[RegFile.scala 66:20:@49982.4]
  wire  regs_18_reset; // @[RegFile.scala 66:20:@49982.4]
  wire [63:0] regs_18_io_in; // @[RegFile.scala 66:20:@49982.4]
  wire  regs_18_io_reset; // @[RegFile.scala 66:20:@49982.4]
  wire [63:0] regs_18_io_out; // @[RegFile.scala 66:20:@49982.4]
  wire  regs_18_io_enable; // @[RegFile.scala 66:20:@49982.4]
  wire  regs_19_clock; // @[RegFile.scala 66:20:@49996.4]
  wire  regs_19_reset; // @[RegFile.scala 66:20:@49996.4]
  wire [63:0] regs_19_io_in; // @[RegFile.scala 66:20:@49996.4]
  wire  regs_19_io_reset; // @[RegFile.scala 66:20:@49996.4]
  wire [63:0] regs_19_io_out; // @[RegFile.scala 66:20:@49996.4]
  wire  regs_19_io_enable; // @[RegFile.scala 66:20:@49996.4]
  wire  regs_20_clock; // @[RegFile.scala 66:20:@50010.4]
  wire  regs_20_reset; // @[RegFile.scala 66:20:@50010.4]
  wire [63:0] regs_20_io_in; // @[RegFile.scala 66:20:@50010.4]
  wire  regs_20_io_reset; // @[RegFile.scala 66:20:@50010.4]
  wire [63:0] regs_20_io_out; // @[RegFile.scala 66:20:@50010.4]
  wire  regs_20_io_enable; // @[RegFile.scala 66:20:@50010.4]
  wire  regs_21_clock; // @[RegFile.scala 66:20:@50024.4]
  wire  regs_21_reset; // @[RegFile.scala 66:20:@50024.4]
  wire [63:0] regs_21_io_in; // @[RegFile.scala 66:20:@50024.4]
  wire  regs_21_io_reset; // @[RegFile.scala 66:20:@50024.4]
  wire [63:0] regs_21_io_out; // @[RegFile.scala 66:20:@50024.4]
  wire  regs_21_io_enable; // @[RegFile.scala 66:20:@50024.4]
  wire  regs_22_clock; // @[RegFile.scala 66:20:@50038.4]
  wire  regs_22_reset; // @[RegFile.scala 66:20:@50038.4]
  wire [63:0] regs_22_io_in; // @[RegFile.scala 66:20:@50038.4]
  wire  regs_22_io_reset; // @[RegFile.scala 66:20:@50038.4]
  wire [63:0] regs_22_io_out; // @[RegFile.scala 66:20:@50038.4]
  wire  regs_22_io_enable; // @[RegFile.scala 66:20:@50038.4]
  wire  regs_23_clock; // @[RegFile.scala 66:20:@50052.4]
  wire  regs_23_reset; // @[RegFile.scala 66:20:@50052.4]
  wire [63:0] regs_23_io_in; // @[RegFile.scala 66:20:@50052.4]
  wire  regs_23_io_reset; // @[RegFile.scala 66:20:@50052.4]
  wire [63:0] regs_23_io_out; // @[RegFile.scala 66:20:@50052.4]
  wire  regs_23_io_enable; // @[RegFile.scala 66:20:@50052.4]
  wire  regs_24_clock; // @[RegFile.scala 66:20:@50066.4]
  wire  regs_24_reset; // @[RegFile.scala 66:20:@50066.4]
  wire [63:0] regs_24_io_in; // @[RegFile.scala 66:20:@50066.4]
  wire  regs_24_io_reset; // @[RegFile.scala 66:20:@50066.4]
  wire [63:0] regs_24_io_out; // @[RegFile.scala 66:20:@50066.4]
  wire  regs_24_io_enable; // @[RegFile.scala 66:20:@50066.4]
  wire  regs_25_clock; // @[RegFile.scala 66:20:@50080.4]
  wire  regs_25_reset; // @[RegFile.scala 66:20:@50080.4]
  wire [63:0] regs_25_io_in; // @[RegFile.scala 66:20:@50080.4]
  wire  regs_25_io_reset; // @[RegFile.scala 66:20:@50080.4]
  wire [63:0] regs_25_io_out; // @[RegFile.scala 66:20:@50080.4]
  wire  regs_25_io_enable; // @[RegFile.scala 66:20:@50080.4]
  wire  regs_26_clock; // @[RegFile.scala 66:20:@50094.4]
  wire  regs_26_reset; // @[RegFile.scala 66:20:@50094.4]
  wire [63:0] regs_26_io_in; // @[RegFile.scala 66:20:@50094.4]
  wire  regs_26_io_reset; // @[RegFile.scala 66:20:@50094.4]
  wire [63:0] regs_26_io_out; // @[RegFile.scala 66:20:@50094.4]
  wire  regs_26_io_enable; // @[RegFile.scala 66:20:@50094.4]
  wire  regs_27_clock; // @[RegFile.scala 66:20:@50108.4]
  wire  regs_27_reset; // @[RegFile.scala 66:20:@50108.4]
  wire [63:0] regs_27_io_in; // @[RegFile.scala 66:20:@50108.4]
  wire  regs_27_io_reset; // @[RegFile.scala 66:20:@50108.4]
  wire [63:0] regs_27_io_out; // @[RegFile.scala 66:20:@50108.4]
  wire  regs_27_io_enable; // @[RegFile.scala 66:20:@50108.4]
  wire  regs_28_clock; // @[RegFile.scala 66:20:@50122.4]
  wire  regs_28_reset; // @[RegFile.scala 66:20:@50122.4]
  wire [63:0] regs_28_io_in; // @[RegFile.scala 66:20:@50122.4]
  wire  regs_28_io_reset; // @[RegFile.scala 66:20:@50122.4]
  wire [63:0] regs_28_io_out; // @[RegFile.scala 66:20:@50122.4]
  wire  regs_28_io_enable; // @[RegFile.scala 66:20:@50122.4]
  wire  regs_29_clock; // @[RegFile.scala 66:20:@50136.4]
  wire  regs_29_reset; // @[RegFile.scala 66:20:@50136.4]
  wire [63:0] regs_29_io_in; // @[RegFile.scala 66:20:@50136.4]
  wire  regs_29_io_reset; // @[RegFile.scala 66:20:@50136.4]
  wire [63:0] regs_29_io_out; // @[RegFile.scala 66:20:@50136.4]
  wire  regs_29_io_enable; // @[RegFile.scala 66:20:@50136.4]
  wire  regs_30_clock; // @[RegFile.scala 66:20:@50150.4]
  wire  regs_30_reset; // @[RegFile.scala 66:20:@50150.4]
  wire [63:0] regs_30_io_in; // @[RegFile.scala 66:20:@50150.4]
  wire  regs_30_io_reset; // @[RegFile.scala 66:20:@50150.4]
  wire [63:0] regs_30_io_out; // @[RegFile.scala 66:20:@50150.4]
  wire  regs_30_io_enable; // @[RegFile.scala 66:20:@50150.4]
  wire  regs_31_clock; // @[RegFile.scala 66:20:@50164.4]
  wire  regs_31_reset; // @[RegFile.scala 66:20:@50164.4]
  wire [63:0] regs_31_io_in; // @[RegFile.scala 66:20:@50164.4]
  wire  regs_31_io_reset; // @[RegFile.scala 66:20:@50164.4]
  wire [63:0] regs_31_io_out; // @[RegFile.scala 66:20:@50164.4]
  wire  regs_31_io_enable; // @[RegFile.scala 66:20:@50164.4]
  wire  regs_32_clock; // @[RegFile.scala 66:20:@50178.4]
  wire  regs_32_reset; // @[RegFile.scala 66:20:@50178.4]
  wire [63:0] regs_32_io_in; // @[RegFile.scala 66:20:@50178.4]
  wire  regs_32_io_reset; // @[RegFile.scala 66:20:@50178.4]
  wire [63:0] regs_32_io_out; // @[RegFile.scala 66:20:@50178.4]
  wire  regs_32_io_enable; // @[RegFile.scala 66:20:@50178.4]
  wire  regs_33_clock; // @[RegFile.scala 66:20:@50192.4]
  wire  regs_33_reset; // @[RegFile.scala 66:20:@50192.4]
  wire [63:0] regs_33_io_in; // @[RegFile.scala 66:20:@50192.4]
  wire  regs_33_io_reset; // @[RegFile.scala 66:20:@50192.4]
  wire [63:0] regs_33_io_out; // @[RegFile.scala 66:20:@50192.4]
  wire  regs_33_io_enable; // @[RegFile.scala 66:20:@50192.4]
  wire  regs_34_clock; // @[RegFile.scala 66:20:@50206.4]
  wire  regs_34_reset; // @[RegFile.scala 66:20:@50206.4]
  wire [63:0] regs_34_io_in; // @[RegFile.scala 66:20:@50206.4]
  wire  regs_34_io_reset; // @[RegFile.scala 66:20:@50206.4]
  wire [63:0] regs_34_io_out; // @[RegFile.scala 66:20:@50206.4]
  wire  regs_34_io_enable; // @[RegFile.scala 66:20:@50206.4]
  wire  regs_35_clock; // @[RegFile.scala 66:20:@50220.4]
  wire  regs_35_reset; // @[RegFile.scala 66:20:@50220.4]
  wire [63:0] regs_35_io_in; // @[RegFile.scala 66:20:@50220.4]
  wire  regs_35_io_reset; // @[RegFile.scala 66:20:@50220.4]
  wire [63:0] regs_35_io_out; // @[RegFile.scala 66:20:@50220.4]
  wire  regs_35_io_enable; // @[RegFile.scala 66:20:@50220.4]
  wire  regs_36_clock; // @[RegFile.scala 66:20:@50234.4]
  wire  regs_36_reset; // @[RegFile.scala 66:20:@50234.4]
  wire [63:0] regs_36_io_in; // @[RegFile.scala 66:20:@50234.4]
  wire  regs_36_io_reset; // @[RegFile.scala 66:20:@50234.4]
  wire [63:0] regs_36_io_out; // @[RegFile.scala 66:20:@50234.4]
  wire  regs_36_io_enable; // @[RegFile.scala 66:20:@50234.4]
  wire  regs_37_clock; // @[RegFile.scala 66:20:@50248.4]
  wire  regs_37_reset; // @[RegFile.scala 66:20:@50248.4]
  wire [63:0] regs_37_io_in; // @[RegFile.scala 66:20:@50248.4]
  wire  regs_37_io_reset; // @[RegFile.scala 66:20:@50248.4]
  wire [63:0] regs_37_io_out; // @[RegFile.scala 66:20:@50248.4]
  wire  regs_37_io_enable; // @[RegFile.scala 66:20:@50248.4]
  wire  regs_38_clock; // @[RegFile.scala 66:20:@50262.4]
  wire  regs_38_reset; // @[RegFile.scala 66:20:@50262.4]
  wire [63:0] regs_38_io_in; // @[RegFile.scala 66:20:@50262.4]
  wire  regs_38_io_reset; // @[RegFile.scala 66:20:@50262.4]
  wire [63:0] regs_38_io_out; // @[RegFile.scala 66:20:@50262.4]
  wire  regs_38_io_enable; // @[RegFile.scala 66:20:@50262.4]
  wire  regs_39_clock; // @[RegFile.scala 66:20:@50276.4]
  wire  regs_39_reset; // @[RegFile.scala 66:20:@50276.4]
  wire [63:0] regs_39_io_in; // @[RegFile.scala 66:20:@50276.4]
  wire  regs_39_io_reset; // @[RegFile.scala 66:20:@50276.4]
  wire [63:0] regs_39_io_out; // @[RegFile.scala 66:20:@50276.4]
  wire  regs_39_io_enable; // @[RegFile.scala 66:20:@50276.4]
  wire  regs_40_clock; // @[RegFile.scala 66:20:@50290.4]
  wire  regs_40_reset; // @[RegFile.scala 66:20:@50290.4]
  wire [63:0] regs_40_io_in; // @[RegFile.scala 66:20:@50290.4]
  wire  regs_40_io_reset; // @[RegFile.scala 66:20:@50290.4]
  wire [63:0] regs_40_io_out; // @[RegFile.scala 66:20:@50290.4]
  wire  regs_40_io_enable; // @[RegFile.scala 66:20:@50290.4]
  wire  regs_41_clock; // @[RegFile.scala 66:20:@50304.4]
  wire  regs_41_reset; // @[RegFile.scala 66:20:@50304.4]
  wire [63:0] regs_41_io_in; // @[RegFile.scala 66:20:@50304.4]
  wire  regs_41_io_reset; // @[RegFile.scala 66:20:@50304.4]
  wire [63:0] regs_41_io_out; // @[RegFile.scala 66:20:@50304.4]
  wire  regs_41_io_enable; // @[RegFile.scala 66:20:@50304.4]
  wire  regs_42_clock; // @[RegFile.scala 66:20:@50318.4]
  wire  regs_42_reset; // @[RegFile.scala 66:20:@50318.4]
  wire [63:0] regs_42_io_in; // @[RegFile.scala 66:20:@50318.4]
  wire  regs_42_io_reset; // @[RegFile.scala 66:20:@50318.4]
  wire [63:0] regs_42_io_out; // @[RegFile.scala 66:20:@50318.4]
  wire  regs_42_io_enable; // @[RegFile.scala 66:20:@50318.4]
  wire  regs_43_clock; // @[RegFile.scala 66:20:@50332.4]
  wire  regs_43_reset; // @[RegFile.scala 66:20:@50332.4]
  wire [63:0] regs_43_io_in; // @[RegFile.scala 66:20:@50332.4]
  wire  regs_43_io_reset; // @[RegFile.scala 66:20:@50332.4]
  wire [63:0] regs_43_io_out; // @[RegFile.scala 66:20:@50332.4]
  wire  regs_43_io_enable; // @[RegFile.scala 66:20:@50332.4]
  wire  regs_44_clock; // @[RegFile.scala 66:20:@50346.4]
  wire  regs_44_reset; // @[RegFile.scala 66:20:@50346.4]
  wire [63:0] regs_44_io_in; // @[RegFile.scala 66:20:@50346.4]
  wire  regs_44_io_reset; // @[RegFile.scala 66:20:@50346.4]
  wire [63:0] regs_44_io_out; // @[RegFile.scala 66:20:@50346.4]
  wire  regs_44_io_enable; // @[RegFile.scala 66:20:@50346.4]
  wire  regs_45_clock; // @[RegFile.scala 66:20:@50360.4]
  wire  regs_45_reset; // @[RegFile.scala 66:20:@50360.4]
  wire [63:0] regs_45_io_in; // @[RegFile.scala 66:20:@50360.4]
  wire  regs_45_io_reset; // @[RegFile.scala 66:20:@50360.4]
  wire [63:0] regs_45_io_out; // @[RegFile.scala 66:20:@50360.4]
  wire  regs_45_io_enable; // @[RegFile.scala 66:20:@50360.4]
  wire  regs_46_clock; // @[RegFile.scala 66:20:@50374.4]
  wire  regs_46_reset; // @[RegFile.scala 66:20:@50374.4]
  wire [63:0] regs_46_io_in; // @[RegFile.scala 66:20:@50374.4]
  wire  regs_46_io_reset; // @[RegFile.scala 66:20:@50374.4]
  wire [63:0] regs_46_io_out; // @[RegFile.scala 66:20:@50374.4]
  wire  regs_46_io_enable; // @[RegFile.scala 66:20:@50374.4]
  wire  regs_47_clock; // @[RegFile.scala 66:20:@50388.4]
  wire  regs_47_reset; // @[RegFile.scala 66:20:@50388.4]
  wire [63:0] regs_47_io_in; // @[RegFile.scala 66:20:@50388.4]
  wire  regs_47_io_reset; // @[RegFile.scala 66:20:@50388.4]
  wire [63:0] regs_47_io_out; // @[RegFile.scala 66:20:@50388.4]
  wire  regs_47_io_enable; // @[RegFile.scala 66:20:@50388.4]
  wire  regs_48_clock; // @[RegFile.scala 66:20:@50402.4]
  wire  regs_48_reset; // @[RegFile.scala 66:20:@50402.4]
  wire [63:0] regs_48_io_in; // @[RegFile.scala 66:20:@50402.4]
  wire  regs_48_io_reset; // @[RegFile.scala 66:20:@50402.4]
  wire [63:0] regs_48_io_out; // @[RegFile.scala 66:20:@50402.4]
  wire  regs_48_io_enable; // @[RegFile.scala 66:20:@50402.4]
  wire  regs_49_clock; // @[RegFile.scala 66:20:@50416.4]
  wire  regs_49_reset; // @[RegFile.scala 66:20:@50416.4]
  wire [63:0] regs_49_io_in; // @[RegFile.scala 66:20:@50416.4]
  wire  regs_49_io_reset; // @[RegFile.scala 66:20:@50416.4]
  wire [63:0] regs_49_io_out; // @[RegFile.scala 66:20:@50416.4]
  wire  regs_49_io_enable; // @[RegFile.scala 66:20:@50416.4]
  wire  regs_50_clock; // @[RegFile.scala 66:20:@50430.4]
  wire  regs_50_reset; // @[RegFile.scala 66:20:@50430.4]
  wire [63:0] regs_50_io_in; // @[RegFile.scala 66:20:@50430.4]
  wire  regs_50_io_reset; // @[RegFile.scala 66:20:@50430.4]
  wire [63:0] regs_50_io_out; // @[RegFile.scala 66:20:@50430.4]
  wire  regs_50_io_enable; // @[RegFile.scala 66:20:@50430.4]
  wire  regs_51_clock; // @[RegFile.scala 66:20:@50444.4]
  wire  regs_51_reset; // @[RegFile.scala 66:20:@50444.4]
  wire [63:0] regs_51_io_in; // @[RegFile.scala 66:20:@50444.4]
  wire  regs_51_io_reset; // @[RegFile.scala 66:20:@50444.4]
  wire [63:0] regs_51_io_out; // @[RegFile.scala 66:20:@50444.4]
  wire  regs_51_io_enable; // @[RegFile.scala 66:20:@50444.4]
  wire  regs_52_clock; // @[RegFile.scala 66:20:@50458.4]
  wire  regs_52_reset; // @[RegFile.scala 66:20:@50458.4]
  wire [63:0] regs_52_io_in; // @[RegFile.scala 66:20:@50458.4]
  wire  regs_52_io_reset; // @[RegFile.scala 66:20:@50458.4]
  wire [63:0] regs_52_io_out; // @[RegFile.scala 66:20:@50458.4]
  wire  regs_52_io_enable; // @[RegFile.scala 66:20:@50458.4]
  wire  regs_53_clock; // @[RegFile.scala 66:20:@50472.4]
  wire  regs_53_reset; // @[RegFile.scala 66:20:@50472.4]
  wire [63:0] regs_53_io_in; // @[RegFile.scala 66:20:@50472.4]
  wire  regs_53_io_reset; // @[RegFile.scala 66:20:@50472.4]
  wire [63:0] regs_53_io_out; // @[RegFile.scala 66:20:@50472.4]
  wire  regs_53_io_enable; // @[RegFile.scala 66:20:@50472.4]
  wire  regs_54_clock; // @[RegFile.scala 66:20:@50486.4]
  wire  regs_54_reset; // @[RegFile.scala 66:20:@50486.4]
  wire [63:0] regs_54_io_in; // @[RegFile.scala 66:20:@50486.4]
  wire  regs_54_io_reset; // @[RegFile.scala 66:20:@50486.4]
  wire [63:0] regs_54_io_out; // @[RegFile.scala 66:20:@50486.4]
  wire  regs_54_io_enable; // @[RegFile.scala 66:20:@50486.4]
  wire  regs_55_clock; // @[RegFile.scala 66:20:@50500.4]
  wire  regs_55_reset; // @[RegFile.scala 66:20:@50500.4]
  wire [63:0] regs_55_io_in; // @[RegFile.scala 66:20:@50500.4]
  wire  regs_55_io_reset; // @[RegFile.scala 66:20:@50500.4]
  wire [63:0] regs_55_io_out; // @[RegFile.scala 66:20:@50500.4]
  wire  regs_55_io_enable; // @[RegFile.scala 66:20:@50500.4]
  wire  regs_56_clock; // @[RegFile.scala 66:20:@50514.4]
  wire  regs_56_reset; // @[RegFile.scala 66:20:@50514.4]
  wire [63:0] regs_56_io_in; // @[RegFile.scala 66:20:@50514.4]
  wire  regs_56_io_reset; // @[RegFile.scala 66:20:@50514.4]
  wire [63:0] regs_56_io_out; // @[RegFile.scala 66:20:@50514.4]
  wire  regs_56_io_enable; // @[RegFile.scala 66:20:@50514.4]
  wire  regs_57_clock; // @[RegFile.scala 66:20:@50528.4]
  wire  regs_57_reset; // @[RegFile.scala 66:20:@50528.4]
  wire [63:0] regs_57_io_in; // @[RegFile.scala 66:20:@50528.4]
  wire  regs_57_io_reset; // @[RegFile.scala 66:20:@50528.4]
  wire [63:0] regs_57_io_out; // @[RegFile.scala 66:20:@50528.4]
  wire  regs_57_io_enable; // @[RegFile.scala 66:20:@50528.4]
  wire  regs_58_clock; // @[RegFile.scala 66:20:@50542.4]
  wire  regs_58_reset; // @[RegFile.scala 66:20:@50542.4]
  wire [63:0] regs_58_io_in; // @[RegFile.scala 66:20:@50542.4]
  wire  regs_58_io_reset; // @[RegFile.scala 66:20:@50542.4]
  wire [63:0] regs_58_io_out; // @[RegFile.scala 66:20:@50542.4]
  wire  regs_58_io_enable; // @[RegFile.scala 66:20:@50542.4]
  wire  regs_59_clock; // @[RegFile.scala 66:20:@50556.4]
  wire  regs_59_reset; // @[RegFile.scala 66:20:@50556.4]
  wire [63:0] regs_59_io_in; // @[RegFile.scala 66:20:@50556.4]
  wire  regs_59_io_reset; // @[RegFile.scala 66:20:@50556.4]
  wire [63:0] regs_59_io_out; // @[RegFile.scala 66:20:@50556.4]
  wire  regs_59_io_enable; // @[RegFile.scala 66:20:@50556.4]
  wire  regs_60_clock; // @[RegFile.scala 66:20:@50570.4]
  wire  regs_60_reset; // @[RegFile.scala 66:20:@50570.4]
  wire [63:0] regs_60_io_in; // @[RegFile.scala 66:20:@50570.4]
  wire  regs_60_io_reset; // @[RegFile.scala 66:20:@50570.4]
  wire [63:0] regs_60_io_out; // @[RegFile.scala 66:20:@50570.4]
  wire  regs_60_io_enable; // @[RegFile.scala 66:20:@50570.4]
  wire  regs_61_clock; // @[RegFile.scala 66:20:@50584.4]
  wire  regs_61_reset; // @[RegFile.scala 66:20:@50584.4]
  wire [63:0] regs_61_io_in; // @[RegFile.scala 66:20:@50584.4]
  wire  regs_61_io_reset; // @[RegFile.scala 66:20:@50584.4]
  wire [63:0] regs_61_io_out; // @[RegFile.scala 66:20:@50584.4]
  wire  regs_61_io_enable; // @[RegFile.scala 66:20:@50584.4]
  wire  regs_62_clock; // @[RegFile.scala 66:20:@50598.4]
  wire  regs_62_reset; // @[RegFile.scala 66:20:@50598.4]
  wire [63:0] regs_62_io_in; // @[RegFile.scala 66:20:@50598.4]
  wire  regs_62_io_reset; // @[RegFile.scala 66:20:@50598.4]
  wire [63:0] regs_62_io_out; // @[RegFile.scala 66:20:@50598.4]
  wire  regs_62_io_enable; // @[RegFile.scala 66:20:@50598.4]
  wire  regs_63_clock; // @[RegFile.scala 66:20:@50612.4]
  wire  regs_63_reset; // @[RegFile.scala 66:20:@50612.4]
  wire [63:0] regs_63_io_in; // @[RegFile.scala 66:20:@50612.4]
  wire  regs_63_io_reset; // @[RegFile.scala 66:20:@50612.4]
  wire [63:0] regs_63_io_out; // @[RegFile.scala 66:20:@50612.4]
  wire  regs_63_io_enable; // @[RegFile.scala 66:20:@50612.4]
  wire  regs_64_clock; // @[RegFile.scala 66:20:@50626.4]
  wire  regs_64_reset; // @[RegFile.scala 66:20:@50626.4]
  wire [63:0] regs_64_io_in; // @[RegFile.scala 66:20:@50626.4]
  wire  regs_64_io_reset; // @[RegFile.scala 66:20:@50626.4]
  wire [63:0] regs_64_io_out; // @[RegFile.scala 66:20:@50626.4]
  wire  regs_64_io_enable; // @[RegFile.scala 66:20:@50626.4]
  wire  regs_65_clock; // @[RegFile.scala 66:20:@50640.4]
  wire  regs_65_reset; // @[RegFile.scala 66:20:@50640.4]
  wire [63:0] regs_65_io_in; // @[RegFile.scala 66:20:@50640.4]
  wire  regs_65_io_reset; // @[RegFile.scala 66:20:@50640.4]
  wire [63:0] regs_65_io_out; // @[RegFile.scala 66:20:@50640.4]
  wire  regs_65_io_enable; // @[RegFile.scala 66:20:@50640.4]
  wire  regs_66_clock; // @[RegFile.scala 66:20:@50654.4]
  wire  regs_66_reset; // @[RegFile.scala 66:20:@50654.4]
  wire [63:0] regs_66_io_in; // @[RegFile.scala 66:20:@50654.4]
  wire  regs_66_io_reset; // @[RegFile.scala 66:20:@50654.4]
  wire [63:0] regs_66_io_out; // @[RegFile.scala 66:20:@50654.4]
  wire  regs_66_io_enable; // @[RegFile.scala 66:20:@50654.4]
  wire  regs_67_clock; // @[RegFile.scala 66:20:@50668.4]
  wire  regs_67_reset; // @[RegFile.scala 66:20:@50668.4]
  wire [63:0] regs_67_io_in; // @[RegFile.scala 66:20:@50668.4]
  wire  regs_67_io_reset; // @[RegFile.scala 66:20:@50668.4]
  wire [63:0] regs_67_io_out; // @[RegFile.scala 66:20:@50668.4]
  wire  regs_67_io_enable; // @[RegFile.scala 66:20:@50668.4]
  wire  regs_68_clock; // @[RegFile.scala 66:20:@50682.4]
  wire  regs_68_reset; // @[RegFile.scala 66:20:@50682.4]
  wire [63:0] regs_68_io_in; // @[RegFile.scala 66:20:@50682.4]
  wire  regs_68_io_reset; // @[RegFile.scala 66:20:@50682.4]
  wire [63:0] regs_68_io_out; // @[RegFile.scala 66:20:@50682.4]
  wire  regs_68_io_enable; // @[RegFile.scala 66:20:@50682.4]
  wire  regs_69_clock; // @[RegFile.scala 66:20:@50696.4]
  wire  regs_69_reset; // @[RegFile.scala 66:20:@50696.4]
  wire [63:0] regs_69_io_in; // @[RegFile.scala 66:20:@50696.4]
  wire  regs_69_io_reset; // @[RegFile.scala 66:20:@50696.4]
  wire [63:0] regs_69_io_out; // @[RegFile.scala 66:20:@50696.4]
  wire  regs_69_io_enable; // @[RegFile.scala 66:20:@50696.4]
  wire  regs_70_clock; // @[RegFile.scala 66:20:@50710.4]
  wire  regs_70_reset; // @[RegFile.scala 66:20:@50710.4]
  wire [63:0] regs_70_io_in; // @[RegFile.scala 66:20:@50710.4]
  wire  regs_70_io_reset; // @[RegFile.scala 66:20:@50710.4]
  wire [63:0] regs_70_io_out; // @[RegFile.scala 66:20:@50710.4]
  wire  regs_70_io_enable; // @[RegFile.scala 66:20:@50710.4]
  wire  regs_71_clock; // @[RegFile.scala 66:20:@50724.4]
  wire  regs_71_reset; // @[RegFile.scala 66:20:@50724.4]
  wire [63:0] regs_71_io_in; // @[RegFile.scala 66:20:@50724.4]
  wire  regs_71_io_reset; // @[RegFile.scala 66:20:@50724.4]
  wire [63:0] regs_71_io_out; // @[RegFile.scala 66:20:@50724.4]
  wire  regs_71_io_enable; // @[RegFile.scala 66:20:@50724.4]
  wire  regs_72_clock; // @[RegFile.scala 66:20:@50738.4]
  wire  regs_72_reset; // @[RegFile.scala 66:20:@50738.4]
  wire [63:0] regs_72_io_in; // @[RegFile.scala 66:20:@50738.4]
  wire  regs_72_io_reset; // @[RegFile.scala 66:20:@50738.4]
  wire [63:0] regs_72_io_out; // @[RegFile.scala 66:20:@50738.4]
  wire  regs_72_io_enable; // @[RegFile.scala 66:20:@50738.4]
  wire  regs_73_clock; // @[RegFile.scala 66:20:@50752.4]
  wire  regs_73_reset; // @[RegFile.scala 66:20:@50752.4]
  wire [63:0] regs_73_io_in; // @[RegFile.scala 66:20:@50752.4]
  wire  regs_73_io_reset; // @[RegFile.scala 66:20:@50752.4]
  wire [63:0] regs_73_io_out; // @[RegFile.scala 66:20:@50752.4]
  wire  regs_73_io_enable; // @[RegFile.scala 66:20:@50752.4]
  wire  regs_74_clock; // @[RegFile.scala 66:20:@50766.4]
  wire  regs_74_reset; // @[RegFile.scala 66:20:@50766.4]
  wire [63:0] regs_74_io_in; // @[RegFile.scala 66:20:@50766.4]
  wire  regs_74_io_reset; // @[RegFile.scala 66:20:@50766.4]
  wire [63:0] regs_74_io_out; // @[RegFile.scala 66:20:@50766.4]
  wire  regs_74_io_enable; // @[RegFile.scala 66:20:@50766.4]
  wire  regs_75_clock; // @[RegFile.scala 66:20:@50780.4]
  wire  regs_75_reset; // @[RegFile.scala 66:20:@50780.4]
  wire [63:0] regs_75_io_in; // @[RegFile.scala 66:20:@50780.4]
  wire  regs_75_io_reset; // @[RegFile.scala 66:20:@50780.4]
  wire [63:0] regs_75_io_out; // @[RegFile.scala 66:20:@50780.4]
  wire  regs_75_io_enable; // @[RegFile.scala 66:20:@50780.4]
  wire  regs_76_clock; // @[RegFile.scala 66:20:@50794.4]
  wire  regs_76_reset; // @[RegFile.scala 66:20:@50794.4]
  wire [63:0] regs_76_io_in; // @[RegFile.scala 66:20:@50794.4]
  wire  regs_76_io_reset; // @[RegFile.scala 66:20:@50794.4]
  wire [63:0] regs_76_io_out; // @[RegFile.scala 66:20:@50794.4]
  wire  regs_76_io_enable; // @[RegFile.scala 66:20:@50794.4]
  wire  regs_77_clock; // @[RegFile.scala 66:20:@50808.4]
  wire  regs_77_reset; // @[RegFile.scala 66:20:@50808.4]
  wire [63:0] regs_77_io_in; // @[RegFile.scala 66:20:@50808.4]
  wire  regs_77_io_reset; // @[RegFile.scala 66:20:@50808.4]
  wire [63:0] regs_77_io_out; // @[RegFile.scala 66:20:@50808.4]
  wire  regs_77_io_enable; // @[RegFile.scala 66:20:@50808.4]
  wire  regs_78_clock; // @[RegFile.scala 66:20:@50822.4]
  wire  regs_78_reset; // @[RegFile.scala 66:20:@50822.4]
  wire [63:0] regs_78_io_in; // @[RegFile.scala 66:20:@50822.4]
  wire  regs_78_io_reset; // @[RegFile.scala 66:20:@50822.4]
  wire [63:0] regs_78_io_out; // @[RegFile.scala 66:20:@50822.4]
  wire  regs_78_io_enable; // @[RegFile.scala 66:20:@50822.4]
  wire  regs_79_clock; // @[RegFile.scala 66:20:@50836.4]
  wire  regs_79_reset; // @[RegFile.scala 66:20:@50836.4]
  wire [63:0] regs_79_io_in; // @[RegFile.scala 66:20:@50836.4]
  wire  regs_79_io_reset; // @[RegFile.scala 66:20:@50836.4]
  wire [63:0] regs_79_io_out; // @[RegFile.scala 66:20:@50836.4]
  wire  regs_79_io_enable; // @[RegFile.scala 66:20:@50836.4]
  wire  regs_80_clock; // @[RegFile.scala 66:20:@50850.4]
  wire  regs_80_reset; // @[RegFile.scala 66:20:@50850.4]
  wire [63:0] regs_80_io_in; // @[RegFile.scala 66:20:@50850.4]
  wire  regs_80_io_reset; // @[RegFile.scala 66:20:@50850.4]
  wire [63:0] regs_80_io_out; // @[RegFile.scala 66:20:@50850.4]
  wire  regs_80_io_enable; // @[RegFile.scala 66:20:@50850.4]
  wire  regs_81_clock; // @[RegFile.scala 66:20:@50864.4]
  wire  regs_81_reset; // @[RegFile.scala 66:20:@50864.4]
  wire [63:0] regs_81_io_in; // @[RegFile.scala 66:20:@50864.4]
  wire  regs_81_io_reset; // @[RegFile.scala 66:20:@50864.4]
  wire [63:0] regs_81_io_out; // @[RegFile.scala 66:20:@50864.4]
  wire  regs_81_io_enable; // @[RegFile.scala 66:20:@50864.4]
  wire  regs_82_clock; // @[RegFile.scala 66:20:@50878.4]
  wire  regs_82_reset; // @[RegFile.scala 66:20:@50878.4]
  wire [63:0] regs_82_io_in; // @[RegFile.scala 66:20:@50878.4]
  wire  regs_82_io_reset; // @[RegFile.scala 66:20:@50878.4]
  wire [63:0] regs_82_io_out; // @[RegFile.scala 66:20:@50878.4]
  wire  regs_82_io_enable; // @[RegFile.scala 66:20:@50878.4]
  wire  regs_83_clock; // @[RegFile.scala 66:20:@50892.4]
  wire  regs_83_reset; // @[RegFile.scala 66:20:@50892.4]
  wire [63:0] regs_83_io_in; // @[RegFile.scala 66:20:@50892.4]
  wire  regs_83_io_reset; // @[RegFile.scala 66:20:@50892.4]
  wire [63:0] regs_83_io_out; // @[RegFile.scala 66:20:@50892.4]
  wire  regs_83_io_enable; // @[RegFile.scala 66:20:@50892.4]
  wire  regs_84_clock; // @[RegFile.scala 66:20:@50906.4]
  wire  regs_84_reset; // @[RegFile.scala 66:20:@50906.4]
  wire [63:0] regs_84_io_in; // @[RegFile.scala 66:20:@50906.4]
  wire  regs_84_io_reset; // @[RegFile.scala 66:20:@50906.4]
  wire [63:0] regs_84_io_out; // @[RegFile.scala 66:20:@50906.4]
  wire  regs_84_io_enable; // @[RegFile.scala 66:20:@50906.4]
  wire  regs_85_clock; // @[RegFile.scala 66:20:@50920.4]
  wire  regs_85_reset; // @[RegFile.scala 66:20:@50920.4]
  wire [63:0] regs_85_io_in; // @[RegFile.scala 66:20:@50920.4]
  wire  regs_85_io_reset; // @[RegFile.scala 66:20:@50920.4]
  wire [63:0] regs_85_io_out; // @[RegFile.scala 66:20:@50920.4]
  wire  regs_85_io_enable; // @[RegFile.scala 66:20:@50920.4]
  wire  regs_86_clock; // @[RegFile.scala 66:20:@50934.4]
  wire  regs_86_reset; // @[RegFile.scala 66:20:@50934.4]
  wire [63:0] regs_86_io_in; // @[RegFile.scala 66:20:@50934.4]
  wire  regs_86_io_reset; // @[RegFile.scala 66:20:@50934.4]
  wire [63:0] regs_86_io_out; // @[RegFile.scala 66:20:@50934.4]
  wire  regs_86_io_enable; // @[RegFile.scala 66:20:@50934.4]
  wire  regs_87_clock; // @[RegFile.scala 66:20:@50948.4]
  wire  regs_87_reset; // @[RegFile.scala 66:20:@50948.4]
  wire [63:0] regs_87_io_in; // @[RegFile.scala 66:20:@50948.4]
  wire  regs_87_io_reset; // @[RegFile.scala 66:20:@50948.4]
  wire [63:0] regs_87_io_out; // @[RegFile.scala 66:20:@50948.4]
  wire  regs_87_io_enable; // @[RegFile.scala 66:20:@50948.4]
  wire  regs_88_clock; // @[RegFile.scala 66:20:@50962.4]
  wire  regs_88_reset; // @[RegFile.scala 66:20:@50962.4]
  wire [63:0] regs_88_io_in; // @[RegFile.scala 66:20:@50962.4]
  wire  regs_88_io_reset; // @[RegFile.scala 66:20:@50962.4]
  wire [63:0] regs_88_io_out; // @[RegFile.scala 66:20:@50962.4]
  wire  regs_88_io_enable; // @[RegFile.scala 66:20:@50962.4]
  wire  regs_89_clock; // @[RegFile.scala 66:20:@50976.4]
  wire  regs_89_reset; // @[RegFile.scala 66:20:@50976.4]
  wire [63:0] regs_89_io_in; // @[RegFile.scala 66:20:@50976.4]
  wire  regs_89_io_reset; // @[RegFile.scala 66:20:@50976.4]
  wire [63:0] regs_89_io_out; // @[RegFile.scala 66:20:@50976.4]
  wire  regs_89_io_enable; // @[RegFile.scala 66:20:@50976.4]
  wire  regs_90_clock; // @[RegFile.scala 66:20:@50990.4]
  wire  regs_90_reset; // @[RegFile.scala 66:20:@50990.4]
  wire [63:0] regs_90_io_in; // @[RegFile.scala 66:20:@50990.4]
  wire  regs_90_io_reset; // @[RegFile.scala 66:20:@50990.4]
  wire [63:0] regs_90_io_out; // @[RegFile.scala 66:20:@50990.4]
  wire  regs_90_io_enable; // @[RegFile.scala 66:20:@50990.4]
  wire  regs_91_clock; // @[RegFile.scala 66:20:@51004.4]
  wire  regs_91_reset; // @[RegFile.scala 66:20:@51004.4]
  wire [63:0] regs_91_io_in; // @[RegFile.scala 66:20:@51004.4]
  wire  regs_91_io_reset; // @[RegFile.scala 66:20:@51004.4]
  wire [63:0] regs_91_io_out; // @[RegFile.scala 66:20:@51004.4]
  wire  regs_91_io_enable; // @[RegFile.scala 66:20:@51004.4]
  wire  regs_92_clock; // @[RegFile.scala 66:20:@51018.4]
  wire  regs_92_reset; // @[RegFile.scala 66:20:@51018.4]
  wire [63:0] regs_92_io_in; // @[RegFile.scala 66:20:@51018.4]
  wire  regs_92_io_reset; // @[RegFile.scala 66:20:@51018.4]
  wire [63:0] regs_92_io_out; // @[RegFile.scala 66:20:@51018.4]
  wire  regs_92_io_enable; // @[RegFile.scala 66:20:@51018.4]
  wire  regs_93_clock; // @[RegFile.scala 66:20:@51032.4]
  wire  regs_93_reset; // @[RegFile.scala 66:20:@51032.4]
  wire [63:0] regs_93_io_in; // @[RegFile.scala 66:20:@51032.4]
  wire  regs_93_io_reset; // @[RegFile.scala 66:20:@51032.4]
  wire [63:0] regs_93_io_out; // @[RegFile.scala 66:20:@51032.4]
  wire  regs_93_io_enable; // @[RegFile.scala 66:20:@51032.4]
  wire  regs_94_clock; // @[RegFile.scala 66:20:@51046.4]
  wire  regs_94_reset; // @[RegFile.scala 66:20:@51046.4]
  wire [63:0] regs_94_io_in; // @[RegFile.scala 66:20:@51046.4]
  wire  regs_94_io_reset; // @[RegFile.scala 66:20:@51046.4]
  wire [63:0] regs_94_io_out; // @[RegFile.scala 66:20:@51046.4]
  wire  regs_94_io_enable; // @[RegFile.scala 66:20:@51046.4]
  wire  regs_95_clock; // @[RegFile.scala 66:20:@51060.4]
  wire  regs_95_reset; // @[RegFile.scala 66:20:@51060.4]
  wire [63:0] regs_95_io_in; // @[RegFile.scala 66:20:@51060.4]
  wire  regs_95_io_reset; // @[RegFile.scala 66:20:@51060.4]
  wire [63:0] regs_95_io_out; // @[RegFile.scala 66:20:@51060.4]
  wire  regs_95_io_enable; // @[RegFile.scala 66:20:@51060.4]
  wire  regs_96_clock; // @[RegFile.scala 66:20:@51074.4]
  wire  regs_96_reset; // @[RegFile.scala 66:20:@51074.4]
  wire [63:0] regs_96_io_in; // @[RegFile.scala 66:20:@51074.4]
  wire  regs_96_io_reset; // @[RegFile.scala 66:20:@51074.4]
  wire [63:0] regs_96_io_out; // @[RegFile.scala 66:20:@51074.4]
  wire  regs_96_io_enable; // @[RegFile.scala 66:20:@51074.4]
  wire  regs_97_clock; // @[RegFile.scala 66:20:@51088.4]
  wire  regs_97_reset; // @[RegFile.scala 66:20:@51088.4]
  wire [63:0] regs_97_io_in; // @[RegFile.scala 66:20:@51088.4]
  wire  regs_97_io_reset; // @[RegFile.scala 66:20:@51088.4]
  wire [63:0] regs_97_io_out; // @[RegFile.scala 66:20:@51088.4]
  wire  regs_97_io_enable; // @[RegFile.scala 66:20:@51088.4]
  wire  regs_98_clock; // @[RegFile.scala 66:20:@51102.4]
  wire  regs_98_reset; // @[RegFile.scala 66:20:@51102.4]
  wire [63:0] regs_98_io_in; // @[RegFile.scala 66:20:@51102.4]
  wire  regs_98_io_reset; // @[RegFile.scala 66:20:@51102.4]
  wire [63:0] regs_98_io_out; // @[RegFile.scala 66:20:@51102.4]
  wire  regs_98_io_enable; // @[RegFile.scala 66:20:@51102.4]
  wire  regs_99_clock; // @[RegFile.scala 66:20:@51116.4]
  wire  regs_99_reset; // @[RegFile.scala 66:20:@51116.4]
  wire [63:0] regs_99_io_in; // @[RegFile.scala 66:20:@51116.4]
  wire  regs_99_io_reset; // @[RegFile.scala 66:20:@51116.4]
  wire [63:0] regs_99_io_out; // @[RegFile.scala 66:20:@51116.4]
  wire  regs_99_io_enable; // @[RegFile.scala 66:20:@51116.4]
  wire  regs_100_clock; // @[RegFile.scala 66:20:@51130.4]
  wire  regs_100_reset; // @[RegFile.scala 66:20:@51130.4]
  wire [63:0] regs_100_io_in; // @[RegFile.scala 66:20:@51130.4]
  wire  regs_100_io_reset; // @[RegFile.scala 66:20:@51130.4]
  wire [63:0] regs_100_io_out; // @[RegFile.scala 66:20:@51130.4]
  wire  regs_100_io_enable; // @[RegFile.scala 66:20:@51130.4]
  wire  regs_101_clock; // @[RegFile.scala 66:20:@51144.4]
  wire  regs_101_reset; // @[RegFile.scala 66:20:@51144.4]
  wire [63:0] regs_101_io_in; // @[RegFile.scala 66:20:@51144.4]
  wire  regs_101_io_reset; // @[RegFile.scala 66:20:@51144.4]
  wire [63:0] regs_101_io_out; // @[RegFile.scala 66:20:@51144.4]
  wire  regs_101_io_enable; // @[RegFile.scala 66:20:@51144.4]
  wire  regs_102_clock; // @[RegFile.scala 66:20:@51158.4]
  wire  regs_102_reset; // @[RegFile.scala 66:20:@51158.4]
  wire [63:0] regs_102_io_in; // @[RegFile.scala 66:20:@51158.4]
  wire  regs_102_io_reset; // @[RegFile.scala 66:20:@51158.4]
  wire [63:0] regs_102_io_out; // @[RegFile.scala 66:20:@51158.4]
  wire  regs_102_io_enable; // @[RegFile.scala 66:20:@51158.4]
  wire  regs_103_clock; // @[RegFile.scala 66:20:@51172.4]
  wire  regs_103_reset; // @[RegFile.scala 66:20:@51172.4]
  wire [63:0] regs_103_io_in; // @[RegFile.scala 66:20:@51172.4]
  wire  regs_103_io_reset; // @[RegFile.scala 66:20:@51172.4]
  wire [63:0] regs_103_io_out; // @[RegFile.scala 66:20:@51172.4]
  wire  regs_103_io_enable; // @[RegFile.scala 66:20:@51172.4]
  wire  regs_104_clock; // @[RegFile.scala 66:20:@51186.4]
  wire  regs_104_reset; // @[RegFile.scala 66:20:@51186.4]
  wire [63:0] regs_104_io_in; // @[RegFile.scala 66:20:@51186.4]
  wire  regs_104_io_reset; // @[RegFile.scala 66:20:@51186.4]
  wire [63:0] regs_104_io_out; // @[RegFile.scala 66:20:@51186.4]
  wire  regs_104_io_enable; // @[RegFile.scala 66:20:@51186.4]
  wire  regs_105_clock; // @[RegFile.scala 66:20:@51200.4]
  wire  regs_105_reset; // @[RegFile.scala 66:20:@51200.4]
  wire [63:0] regs_105_io_in; // @[RegFile.scala 66:20:@51200.4]
  wire  regs_105_io_reset; // @[RegFile.scala 66:20:@51200.4]
  wire [63:0] regs_105_io_out; // @[RegFile.scala 66:20:@51200.4]
  wire  regs_105_io_enable; // @[RegFile.scala 66:20:@51200.4]
  wire  regs_106_clock; // @[RegFile.scala 66:20:@51214.4]
  wire  regs_106_reset; // @[RegFile.scala 66:20:@51214.4]
  wire [63:0] regs_106_io_in; // @[RegFile.scala 66:20:@51214.4]
  wire  regs_106_io_reset; // @[RegFile.scala 66:20:@51214.4]
  wire [63:0] regs_106_io_out; // @[RegFile.scala 66:20:@51214.4]
  wire  regs_106_io_enable; // @[RegFile.scala 66:20:@51214.4]
  wire  regs_107_clock; // @[RegFile.scala 66:20:@51228.4]
  wire  regs_107_reset; // @[RegFile.scala 66:20:@51228.4]
  wire [63:0] regs_107_io_in; // @[RegFile.scala 66:20:@51228.4]
  wire  regs_107_io_reset; // @[RegFile.scala 66:20:@51228.4]
  wire [63:0] regs_107_io_out; // @[RegFile.scala 66:20:@51228.4]
  wire  regs_107_io_enable; // @[RegFile.scala 66:20:@51228.4]
  wire  regs_108_clock; // @[RegFile.scala 66:20:@51242.4]
  wire  regs_108_reset; // @[RegFile.scala 66:20:@51242.4]
  wire [63:0] regs_108_io_in; // @[RegFile.scala 66:20:@51242.4]
  wire  regs_108_io_reset; // @[RegFile.scala 66:20:@51242.4]
  wire [63:0] regs_108_io_out; // @[RegFile.scala 66:20:@51242.4]
  wire  regs_108_io_enable; // @[RegFile.scala 66:20:@51242.4]
  wire  regs_109_clock; // @[RegFile.scala 66:20:@51256.4]
  wire  regs_109_reset; // @[RegFile.scala 66:20:@51256.4]
  wire [63:0] regs_109_io_in; // @[RegFile.scala 66:20:@51256.4]
  wire  regs_109_io_reset; // @[RegFile.scala 66:20:@51256.4]
  wire [63:0] regs_109_io_out; // @[RegFile.scala 66:20:@51256.4]
  wire  regs_109_io_enable; // @[RegFile.scala 66:20:@51256.4]
  wire  regs_110_clock; // @[RegFile.scala 66:20:@51270.4]
  wire  regs_110_reset; // @[RegFile.scala 66:20:@51270.4]
  wire [63:0] regs_110_io_in; // @[RegFile.scala 66:20:@51270.4]
  wire  regs_110_io_reset; // @[RegFile.scala 66:20:@51270.4]
  wire [63:0] regs_110_io_out; // @[RegFile.scala 66:20:@51270.4]
  wire  regs_110_io_enable; // @[RegFile.scala 66:20:@51270.4]
  wire  regs_111_clock; // @[RegFile.scala 66:20:@51284.4]
  wire  regs_111_reset; // @[RegFile.scala 66:20:@51284.4]
  wire [63:0] regs_111_io_in; // @[RegFile.scala 66:20:@51284.4]
  wire  regs_111_io_reset; // @[RegFile.scala 66:20:@51284.4]
  wire [63:0] regs_111_io_out; // @[RegFile.scala 66:20:@51284.4]
  wire  regs_111_io_enable; // @[RegFile.scala 66:20:@51284.4]
  wire  regs_112_clock; // @[RegFile.scala 66:20:@51298.4]
  wire  regs_112_reset; // @[RegFile.scala 66:20:@51298.4]
  wire [63:0] regs_112_io_in; // @[RegFile.scala 66:20:@51298.4]
  wire  regs_112_io_reset; // @[RegFile.scala 66:20:@51298.4]
  wire [63:0] regs_112_io_out; // @[RegFile.scala 66:20:@51298.4]
  wire  regs_112_io_enable; // @[RegFile.scala 66:20:@51298.4]
  wire  regs_113_clock; // @[RegFile.scala 66:20:@51312.4]
  wire  regs_113_reset; // @[RegFile.scala 66:20:@51312.4]
  wire [63:0] regs_113_io_in; // @[RegFile.scala 66:20:@51312.4]
  wire  regs_113_io_reset; // @[RegFile.scala 66:20:@51312.4]
  wire [63:0] regs_113_io_out; // @[RegFile.scala 66:20:@51312.4]
  wire  regs_113_io_enable; // @[RegFile.scala 66:20:@51312.4]
  wire  regs_114_clock; // @[RegFile.scala 66:20:@51326.4]
  wire  regs_114_reset; // @[RegFile.scala 66:20:@51326.4]
  wire [63:0] regs_114_io_in; // @[RegFile.scala 66:20:@51326.4]
  wire  regs_114_io_reset; // @[RegFile.scala 66:20:@51326.4]
  wire [63:0] regs_114_io_out; // @[RegFile.scala 66:20:@51326.4]
  wire  regs_114_io_enable; // @[RegFile.scala 66:20:@51326.4]
  wire  regs_115_clock; // @[RegFile.scala 66:20:@51340.4]
  wire  regs_115_reset; // @[RegFile.scala 66:20:@51340.4]
  wire [63:0] regs_115_io_in; // @[RegFile.scala 66:20:@51340.4]
  wire  regs_115_io_reset; // @[RegFile.scala 66:20:@51340.4]
  wire [63:0] regs_115_io_out; // @[RegFile.scala 66:20:@51340.4]
  wire  regs_115_io_enable; // @[RegFile.scala 66:20:@51340.4]
  wire  regs_116_clock; // @[RegFile.scala 66:20:@51354.4]
  wire  regs_116_reset; // @[RegFile.scala 66:20:@51354.4]
  wire [63:0] regs_116_io_in; // @[RegFile.scala 66:20:@51354.4]
  wire  regs_116_io_reset; // @[RegFile.scala 66:20:@51354.4]
  wire [63:0] regs_116_io_out; // @[RegFile.scala 66:20:@51354.4]
  wire  regs_116_io_enable; // @[RegFile.scala 66:20:@51354.4]
  wire  regs_117_clock; // @[RegFile.scala 66:20:@51368.4]
  wire  regs_117_reset; // @[RegFile.scala 66:20:@51368.4]
  wire [63:0] regs_117_io_in; // @[RegFile.scala 66:20:@51368.4]
  wire  regs_117_io_reset; // @[RegFile.scala 66:20:@51368.4]
  wire [63:0] regs_117_io_out; // @[RegFile.scala 66:20:@51368.4]
  wire  regs_117_io_enable; // @[RegFile.scala 66:20:@51368.4]
  wire  regs_118_clock; // @[RegFile.scala 66:20:@51382.4]
  wire  regs_118_reset; // @[RegFile.scala 66:20:@51382.4]
  wire [63:0] regs_118_io_in; // @[RegFile.scala 66:20:@51382.4]
  wire  regs_118_io_reset; // @[RegFile.scala 66:20:@51382.4]
  wire [63:0] regs_118_io_out; // @[RegFile.scala 66:20:@51382.4]
  wire  regs_118_io_enable; // @[RegFile.scala 66:20:@51382.4]
  wire  regs_119_clock; // @[RegFile.scala 66:20:@51396.4]
  wire  regs_119_reset; // @[RegFile.scala 66:20:@51396.4]
  wire [63:0] regs_119_io_in; // @[RegFile.scala 66:20:@51396.4]
  wire  regs_119_io_reset; // @[RegFile.scala 66:20:@51396.4]
  wire [63:0] regs_119_io_out; // @[RegFile.scala 66:20:@51396.4]
  wire  regs_119_io_enable; // @[RegFile.scala 66:20:@51396.4]
  wire  regs_120_clock; // @[RegFile.scala 66:20:@51410.4]
  wire  regs_120_reset; // @[RegFile.scala 66:20:@51410.4]
  wire [63:0] regs_120_io_in; // @[RegFile.scala 66:20:@51410.4]
  wire  regs_120_io_reset; // @[RegFile.scala 66:20:@51410.4]
  wire [63:0] regs_120_io_out; // @[RegFile.scala 66:20:@51410.4]
  wire  regs_120_io_enable; // @[RegFile.scala 66:20:@51410.4]
  wire  regs_121_clock; // @[RegFile.scala 66:20:@51424.4]
  wire  regs_121_reset; // @[RegFile.scala 66:20:@51424.4]
  wire [63:0] regs_121_io_in; // @[RegFile.scala 66:20:@51424.4]
  wire  regs_121_io_reset; // @[RegFile.scala 66:20:@51424.4]
  wire [63:0] regs_121_io_out; // @[RegFile.scala 66:20:@51424.4]
  wire  regs_121_io_enable; // @[RegFile.scala 66:20:@51424.4]
  wire  regs_122_clock; // @[RegFile.scala 66:20:@51438.4]
  wire  regs_122_reset; // @[RegFile.scala 66:20:@51438.4]
  wire [63:0] regs_122_io_in; // @[RegFile.scala 66:20:@51438.4]
  wire  regs_122_io_reset; // @[RegFile.scala 66:20:@51438.4]
  wire [63:0] regs_122_io_out; // @[RegFile.scala 66:20:@51438.4]
  wire  regs_122_io_enable; // @[RegFile.scala 66:20:@51438.4]
  wire  regs_123_clock; // @[RegFile.scala 66:20:@51452.4]
  wire  regs_123_reset; // @[RegFile.scala 66:20:@51452.4]
  wire [63:0] regs_123_io_in; // @[RegFile.scala 66:20:@51452.4]
  wire  regs_123_io_reset; // @[RegFile.scala 66:20:@51452.4]
  wire [63:0] regs_123_io_out; // @[RegFile.scala 66:20:@51452.4]
  wire  regs_123_io_enable; // @[RegFile.scala 66:20:@51452.4]
  wire  regs_124_clock; // @[RegFile.scala 66:20:@51466.4]
  wire  regs_124_reset; // @[RegFile.scala 66:20:@51466.4]
  wire [63:0] regs_124_io_in; // @[RegFile.scala 66:20:@51466.4]
  wire  regs_124_io_reset; // @[RegFile.scala 66:20:@51466.4]
  wire [63:0] regs_124_io_out; // @[RegFile.scala 66:20:@51466.4]
  wire  regs_124_io_enable; // @[RegFile.scala 66:20:@51466.4]
  wire  regs_125_clock; // @[RegFile.scala 66:20:@51480.4]
  wire  regs_125_reset; // @[RegFile.scala 66:20:@51480.4]
  wire [63:0] regs_125_io_in; // @[RegFile.scala 66:20:@51480.4]
  wire  regs_125_io_reset; // @[RegFile.scala 66:20:@51480.4]
  wire [63:0] regs_125_io_out; // @[RegFile.scala 66:20:@51480.4]
  wire  regs_125_io_enable; // @[RegFile.scala 66:20:@51480.4]
  wire  regs_126_clock; // @[RegFile.scala 66:20:@51494.4]
  wire  regs_126_reset; // @[RegFile.scala 66:20:@51494.4]
  wire [63:0] regs_126_io_in; // @[RegFile.scala 66:20:@51494.4]
  wire  regs_126_io_reset; // @[RegFile.scala 66:20:@51494.4]
  wire [63:0] regs_126_io_out; // @[RegFile.scala 66:20:@51494.4]
  wire  regs_126_io_enable; // @[RegFile.scala 66:20:@51494.4]
  wire  regs_127_clock; // @[RegFile.scala 66:20:@51508.4]
  wire  regs_127_reset; // @[RegFile.scala 66:20:@51508.4]
  wire [63:0] regs_127_io_in; // @[RegFile.scala 66:20:@51508.4]
  wire  regs_127_io_reset; // @[RegFile.scala 66:20:@51508.4]
  wire [63:0] regs_127_io_out; // @[RegFile.scala 66:20:@51508.4]
  wire  regs_127_io_enable; // @[RegFile.scala 66:20:@51508.4]
  wire  regs_128_clock; // @[RegFile.scala 66:20:@51522.4]
  wire  regs_128_reset; // @[RegFile.scala 66:20:@51522.4]
  wire [63:0] regs_128_io_in; // @[RegFile.scala 66:20:@51522.4]
  wire  regs_128_io_reset; // @[RegFile.scala 66:20:@51522.4]
  wire [63:0] regs_128_io_out; // @[RegFile.scala 66:20:@51522.4]
  wire  regs_128_io_enable; // @[RegFile.scala 66:20:@51522.4]
  wire  regs_129_clock; // @[RegFile.scala 66:20:@51536.4]
  wire  regs_129_reset; // @[RegFile.scala 66:20:@51536.4]
  wire [63:0] regs_129_io_in; // @[RegFile.scala 66:20:@51536.4]
  wire  regs_129_io_reset; // @[RegFile.scala 66:20:@51536.4]
  wire [63:0] regs_129_io_out; // @[RegFile.scala 66:20:@51536.4]
  wire  regs_129_io_enable; // @[RegFile.scala 66:20:@51536.4]
  wire  regs_130_clock; // @[RegFile.scala 66:20:@51550.4]
  wire  regs_130_reset; // @[RegFile.scala 66:20:@51550.4]
  wire [63:0] regs_130_io_in; // @[RegFile.scala 66:20:@51550.4]
  wire  regs_130_io_reset; // @[RegFile.scala 66:20:@51550.4]
  wire [63:0] regs_130_io_out; // @[RegFile.scala 66:20:@51550.4]
  wire  regs_130_io_enable; // @[RegFile.scala 66:20:@51550.4]
  wire  regs_131_clock; // @[RegFile.scala 66:20:@51564.4]
  wire  regs_131_reset; // @[RegFile.scala 66:20:@51564.4]
  wire [63:0] regs_131_io_in; // @[RegFile.scala 66:20:@51564.4]
  wire  regs_131_io_reset; // @[RegFile.scala 66:20:@51564.4]
  wire [63:0] regs_131_io_out; // @[RegFile.scala 66:20:@51564.4]
  wire  regs_131_io_enable; // @[RegFile.scala 66:20:@51564.4]
  wire  regs_132_clock; // @[RegFile.scala 66:20:@51578.4]
  wire  regs_132_reset; // @[RegFile.scala 66:20:@51578.4]
  wire [63:0] regs_132_io_in; // @[RegFile.scala 66:20:@51578.4]
  wire  regs_132_io_reset; // @[RegFile.scala 66:20:@51578.4]
  wire [63:0] regs_132_io_out; // @[RegFile.scala 66:20:@51578.4]
  wire  regs_132_io_enable; // @[RegFile.scala 66:20:@51578.4]
  wire  regs_133_clock; // @[RegFile.scala 66:20:@51592.4]
  wire  regs_133_reset; // @[RegFile.scala 66:20:@51592.4]
  wire [63:0] regs_133_io_in; // @[RegFile.scala 66:20:@51592.4]
  wire  regs_133_io_reset; // @[RegFile.scala 66:20:@51592.4]
  wire [63:0] regs_133_io_out; // @[RegFile.scala 66:20:@51592.4]
  wire  regs_133_io_enable; // @[RegFile.scala 66:20:@51592.4]
  wire  regs_134_clock; // @[RegFile.scala 66:20:@51606.4]
  wire  regs_134_reset; // @[RegFile.scala 66:20:@51606.4]
  wire [63:0] regs_134_io_in; // @[RegFile.scala 66:20:@51606.4]
  wire  regs_134_io_reset; // @[RegFile.scala 66:20:@51606.4]
  wire [63:0] regs_134_io_out; // @[RegFile.scala 66:20:@51606.4]
  wire  regs_134_io_enable; // @[RegFile.scala 66:20:@51606.4]
  wire  regs_135_clock; // @[RegFile.scala 66:20:@51620.4]
  wire  regs_135_reset; // @[RegFile.scala 66:20:@51620.4]
  wire [63:0] regs_135_io_in; // @[RegFile.scala 66:20:@51620.4]
  wire  regs_135_io_reset; // @[RegFile.scala 66:20:@51620.4]
  wire [63:0] regs_135_io_out; // @[RegFile.scala 66:20:@51620.4]
  wire  regs_135_io_enable; // @[RegFile.scala 66:20:@51620.4]
  wire  regs_136_clock; // @[RegFile.scala 66:20:@51634.4]
  wire  regs_136_reset; // @[RegFile.scala 66:20:@51634.4]
  wire [63:0] regs_136_io_in; // @[RegFile.scala 66:20:@51634.4]
  wire  regs_136_io_reset; // @[RegFile.scala 66:20:@51634.4]
  wire [63:0] regs_136_io_out; // @[RegFile.scala 66:20:@51634.4]
  wire  regs_136_io_enable; // @[RegFile.scala 66:20:@51634.4]
  wire  regs_137_clock; // @[RegFile.scala 66:20:@51648.4]
  wire  regs_137_reset; // @[RegFile.scala 66:20:@51648.4]
  wire [63:0] regs_137_io_in; // @[RegFile.scala 66:20:@51648.4]
  wire  regs_137_io_reset; // @[RegFile.scala 66:20:@51648.4]
  wire [63:0] regs_137_io_out; // @[RegFile.scala 66:20:@51648.4]
  wire  regs_137_io_enable; // @[RegFile.scala 66:20:@51648.4]
  wire  regs_138_clock; // @[RegFile.scala 66:20:@51662.4]
  wire  regs_138_reset; // @[RegFile.scala 66:20:@51662.4]
  wire [63:0] regs_138_io_in; // @[RegFile.scala 66:20:@51662.4]
  wire  regs_138_io_reset; // @[RegFile.scala 66:20:@51662.4]
  wire [63:0] regs_138_io_out; // @[RegFile.scala 66:20:@51662.4]
  wire  regs_138_io_enable; // @[RegFile.scala 66:20:@51662.4]
  wire  regs_139_clock; // @[RegFile.scala 66:20:@51676.4]
  wire  regs_139_reset; // @[RegFile.scala 66:20:@51676.4]
  wire [63:0] regs_139_io_in; // @[RegFile.scala 66:20:@51676.4]
  wire  regs_139_io_reset; // @[RegFile.scala 66:20:@51676.4]
  wire [63:0] regs_139_io_out; // @[RegFile.scala 66:20:@51676.4]
  wire  regs_139_io_enable; // @[RegFile.scala 66:20:@51676.4]
  wire  regs_140_clock; // @[RegFile.scala 66:20:@51690.4]
  wire  regs_140_reset; // @[RegFile.scala 66:20:@51690.4]
  wire [63:0] regs_140_io_in; // @[RegFile.scala 66:20:@51690.4]
  wire  regs_140_io_reset; // @[RegFile.scala 66:20:@51690.4]
  wire [63:0] regs_140_io_out; // @[RegFile.scala 66:20:@51690.4]
  wire  regs_140_io_enable; // @[RegFile.scala 66:20:@51690.4]
  wire  regs_141_clock; // @[RegFile.scala 66:20:@51704.4]
  wire  regs_141_reset; // @[RegFile.scala 66:20:@51704.4]
  wire [63:0] regs_141_io_in; // @[RegFile.scala 66:20:@51704.4]
  wire  regs_141_io_reset; // @[RegFile.scala 66:20:@51704.4]
  wire [63:0] regs_141_io_out; // @[RegFile.scala 66:20:@51704.4]
  wire  regs_141_io_enable; // @[RegFile.scala 66:20:@51704.4]
  wire  regs_142_clock; // @[RegFile.scala 66:20:@51718.4]
  wire  regs_142_reset; // @[RegFile.scala 66:20:@51718.4]
  wire [63:0] regs_142_io_in; // @[RegFile.scala 66:20:@51718.4]
  wire  regs_142_io_reset; // @[RegFile.scala 66:20:@51718.4]
  wire [63:0] regs_142_io_out; // @[RegFile.scala 66:20:@51718.4]
  wire  regs_142_io_enable; // @[RegFile.scala 66:20:@51718.4]
  wire  regs_143_clock; // @[RegFile.scala 66:20:@51732.4]
  wire  regs_143_reset; // @[RegFile.scala 66:20:@51732.4]
  wire [63:0] regs_143_io_in; // @[RegFile.scala 66:20:@51732.4]
  wire  regs_143_io_reset; // @[RegFile.scala 66:20:@51732.4]
  wire [63:0] regs_143_io_out; // @[RegFile.scala 66:20:@51732.4]
  wire  regs_143_io_enable; // @[RegFile.scala 66:20:@51732.4]
  wire  regs_144_clock; // @[RegFile.scala 66:20:@51746.4]
  wire  regs_144_reset; // @[RegFile.scala 66:20:@51746.4]
  wire [63:0] regs_144_io_in; // @[RegFile.scala 66:20:@51746.4]
  wire  regs_144_io_reset; // @[RegFile.scala 66:20:@51746.4]
  wire [63:0] regs_144_io_out; // @[RegFile.scala 66:20:@51746.4]
  wire  regs_144_io_enable; // @[RegFile.scala 66:20:@51746.4]
  wire  regs_145_clock; // @[RegFile.scala 66:20:@51760.4]
  wire  regs_145_reset; // @[RegFile.scala 66:20:@51760.4]
  wire [63:0] regs_145_io_in; // @[RegFile.scala 66:20:@51760.4]
  wire  regs_145_io_reset; // @[RegFile.scala 66:20:@51760.4]
  wire [63:0] regs_145_io_out; // @[RegFile.scala 66:20:@51760.4]
  wire  regs_145_io_enable; // @[RegFile.scala 66:20:@51760.4]
  wire  regs_146_clock; // @[RegFile.scala 66:20:@51774.4]
  wire  regs_146_reset; // @[RegFile.scala 66:20:@51774.4]
  wire [63:0] regs_146_io_in; // @[RegFile.scala 66:20:@51774.4]
  wire  regs_146_io_reset; // @[RegFile.scala 66:20:@51774.4]
  wire [63:0] regs_146_io_out; // @[RegFile.scala 66:20:@51774.4]
  wire  regs_146_io_enable; // @[RegFile.scala 66:20:@51774.4]
  wire  regs_147_clock; // @[RegFile.scala 66:20:@51788.4]
  wire  regs_147_reset; // @[RegFile.scala 66:20:@51788.4]
  wire [63:0] regs_147_io_in; // @[RegFile.scala 66:20:@51788.4]
  wire  regs_147_io_reset; // @[RegFile.scala 66:20:@51788.4]
  wire [63:0] regs_147_io_out; // @[RegFile.scala 66:20:@51788.4]
  wire  regs_147_io_enable; // @[RegFile.scala 66:20:@51788.4]
  wire  regs_148_clock; // @[RegFile.scala 66:20:@51802.4]
  wire  regs_148_reset; // @[RegFile.scala 66:20:@51802.4]
  wire [63:0] regs_148_io_in; // @[RegFile.scala 66:20:@51802.4]
  wire  regs_148_io_reset; // @[RegFile.scala 66:20:@51802.4]
  wire [63:0] regs_148_io_out; // @[RegFile.scala 66:20:@51802.4]
  wire  regs_148_io_enable; // @[RegFile.scala 66:20:@51802.4]
  wire  regs_149_clock; // @[RegFile.scala 66:20:@51816.4]
  wire  regs_149_reset; // @[RegFile.scala 66:20:@51816.4]
  wire [63:0] regs_149_io_in; // @[RegFile.scala 66:20:@51816.4]
  wire  regs_149_io_reset; // @[RegFile.scala 66:20:@51816.4]
  wire [63:0] regs_149_io_out; // @[RegFile.scala 66:20:@51816.4]
  wire  regs_149_io_enable; // @[RegFile.scala 66:20:@51816.4]
  wire  regs_150_clock; // @[RegFile.scala 66:20:@51830.4]
  wire  regs_150_reset; // @[RegFile.scala 66:20:@51830.4]
  wire [63:0] regs_150_io_in; // @[RegFile.scala 66:20:@51830.4]
  wire  regs_150_io_reset; // @[RegFile.scala 66:20:@51830.4]
  wire [63:0] regs_150_io_out; // @[RegFile.scala 66:20:@51830.4]
  wire  regs_150_io_enable; // @[RegFile.scala 66:20:@51830.4]
  wire  regs_151_clock; // @[RegFile.scala 66:20:@51844.4]
  wire  regs_151_reset; // @[RegFile.scala 66:20:@51844.4]
  wire [63:0] regs_151_io_in; // @[RegFile.scala 66:20:@51844.4]
  wire  regs_151_io_reset; // @[RegFile.scala 66:20:@51844.4]
  wire [63:0] regs_151_io_out; // @[RegFile.scala 66:20:@51844.4]
  wire  regs_151_io_enable; // @[RegFile.scala 66:20:@51844.4]
  wire  regs_152_clock; // @[RegFile.scala 66:20:@51858.4]
  wire  regs_152_reset; // @[RegFile.scala 66:20:@51858.4]
  wire [63:0] regs_152_io_in; // @[RegFile.scala 66:20:@51858.4]
  wire  regs_152_io_reset; // @[RegFile.scala 66:20:@51858.4]
  wire [63:0] regs_152_io_out; // @[RegFile.scala 66:20:@51858.4]
  wire  regs_152_io_enable; // @[RegFile.scala 66:20:@51858.4]
  wire  regs_153_clock; // @[RegFile.scala 66:20:@51872.4]
  wire  regs_153_reset; // @[RegFile.scala 66:20:@51872.4]
  wire [63:0] regs_153_io_in; // @[RegFile.scala 66:20:@51872.4]
  wire  regs_153_io_reset; // @[RegFile.scala 66:20:@51872.4]
  wire [63:0] regs_153_io_out; // @[RegFile.scala 66:20:@51872.4]
  wire  regs_153_io_enable; // @[RegFile.scala 66:20:@51872.4]
  wire  regs_154_clock; // @[RegFile.scala 66:20:@51886.4]
  wire  regs_154_reset; // @[RegFile.scala 66:20:@51886.4]
  wire [63:0] regs_154_io_in; // @[RegFile.scala 66:20:@51886.4]
  wire  regs_154_io_reset; // @[RegFile.scala 66:20:@51886.4]
  wire [63:0] regs_154_io_out; // @[RegFile.scala 66:20:@51886.4]
  wire  regs_154_io_enable; // @[RegFile.scala 66:20:@51886.4]
  wire  regs_155_clock; // @[RegFile.scala 66:20:@51900.4]
  wire  regs_155_reset; // @[RegFile.scala 66:20:@51900.4]
  wire [63:0] regs_155_io_in; // @[RegFile.scala 66:20:@51900.4]
  wire  regs_155_io_reset; // @[RegFile.scala 66:20:@51900.4]
  wire [63:0] regs_155_io_out; // @[RegFile.scala 66:20:@51900.4]
  wire  regs_155_io_enable; // @[RegFile.scala 66:20:@51900.4]
  wire  regs_156_clock; // @[RegFile.scala 66:20:@51914.4]
  wire  regs_156_reset; // @[RegFile.scala 66:20:@51914.4]
  wire [63:0] regs_156_io_in; // @[RegFile.scala 66:20:@51914.4]
  wire  regs_156_io_reset; // @[RegFile.scala 66:20:@51914.4]
  wire [63:0] regs_156_io_out; // @[RegFile.scala 66:20:@51914.4]
  wire  regs_156_io_enable; // @[RegFile.scala 66:20:@51914.4]
  wire  regs_157_clock; // @[RegFile.scala 66:20:@51928.4]
  wire  regs_157_reset; // @[RegFile.scala 66:20:@51928.4]
  wire [63:0] regs_157_io_in; // @[RegFile.scala 66:20:@51928.4]
  wire  regs_157_io_reset; // @[RegFile.scala 66:20:@51928.4]
  wire [63:0] regs_157_io_out; // @[RegFile.scala 66:20:@51928.4]
  wire  regs_157_io_enable; // @[RegFile.scala 66:20:@51928.4]
  wire  regs_158_clock; // @[RegFile.scala 66:20:@51942.4]
  wire  regs_158_reset; // @[RegFile.scala 66:20:@51942.4]
  wire [63:0] regs_158_io_in; // @[RegFile.scala 66:20:@51942.4]
  wire  regs_158_io_reset; // @[RegFile.scala 66:20:@51942.4]
  wire [63:0] regs_158_io_out; // @[RegFile.scala 66:20:@51942.4]
  wire  regs_158_io_enable; // @[RegFile.scala 66:20:@51942.4]
  wire  regs_159_clock; // @[RegFile.scala 66:20:@51956.4]
  wire  regs_159_reset; // @[RegFile.scala 66:20:@51956.4]
  wire [63:0] regs_159_io_in; // @[RegFile.scala 66:20:@51956.4]
  wire  regs_159_io_reset; // @[RegFile.scala 66:20:@51956.4]
  wire [63:0] regs_159_io_out; // @[RegFile.scala 66:20:@51956.4]
  wire  regs_159_io_enable; // @[RegFile.scala 66:20:@51956.4]
  wire  regs_160_clock; // @[RegFile.scala 66:20:@51970.4]
  wire  regs_160_reset; // @[RegFile.scala 66:20:@51970.4]
  wire [63:0] regs_160_io_in; // @[RegFile.scala 66:20:@51970.4]
  wire  regs_160_io_reset; // @[RegFile.scala 66:20:@51970.4]
  wire [63:0] regs_160_io_out; // @[RegFile.scala 66:20:@51970.4]
  wire  regs_160_io_enable; // @[RegFile.scala 66:20:@51970.4]
  wire  regs_161_clock; // @[RegFile.scala 66:20:@51984.4]
  wire  regs_161_reset; // @[RegFile.scala 66:20:@51984.4]
  wire [63:0] regs_161_io_in; // @[RegFile.scala 66:20:@51984.4]
  wire  regs_161_io_reset; // @[RegFile.scala 66:20:@51984.4]
  wire [63:0] regs_161_io_out; // @[RegFile.scala 66:20:@51984.4]
  wire  regs_161_io_enable; // @[RegFile.scala 66:20:@51984.4]
  wire  regs_162_clock; // @[RegFile.scala 66:20:@51998.4]
  wire  regs_162_reset; // @[RegFile.scala 66:20:@51998.4]
  wire [63:0] regs_162_io_in; // @[RegFile.scala 66:20:@51998.4]
  wire  regs_162_io_reset; // @[RegFile.scala 66:20:@51998.4]
  wire [63:0] regs_162_io_out; // @[RegFile.scala 66:20:@51998.4]
  wire  regs_162_io_enable; // @[RegFile.scala 66:20:@51998.4]
  wire  regs_163_clock; // @[RegFile.scala 66:20:@52012.4]
  wire  regs_163_reset; // @[RegFile.scala 66:20:@52012.4]
  wire [63:0] regs_163_io_in; // @[RegFile.scala 66:20:@52012.4]
  wire  regs_163_io_reset; // @[RegFile.scala 66:20:@52012.4]
  wire [63:0] regs_163_io_out; // @[RegFile.scala 66:20:@52012.4]
  wire  regs_163_io_enable; // @[RegFile.scala 66:20:@52012.4]
  wire  regs_164_clock; // @[RegFile.scala 66:20:@52026.4]
  wire  regs_164_reset; // @[RegFile.scala 66:20:@52026.4]
  wire [63:0] regs_164_io_in; // @[RegFile.scala 66:20:@52026.4]
  wire  regs_164_io_reset; // @[RegFile.scala 66:20:@52026.4]
  wire [63:0] regs_164_io_out; // @[RegFile.scala 66:20:@52026.4]
  wire  regs_164_io_enable; // @[RegFile.scala 66:20:@52026.4]
  wire  regs_165_clock; // @[RegFile.scala 66:20:@52040.4]
  wire  regs_165_reset; // @[RegFile.scala 66:20:@52040.4]
  wire [63:0] regs_165_io_in; // @[RegFile.scala 66:20:@52040.4]
  wire  regs_165_io_reset; // @[RegFile.scala 66:20:@52040.4]
  wire [63:0] regs_165_io_out; // @[RegFile.scala 66:20:@52040.4]
  wire  regs_165_io_enable; // @[RegFile.scala 66:20:@52040.4]
  wire  regs_166_clock; // @[RegFile.scala 66:20:@52054.4]
  wire  regs_166_reset; // @[RegFile.scala 66:20:@52054.4]
  wire [63:0] regs_166_io_in; // @[RegFile.scala 66:20:@52054.4]
  wire  regs_166_io_reset; // @[RegFile.scala 66:20:@52054.4]
  wire [63:0] regs_166_io_out; // @[RegFile.scala 66:20:@52054.4]
  wire  regs_166_io_enable; // @[RegFile.scala 66:20:@52054.4]
  wire  regs_167_clock; // @[RegFile.scala 66:20:@52068.4]
  wire  regs_167_reset; // @[RegFile.scala 66:20:@52068.4]
  wire [63:0] regs_167_io_in; // @[RegFile.scala 66:20:@52068.4]
  wire  regs_167_io_reset; // @[RegFile.scala 66:20:@52068.4]
  wire [63:0] regs_167_io_out; // @[RegFile.scala 66:20:@52068.4]
  wire  regs_167_io_enable; // @[RegFile.scala 66:20:@52068.4]
  wire  regs_168_clock; // @[RegFile.scala 66:20:@52082.4]
  wire  regs_168_reset; // @[RegFile.scala 66:20:@52082.4]
  wire [63:0] regs_168_io_in; // @[RegFile.scala 66:20:@52082.4]
  wire  regs_168_io_reset; // @[RegFile.scala 66:20:@52082.4]
  wire [63:0] regs_168_io_out; // @[RegFile.scala 66:20:@52082.4]
  wire  regs_168_io_enable; // @[RegFile.scala 66:20:@52082.4]
  wire  regs_169_clock; // @[RegFile.scala 66:20:@52096.4]
  wire  regs_169_reset; // @[RegFile.scala 66:20:@52096.4]
  wire [63:0] regs_169_io_in; // @[RegFile.scala 66:20:@52096.4]
  wire  regs_169_io_reset; // @[RegFile.scala 66:20:@52096.4]
  wire [63:0] regs_169_io_out; // @[RegFile.scala 66:20:@52096.4]
  wire  regs_169_io_enable; // @[RegFile.scala 66:20:@52096.4]
  wire  regs_170_clock; // @[RegFile.scala 66:20:@52110.4]
  wire  regs_170_reset; // @[RegFile.scala 66:20:@52110.4]
  wire [63:0] regs_170_io_in; // @[RegFile.scala 66:20:@52110.4]
  wire  regs_170_io_reset; // @[RegFile.scala 66:20:@52110.4]
  wire [63:0] regs_170_io_out; // @[RegFile.scala 66:20:@52110.4]
  wire  regs_170_io_enable; // @[RegFile.scala 66:20:@52110.4]
  wire  regs_171_clock; // @[RegFile.scala 66:20:@52124.4]
  wire  regs_171_reset; // @[RegFile.scala 66:20:@52124.4]
  wire [63:0] regs_171_io_in; // @[RegFile.scala 66:20:@52124.4]
  wire  regs_171_io_reset; // @[RegFile.scala 66:20:@52124.4]
  wire [63:0] regs_171_io_out; // @[RegFile.scala 66:20:@52124.4]
  wire  regs_171_io_enable; // @[RegFile.scala 66:20:@52124.4]
  wire  regs_172_clock; // @[RegFile.scala 66:20:@52138.4]
  wire  regs_172_reset; // @[RegFile.scala 66:20:@52138.4]
  wire [63:0] regs_172_io_in; // @[RegFile.scala 66:20:@52138.4]
  wire  regs_172_io_reset; // @[RegFile.scala 66:20:@52138.4]
  wire [63:0] regs_172_io_out; // @[RegFile.scala 66:20:@52138.4]
  wire  regs_172_io_enable; // @[RegFile.scala 66:20:@52138.4]
  wire  regs_173_clock; // @[RegFile.scala 66:20:@52152.4]
  wire  regs_173_reset; // @[RegFile.scala 66:20:@52152.4]
  wire [63:0] regs_173_io_in; // @[RegFile.scala 66:20:@52152.4]
  wire  regs_173_io_reset; // @[RegFile.scala 66:20:@52152.4]
  wire [63:0] regs_173_io_out; // @[RegFile.scala 66:20:@52152.4]
  wire  regs_173_io_enable; // @[RegFile.scala 66:20:@52152.4]
  wire  regs_174_clock; // @[RegFile.scala 66:20:@52166.4]
  wire  regs_174_reset; // @[RegFile.scala 66:20:@52166.4]
  wire [63:0] regs_174_io_in; // @[RegFile.scala 66:20:@52166.4]
  wire  regs_174_io_reset; // @[RegFile.scala 66:20:@52166.4]
  wire [63:0] regs_174_io_out; // @[RegFile.scala 66:20:@52166.4]
  wire  regs_174_io_enable; // @[RegFile.scala 66:20:@52166.4]
  wire  regs_175_clock; // @[RegFile.scala 66:20:@52180.4]
  wire  regs_175_reset; // @[RegFile.scala 66:20:@52180.4]
  wire [63:0] regs_175_io_in; // @[RegFile.scala 66:20:@52180.4]
  wire  regs_175_io_reset; // @[RegFile.scala 66:20:@52180.4]
  wire [63:0] regs_175_io_out; // @[RegFile.scala 66:20:@52180.4]
  wire  regs_175_io_enable; // @[RegFile.scala 66:20:@52180.4]
  wire  regs_176_clock; // @[RegFile.scala 66:20:@52194.4]
  wire  regs_176_reset; // @[RegFile.scala 66:20:@52194.4]
  wire [63:0] regs_176_io_in; // @[RegFile.scala 66:20:@52194.4]
  wire  regs_176_io_reset; // @[RegFile.scala 66:20:@52194.4]
  wire [63:0] regs_176_io_out; // @[RegFile.scala 66:20:@52194.4]
  wire  regs_176_io_enable; // @[RegFile.scala 66:20:@52194.4]
  wire  regs_177_clock; // @[RegFile.scala 66:20:@52208.4]
  wire  regs_177_reset; // @[RegFile.scala 66:20:@52208.4]
  wire [63:0] regs_177_io_in; // @[RegFile.scala 66:20:@52208.4]
  wire  regs_177_io_reset; // @[RegFile.scala 66:20:@52208.4]
  wire [63:0] regs_177_io_out; // @[RegFile.scala 66:20:@52208.4]
  wire  regs_177_io_enable; // @[RegFile.scala 66:20:@52208.4]
  wire  regs_178_clock; // @[RegFile.scala 66:20:@52222.4]
  wire  regs_178_reset; // @[RegFile.scala 66:20:@52222.4]
  wire [63:0] regs_178_io_in; // @[RegFile.scala 66:20:@52222.4]
  wire  regs_178_io_reset; // @[RegFile.scala 66:20:@52222.4]
  wire [63:0] regs_178_io_out; // @[RegFile.scala 66:20:@52222.4]
  wire  regs_178_io_enable; // @[RegFile.scala 66:20:@52222.4]
  wire  regs_179_clock; // @[RegFile.scala 66:20:@52236.4]
  wire  regs_179_reset; // @[RegFile.scala 66:20:@52236.4]
  wire [63:0] regs_179_io_in; // @[RegFile.scala 66:20:@52236.4]
  wire  regs_179_io_reset; // @[RegFile.scala 66:20:@52236.4]
  wire [63:0] regs_179_io_out; // @[RegFile.scala 66:20:@52236.4]
  wire  regs_179_io_enable; // @[RegFile.scala 66:20:@52236.4]
  wire  regs_180_clock; // @[RegFile.scala 66:20:@52250.4]
  wire  regs_180_reset; // @[RegFile.scala 66:20:@52250.4]
  wire [63:0] regs_180_io_in; // @[RegFile.scala 66:20:@52250.4]
  wire  regs_180_io_reset; // @[RegFile.scala 66:20:@52250.4]
  wire [63:0] regs_180_io_out; // @[RegFile.scala 66:20:@52250.4]
  wire  regs_180_io_enable; // @[RegFile.scala 66:20:@52250.4]
  wire  regs_181_clock; // @[RegFile.scala 66:20:@52264.4]
  wire  regs_181_reset; // @[RegFile.scala 66:20:@52264.4]
  wire [63:0] regs_181_io_in; // @[RegFile.scala 66:20:@52264.4]
  wire  regs_181_io_reset; // @[RegFile.scala 66:20:@52264.4]
  wire [63:0] regs_181_io_out; // @[RegFile.scala 66:20:@52264.4]
  wire  regs_181_io_enable; // @[RegFile.scala 66:20:@52264.4]
  wire  regs_182_clock; // @[RegFile.scala 66:20:@52278.4]
  wire  regs_182_reset; // @[RegFile.scala 66:20:@52278.4]
  wire [63:0] regs_182_io_in; // @[RegFile.scala 66:20:@52278.4]
  wire  regs_182_io_reset; // @[RegFile.scala 66:20:@52278.4]
  wire [63:0] regs_182_io_out; // @[RegFile.scala 66:20:@52278.4]
  wire  regs_182_io_enable; // @[RegFile.scala 66:20:@52278.4]
  wire  regs_183_clock; // @[RegFile.scala 66:20:@52292.4]
  wire  regs_183_reset; // @[RegFile.scala 66:20:@52292.4]
  wire [63:0] regs_183_io_in; // @[RegFile.scala 66:20:@52292.4]
  wire  regs_183_io_reset; // @[RegFile.scala 66:20:@52292.4]
  wire [63:0] regs_183_io_out; // @[RegFile.scala 66:20:@52292.4]
  wire  regs_183_io_enable; // @[RegFile.scala 66:20:@52292.4]
  wire  regs_184_clock; // @[RegFile.scala 66:20:@52306.4]
  wire  regs_184_reset; // @[RegFile.scala 66:20:@52306.4]
  wire [63:0] regs_184_io_in; // @[RegFile.scala 66:20:@52306.4]
  wire  regs_184_io_reset; // @[RegFile.scala 66:20:@52306.4]
  wire [63:0] regs_184_io_out; // @[RegFile.scala 66:20:@52306.4]
  wire  regs_184_io_enable; // @[RegFile.scala 66:20:@52306.4]
  wire  regs_185_clock; // @[RegFile.scala 66:20:@52320.4]
  wire  regs_185_reset; // @[RegFile.scala 66:20:@52320.4]
  wire [63:0] regs_185_io_in; // @[RegFile.scala 66:20:@52320.4]
  wire  regs_185_io_reset; // @[RegFile.scala 66:20:@52320.4]
  wire [63:0] regs_185_io_out; // @[RegFile.scala 66:20:@52320.4]
  wire  regs_185_io_enable; // @[RegFile.scala 66:20:@52320.4]
  wire  regs_186_clock; // @[RegFile.scala 66:20:@52334.4]
  wire  regs_186_reset; // @[RegFile.scala 66:20:@52334.4]
  wire [63:0] regs_186_io_in; // @[RegFile.scala 66:20:@52334.4]
  wire  regs_186_io_reset; // @[RegFile.scala 66:20:@52334.4]
  wire [63:0] regs_186_io_out; // @[RegFile.scala 66:20:@52334.4]
  wire  regs_186_io_enable; // @[RegFile.scala 66:20:@52334.4]
  wire  regs_187_clock; // @[RegFile.scala 66:20:@52348.4]
  wire  regs_187_reset; // @[RegFile.scala 66:20:@52348.4]
  wire [63:0] regs_187_io_in; // @[RegFile.scala 66:20:@52348.4]
  wire  regs_187_io_reset; // @[RegFile.scala 66:20:@52348.4]
  wire [63:0] regs_187_io_out; // @[RegFile.scala 66:20:@52348.4]
  wire  regs_187_io_enable; // @[RegFile.scala 66:20:@52348.4]
  wire  regs_188_clock; // @[RegFile.scala 66:20:@52362.4]
  wire  regs_188_reset; // @[RegFile.scala 66:20:@52362.4]
  wire [63:0] regs_188_io_in; // @[RegFile.scala 66:20:@52362.4]
  wire  regs_188_io_reset; // @[RegFile.scala 66:20:@52362.4]
  wire [63:0] regs_188_io_out; // @[RegFile.scala 66:20:@52362.4]
  wire  regs_188_io_enable; // @[RegFile.scala 66:20:@52362.4]
  wire  regs_189_clock; // @[RegFile.scala 66:20:@52376.4]
  wire  regs_189_reset; // @[RegFile.scala 66:20:@52376.4]
  wire [63:0] regs_189_io_in; // @[RegFile.scala 66:20:@52376.4]
  wire  regs_189_io_reset; // @[RegFile.scala 66:20:@52376.4]
  wire [63:0] regs_189_io_out; // @[RegFile.scala 66:20:@52376.4]
  wire  regs_189_io_enable; // @[RegFile.scala 66:20:@52376.4]
  wire  regs_190_clock; // @[RegFile.scala 66:20:@52390.4]
  wire  regs_190_reset; // @[RegFile.scala 66:20:@52390.4]
  wire [63:0] regs_190_io_in; // @[RegFile.scala 66:20:@52390.4]
  wire  regs_190_io_reset; // @[RegFile.scala 66:20:@52390.4]
  wire [63:0] regs_190_io_out; // @[RegFile.scala 66:20:@52390.4]
  wire  regs_190_io_enable; // @[RegFile.scala 66:20:@52390.4]
  wire  regs_191_clock; // @[RegFile.scala 66:20:@52404.4]
  wire  regs_191_reset; // @[RegFile.scala 66:20:@52404.4]
  wire [63:0] regs_191_io_in; // @[RegFile.scala 66:20:@52404.4]
  wire  regs_191_io_reset; // @[RegFile.scala 66:20:@52404.4]
  wire [63:0] regs_191_io_out; // @[RegFile.scala 66:20:@52404.4]
  wire  regs_191_io_enable; // @[RegFile.scala 66:20:@52404.4]
  wire  regs_192_clock; // @[RegFile.scala 66:20:@52418.4]
  wire  regs_192_reset; // @[RegFile.scala 66:20:@52418.4]
  wire [63:0] regs_192_io_in; // @[RegFile.scala 66:20:@52418.4]
  wire  regs_192_io_reset; // @[RegFile.scala 66:20:@52418.4]
  wire [63:0] regs_192_io_out; // @[RegFile.scala 66:20:@52418.4]
  wire  regs_192_io_enable; // @[RegFile.scala 66:20:@52418.4]
  wire  regs_193_clock; // @[RegFile.scala 66:20:@52432.4]
  wire  regs_193_reset; // @[RegFile.scala 66:20:@52432.4]
  wire [63:0] regs_193_io_in; // @[RegFile.scala 66:20:@52432.4]
  wire  regs_193_io_reset; // @[RegFile.scala 66:20:@52432.4]
  wire [63:0] regs_193_io_out; // @[RegFile.scala 66:20:@52432.4]
  wire  regs_193_io_enable; // @[RegFile.scala 66:20:@52432.4]
  wire  regs_194_clock; // @[RegFile.scala 66:20:@52446.4]
  wire  regs_194_reset; // @[RegFile.scala 66:20:@52446.4]
  wire [63:0] regs_194_io_in; // @[RegFile.scala 66:20:@52446.4]
  wire  regs_194_io_reset; // @[RegFile.scala 66:20:@52446.4]
  wire [63:0] regs_194_io_out; // @[RegFile.scala 66:20:@52446.4]
  wire  regs_194_io_enable; // @[RegFile.scala 66:20:@52446.4]
  wire  regs_195_clock; // @[RegFile.scala 66:20:@52460.4]
  wire  regs_195_reset; // @[RegFile.scala 66:20:@52460.4]
  wire [63:0] regs_195_io_in; // @[RegFile.scala 66:20:@52460.4]
  wire  regs_195_io_reset; // @[RegFile.scala 66:20:@52460.4]
  wire [63:0] regs_195_io_out; // @[RegFile.scala 66:20:@52460.4]
  wire  regs_195_io_enable; // @[RegFile.scala 66:20:@52460.4]
  wire  regs_196_clock; // @[RegFile.scala 66:20:@52474.4]
  wire  regs_196_reset; // @[RegFile.scala 66:20:@52474.4]
  wire [63:0] regs_196_io_in; // @[RegFile.scala 66:20:@52474.4]
  wire  regs_196_io_reset; // @[RegFile.scala 66:20:@52474.4]
  wire [63:0] regs_196_io_out; // @[RegFile.scala 66:20:@52474.4]
  wire  regs_196_io_enable; // @[RegFile.scala 66:20:@52474.4]
  wire  regs_197_clock; // @[RegFile.scala 66:20:@52488.4]
  wire  regs_197_reset; // @[RegFile.scala 66:20:@52488.4]
  wire [63:0] regs_197_io_in; // @[RegFile.scala 66:20:@52488.4]
  wire  regs_197_io_reset; // @[RegFile.scala 66:20:@52488.4]
  wire [63:0] regs_197_io_out; // @[RegFile.scala 66:20:@52488.4]
  wire  regs_197_io_enable; // @[RegFile.scala 66:20:@52488.4]
  wire  regs_198_clock; // @[RegFile.scala 66:20:@52502.4]
  wire  regs_198_reset; // @[RegFile.scala 66:20:@52502.4]
  wire [63:0] regs_198_io_in; // @[RegFile.scala 66:20:@52502.4]
  wire  regs_198_io_reset; // @[RegFile.scala 66:20:@52502.4]
  wire [63:0] regs_198_io_out; // @[RegFile.scala 66:20:@52502.4]
  wire  regs_198_io_enable; // @[RegFile.scala 66:20:@52502.4]
  wire  regs_199_clock; // @[RegFile.scala 66:20:@52516.4]
  wire  regs_199_reset; // @[RegFile.scala 66:20:@52516.4]
  wire [63:0] regs_199_io_in; // @[RegFile.scala 66:20:@52516.4]
  wire  regs_199_io_reset; // @[RegFile.scala 66:20:@52516.4]
  wire [63:0] regs_199_io_out; // @[RegFile.scala 66:20:@52516.4]
  wire  regs_199_io_enable; // @[RegFile.scala 66:20:@52516.4]
  wire  regs_200_clock; // @[RegFile.scala 66:20:@52530.4]
  wire  regs_200_reset; // @[RegFile.scala 66:20:@52530.4]
  wire [63:0] regs_200_io_in; // @[RegFile.scala 66:20:@52530.4]
  wire  regs_200_io_reset; // @[RegFile.scala 66:20:@52530.4]
  wire [63:0] regs_200_io_out; // @[RegFile.scala 66:20:@52530.4]
  wire  regs_200_io_enable; // @[RegFile.scala 66:20:@52530.4]
  wire  regs_201_clock; // @[RegFile.scala 66:20:@52544.4]
  wire  regs_201_reset; // @[RegFile.scala 66:20:@52544.4]
  wire [63:0] regs_201_io_in; // @[RegFile.scala 66:20:@52544.4]
  wire  regs_201_io_reset; // @[RegFile.scala 66:20:@52544.4]
  wire [63:0] regs_201_io_out; // @[RegFile.scala 66:20:@52544.4]
  wire  regs_201_io_enable; // @[RegFile.scala 66:20:@52544.4]
  wire  regs_202_clock; // @[RegFile.scala 66:20:@52558.4]
  wire  regs_202_reset; // @[RegFile.scala 66:20:@52558.4]
  wire [63:0] regs_202_io_in; // @[RegFile.scala 66:20:@52558.4]
  wire  regs_202_io_reset; // @[RegFile.scala 66:20:@52558.4]
  wire [63:0] regs_202_io_out; // @[RegFile.scala 66:20:@52558.4]
  wire  regs_202_io_enable; // @[RegFile.scala 66:20:@52558.4]
  wire  regs_203_clock; // @[RegFile.scala 66:20:@52572.4]
  wire  regs_203_reset; // @[RegFile.scala 66:20:@52572.4]
  wire [63:0] regs_203_io_in; // @[RegFile.scala 66:20:@52572.4]
  wire  regs_203_io_reset; // @[RegFile.scala 66:20:@52572.4]
  wire [63:0] regs_203_io_out; // @[RegFile.scala 66:20:@52572.4]
  wire  regs_203_io_enable; // @[RegFile.scala 66:20:@52572.4]
  wire  regs_204_clock; // @[RegFile.scala 66:20:@52586.4]
  wire  regs_204_reset; // @[RegFile.scala 66:20:@52586.4]
  wire [63:0] regs_204_io_in; // @[RegFile.scala 66:20:@52586.4]
  wire  regs_204_io_reset; // @[RegFile.scala 66:20:@52586.4]
  wire [63:0] regs_204_io_out; // @[RegFile.scala 66:20:@52586.4]
  wire  regs_204_io_enable; // @[RegFile.scala 66:20:@52586.4]
  wire  regs_205_clock; // @[RegFile.scala 66:20:@52600.4]
  wire  regs_205_reset; // @[RegFile.scala 66:20:@52600.4]
  wire [63:0] regs_205_io_in; // @[RegFile.scala 66:20:@52600.4]
  wire  regs_205_io_reset; // @[RegFile.scala 66:20:@52600.4]
  wire [63:0] regs_205_io_out; // @[RegFile.scala 66:20:@52600.4]
  wire  regs_205_io_enable; // @[RegFile.scala 66:20:@52600.4]
  wire  regs_206_clock; // @[RegFile.scala 66:20:@52614.4]
  wire  regs_206_reset; // @[RegFile.scala 66:20:@52614.4]
  wire [63:0] regs_206_io_in; // @[RegFile.scala 66:20:@52614.4]
  wire  regs_206_io_reset; // @[RegFile.scala 66:20:@52614.4]
  wire [63:0] regs_206_io_out; // @[RegFile.scala 66:20:@52614.4]
  wire  regs_206_io_enable; // @[RegFile.scala 66:20:@52614.4]
  wire  regs_207_clock; // @[RegFile.scala 66:20:@52628.4]
  wire  regs_207_reset; // @[RegFile.scala 66:20:@52628.4]
  wire [63:0] regs_207_io_in; // @[RegFile.scala 66:20:@52628.4]
  wire  regs_207_io_reset; // @[RegFile.scala 66:20:@52628.4]
  wire [63:0] regs_207_io_out; // @[RegFile.scala 66:20:@52628.4]
  wire  regs_207_io_enable; // @[RegFile.scala 66:20:@52628.4]
  wire  regs_208_clock; // @[RegFile.scala 66:20:@52642.4]
  wire  regs_208_reset; // @[RegFile.scala 66:20:@52642.4]
  wire [63:0] regs_208_io_in; // @[RegFile.scala 66:20:@52642.4]
  wire  regs_208_io_reset; // @[RegFile.scala 66:20:@52642.4]
  wire [63:0] regs_208_io_out; // @[RegFile.scala 66:20:@52642.4]
  wire  regs_208_io_enable; // @[RegFile.scala 66:20:@52642.4]
  wire  regs_209_clock; // @[RegFile.scala 66:20:@52656.4]
  wire  regs_209_reset; // @[RegFile.scala 66:20:@52656.4]
  wire [63:0] regs_209_io_in; // @[RegFile.scala 66:20:@52656.4]
  wire  regs_209_io_reset; // @[RegFile.scala 66:20:@52656.4]
  wire [63:0] regs_209_io_out; // @[RegFile.scala 66:20:@52656.4]
  wire  regs_209_io_enable; // @[RegFile.scala 66:20:@52656.4]
  wire  regs_210_clock; // @[RegFile.scala 66:20:@52670.4]
  wire  regs_210_reset; // @[RegFile.scala 66:20:@52670.4]
  wire [63:0] regs_210_io_in; // @[RegFile.scala 66:20:@52670.4]
  wire  regs_210_io_reset; // @[RegFile.scala 66:20:@52670.4]
  wire [63:0] regs_210_io_out; // @[RegFile.scala 66:20:@52670.4]
  wire  regs_210_io_enable; // @[RegFile.scala 66:20:@52670.4]
  wire  regs_211_clock; // @[RegFile.scala 66:20:@52684.4]
  wire  regs_211_reset; // @[RegFile.scala 66:20:@52684.4]
  wire [63:0] regs_211_io_in; // @[RegFile.scala 66:20:@52684.4]
  wire  regs_211_io_reset; // @[RegFile.scala 66:20:@52684.4]
  wire [63:0] regs_211_io_out; // @[RegFile.scala 66:20:@52684.4]
  wire  regs_211_io_enable; // @[RegFile.scala 66:20:@52684.4]
  wire  regs_212_clock; // @[RegFile.scala 66:20:@52698.4]
  wire  regs_212_reset; // @[RegFile.scala 66:20:@52698.4]
  wire [63:0] regs_212_io_in; // @[RegFile.scala 66:20:@52698.4]
  wire  regs_212_io_reset; // @[RegFile.scala 66:20:@52698.4]
  wire [63:0] regs_212_io_out; // @[RegFile.scala 66:20:@52698.4]
  wire  regs_212_io_enable; // @[RegFile.scala 66:20:@52698.4]
  wire  regs_213_clock; // @[RegFile.scala 66:20:@52712.4]
  wire  regs_213_reset; // @[RegFile.scala 66:20:@52712.4]
  wire [63:0] regs_213_io_in; // @[RegFile.scala 66:20:@52712.4]
  wire  regs_213_io_reset; // @[RegFile.scala 66:20:@52712.4]
  wire [63:0] regs_213_io_out; // @[RegFile.scala 66:20:@52712.4]
  wire  regs_213_io_enable; // @[RegFile.scala 66:20:@52712.4]
  wire  regs_214_clock; // @[RegFile.scala 66:20:@52726.4]
  wire  regs_214_reset; // @[RegFile.scala 66:20:@52726.4]
  wire [63:0] regs_214_io_in; // @[RegFile.scala 66:20:@52726.4]
  wire  regs_214_io_reset; // @[RegFile.scala 66:20:@52726.4]
  wire [63:0] regs_214_io_out; // @[RegFile.scala 66:20:@52726.4]
  wire  regs_214_io_enable; // @[RegFile.scala 66:20:@52726.4]
  wire  regs_215_clock; // @[RegFile.scala 66:20:@52740.4]
  wire  regs_215_reset; // @[RegFile.scala 66:20:@52740.4]
  wire [63:0] regs_215_io_in; // @[RegFile.scala 66:20:@52740.4]
  wire  regs_215_io_reset; // @[RegFile.scala 66:20:@52740.4]
  wire [63:0] regs_215_io_out; // @[RegFile.scala 66:20:@52740.4]
  wire  regs_215_io_enable; // @[RegFile.scala 66:20:@52740.4]
  wire  regs_216_clock; // @[RegFile.scala 66:20:@52754.4]
  wire  regs_216_reset; // @[RegFile.scala 66:20:@52754.4]
  wire [63:0] regs_216_io_in; // @[RegFile.scala 66:20:@52754.4]
  wire  regs_216_io_reset; // @[RegFile.scala 66:20:@52754.4]
  wire [63:0] regs_216_io_out; // @[RegFile.scala 66:20:@52754.4]
  wire  regs_216_io_enable; // @[RegFile.scala 66:20:@52754.4]
  wire  regs_217_clock; // @[RegFile.scala 66:20:@52768.4]
  wire  regs_217_reset; // @[RegFile.scala 66:20:@52768.4]
  wire [63:0] regs_217_io_in; // @[RegFile.scala 66:20:@52768.4]
  wire  regs_217_io_reset; // @[RegFile.scala 66:20:@52768.4]
  wire [63:0] regs_217_io_out; // @[RegFile.scala 66:20:@52768.4]
  wire  regs_217_io_enable; // @[RegFile.scala 66:20:@52768.4]
  wire  regs_218_clock; // @[RegFile.scala 66:20:@52782.4]
  wire  regs_218_reset; // @[RegFile.scala 66:20:@52782.4]
  wire [63:0] regs_218_io_in; // @[RegFile.scala 66:20:@52782.4]
  wire  regs_218_io_reset; // @[RegFile.scala 66:20:@52782.4]
  wire [63:0] regs_218_io_out; // @[RegFile.scala 66:20:@52782.4]
  wire  regs_218_io_enable; // @[RegFile.scala 66:20:@52782.4]
  wire  regs_219_clock; // @[RegFile.scala 66:20:@52796.4]
  wire  regs_219_reset; // @[RegFile.scala 66:20:@52796.4]
  wire [63:0] regs_219_io_in; // @[RegFile.scala 66:20:@52796.4]
  wire  regs_219_io_reset; // @[RegFile.scala 66:20:@52796.4]
  wire [63:0] regs_219_io_out; // @[RegFile.scala 66:20:@52796.4]
  wire  regs_219_io_enable; // @[RegFile.scala 66:20:@52796.4]
  wire  regs_220_clock; // @[RegFile.scala 66:20:@52810.4]
  wire  regs_220_reset; // @[RegFile.scala 66:20:@52810.4]
  wire [63:0] regs_220_io_in; // @[RegFile.scala 66:20:@52810.4]
  wire  regs_220_io_reset; // @[RegFile.scala 66:20:@52810.4]
  wire [63:0] regs_220_io_out; // @[RegFile.scala 66:20:@52810.4]
  wire  regs_220_io_enable; // @[RegFile.scala 66:20:@52810.4]
  wire  regs_221_clock; // @[RegFile.scala 66:20:@52824.4]
  wire  regs_221_reset; // @[RegFile.scala 66:20:@52824.4]
  wire [63:0] regs_221_io_in; // @[RegFile.scala 66:20:@52824.4]
  wire  regs_221_io_reset; // @[RegFile.scala 66:20:@52824.4]
  wire [63:0] regs_221_io_out; // @[RegFile.scala 66:20:@52824.4]
  wire  regs_221_io_enable; // @[RegFile.scala 66:20:@52824.4]
  wire  regs_222_clock; // @[RegFile.scala 66:20:@52838.4]
  wire  regs_222_reset; // @[RegFile.scala 66:20:@52838.4]
  wire [63:0] regs_222_io_in; // @[RegFile.scala 66:20:@52838.4]
  wire  regs_222_io_reset; // @[RegFile.scala 66:20:@52838.4]
  wire [63:0] regs_222_io_out; // @[RegFile.scala 66:20:@52838.4]
  wire  regs_222_io_enable; // @[RegFile.scala 66:20:@52838.4]
  wire  regs_223_clock; // @[RegFile.scala 66:20:@52852.4]
  wire  regs_223_reset; // @[RegFile.scala 66:20:@52852.4]
  wire [63:0] regs_223_io_in; // @[RegFile.scala 66:20:@52852.4]
  wire  regs_223_io_reset; // @[RegFile.scala 66:20:@52852.4]
  wire [63:0] regs_223_io_out; // @[RegFile.scala 66:20:@52852.4]
  wire  regs_223_io_enable; // @[RegFile.scala 66:20:@52852.4]
  wire  regs_224_clock; // @[RegFile.scala 66:20:@52866.4]
  wire  regs_224_reset; // @[RegFile.scala 66:20:@52866.4]
  wire [63:0] regs_224_io_in; // @[RegFile.scala 66:20:@52866.4]
  wire  regs_224_io_reset; // @[RegFile.scala 66:20:@52866.4]
  wire [63:0] regs_224_io_out; // @[RegFile.scala 66:20:@52866.4]
  wire  regs_224_io_enable; // @[RegFile.scala 66:20:@52866.4]
  wire  regs_225_clock; // @[RegFile.scala 66:20:@52880.4]
  wire  regs_225_reset; // @[RegFile.scala 66:20:@52880.4]
  wire [63:0] regs_225_io_in; // @[RegFile.scala 66:20:@52880.4]
  wire  regs_225_io_reset; // @[RegFile.scala 66:20:@52880.4]
  wire [63:0] regs_225_io_out; // @[RegFile.scala 66:20:@52880.4]
  wire  regs_225_io_enable; // @[RegFile.scala 66:20:@52880.4]
  wire  regs_226_clock; // @[RegFile.scala 66:20:@52894.4]
  wire  regs_226_reset; // @[RegFile.scala 66:20:@52894.4]
  wire [63:0] regs_226_io_in; // @[RegFile.scala 66:20:@52894.4]
  wire  regs_226_io_reset; // @[RegFile.scala 66:20:@52894.4]
  wire [63:0] regs_226_io_out; // @[RegFile.scala 66:20:@52894.4]
  wire  regs_226_io_enable; // @[RegFile.scala 66:20:@52894.4]
  wire  regs_227_clock; // @[RegFile.scala 66:20:@52908.4]
  wire  regs_227_reset; // @[RegFile.scala 66:20:@52908.4]
  wire [63:0] regs_227_io_in; // @[RegFile.scala 66:20:@52908.4]
  wire  regs_227_io_reset; // @[RegFile.scala 66:20:@52908.4]
  wire [63:0] regs_227_io_out; // @[RegFile.scala 66:20:@52908.4]
  wire  regs_227_io_enable; // @[RegFile.scala 66:20:@52908.4]
  wire  regs_228_clock; // @[RegFile.scala 66:20:@52922.4]
  wire  regs_228_reset; // @[RegFile.scala 66:20:@52922.4]
  wire [63:0] regs_228_io_in; // @[RegFile.scala 66:20:@52922.4]
  wire  regs_228_io_reset; // @[RegFile.scala 66:20:@52922.4]
  wire [63:0] regs_228_io_out; // @[RegFile.scala 66:20:@52922.4]
  wire  regs_228_io_enable; // @[RegFile.scala 66:20:@52922.4]
  wire  regs_229_clock; // @[RegFile.scala 66:20:@52936.4]
  wire  regs_229_reset; // @[RegFile.scala 66:20:@52936.4]
  wire [63:0] regs_229_io_in; // @[RegFile.scala 66:20:@52936.4]
  wire  regs_229_io_reset; // @[RegFile.scala 66:20:@52936.4]
  wire [63:0] regs_229_io_out; // @[RegFile.scala 66:20:@52936.4]
  wire  regs_229_io_enable; // @[RegFile.scala 66:20:@52936.4]
  wire  regs_230_clock; // @[RegFile.scala 66:20:@52950.4]
  wire  regs_230_reset; // @[RegFile.scala 66:20:@52950.4]
  wire [63:0] regs_230_io_in; // @[RegFile.scala 66:20:@52950.4]
  wire  regs_230_io_reset; // @[RegFile.scala 66:20:@52950.4]
  wire [63:0] regs_230_io_out; // @[RegFile.scala 66:20:@52950.4]
  wire  regs_230_io_enable; // @[RegFile.scala 66:20:@52950.4]
  wire  regs_231_clock; // @[RegFile.scala 66:20:@52964.4]
  wire  regs_231_reset; // @[RegFile.scala 66:20:@52964.4]
  wire [63:0] regs_231_io_in; // @[RegFile.scala 66:20:@52964.4]
  wire  regs_231_io_reset; // @[RegFile.scala 66:20:@52964.4]
  wire [63:0] regs_231_io_out; // @[RegFile.scala 66:20:@52964.4]
  wire  regs_231_io_enable; // @[RegFile.scala 66:20:@52964.4]
  wire  regs_232_clock; // @[RegFile.scala 66:20:@52978.4]
  wire  regs_232_reset; // @[RegFile.scala 66:20:@52978.4]
  wire [63:0] regs_232_io_in; // @[RegFile.scala 66:20:@52978.4]
  wire  regs_232_io_reset; // @[RegFile.scala 66:20:@52978.4]
  wire [63:0] regs_232_io_out; // @[RegFile.scala 66:20:@52978.4]
  wire  regs_232_io_enable; // @[RegFile.scala 66:20:@52978.4]
  wire  regs_233_clock; // @[RegFile.scala 66:20:@52992.4]
  wire  regs_233_reset; // @[RegFile.scala 66:20:@52992.4]
  wire [63:0] regs_233_io_in; // @[RegFile.scala 66:20:@52992.4]
  wire  regs_233_io_reset; // @[RegFile.scala 66:20:@52992.4]
  wire [63:0] regs_233_io_out; // @[RegFile.scala 66:20:@52992.4]
  wire  regs_233_io_enable; // @[RegFile.scala 66:20:@52992.4]
  wire  regs_234_clock; // @[RegFile.scala 66:20:@53006.4]
  wire  regs_234_reset; // @[RegFile.scala 66:20:@53006.4]
  wire [63:0] regs_234_io_in; // @[RegFile.scala 66:20:@53006.4]
  wire  regs_234_io_reset; // @[RegFile.scala 66:20:@53006.4]
  wire [63:0] regs_234_io_out; // @[RegFile.scala 66:20:@53006.4]
  wire  regs_234_io_enable; // @[RegFile.scala 66:20:@53006.4]
  wire  regs_235_clock; // @[RegFile.scala 66:20:@53020.4]
  wire  regs_235_reset; // @[RegFile.scala 66:20:@53020.4]
  wire [63:0] regs_235_io_in; // @[RegFile.scala 66:20:@53020.4]
  wire  regs_235_io_reset; // @[RegFile.scala 66:20:@53020.4]
  wire [63:0] regs_235_io_out; // @[RegFile.scala 66:20:@53020.4]
  wire  regs_235_io_enable; // @[RegFile.scala 66:20:@53020.4]
  wire  regs_236_clock; // @[RegFile.scala 66:20:@53034.4]
  wire  regs_236_reset; // @[RegFile.scala 66:20:@53034.4]
  wire [63:0] regs_236_io_in; // @[RegFile.scala 66:20:@53034.4]
  wire  regs_236_io_reset; // @[RegFile.scala 66:20:@53034.4]
  wire [63:0] regs_236_io_out; // @[RegFile.scala 66:20:@53034.4]
  wire  regs_236_io_enable; // @[RegFile.scala 66:20:@53034.4]
  wire  regs_237_clock; // @[RegFile.scala 66:20:@53048.4]
  wire  regs_237_reset; // @[RegFile.scala 66:20:@53048.4]
  wire [63:0] regs_237_io_in; // @[RegFile.scala 66:20:@53048.4]
  wire  regs_237_io_reset; // @[RegFile.scala 66:20:@53048.4]
  wire [63:0] regs_237_io_out; // @[RegFile.scala 66:20:@53048.4]
  wire  regs_237_io_enable; // @[RegFile.scala 66:20:@53048.4]
  wire  regs_238_clock; // @[RegFile.scala 66:20:@53062.4]
  wire  regs_238_reset; // @[RegFile.scala 66:20:@53062.4]
  wire [63:0] regs_238_io_in; // @[RegFile.scala 66:20:@53062.4]
  wire  regs_238_io_reset; // @[RegFile.scala 66:20:@53062.4]
  wire [63:0] regs_238_io_out; // @[RegFile.scala 66:20:@53062.4]
  wire  regs_238_io_enable; // @[RegFile.scala 66:20:@53062.4]
  wire  regs_239_clock; // @[RegFile.scala 66:20:@53076.4]
  wire  regs_239_reset; // @[RegFile.scala 66:20:@53076.4]
  wire [63:0] regs_239_io_in; // @[RegFile.scala 66:20:@53076.4]
  wire  regs_239_io_reset; // @[RegFile.scala 66:20:@53076.4]
  wire [63:0] regs_239_io_out; // @[RegFile.scala 66:20:@53076.4]
  wire  regs_239_io_enable; // @[RegFile.scala 66:20:@53076.4]
  wire  regs_240_clock; // @[RegFile.scala 66:20:@53090.4]
  wire  regs_240_reset; // @[RegFile.scala 66:20:@53090.4]
  wire [63:0] regs_240_io_in; // @[RegFile.scala 66:20:@53090.4]
  wire  regs_240_io_reset; // @[RegFile.scala 66:20:@53090.4]
  wire [63:0] regs_240_io_out; // @[RegFile.scala 66:20:@53090.4]
  wire  regs_240_io_enable; // @[RegFile.scala 66:20:@53090.4]
  wire  regs_241_clock; // @[RegFile.scala 66:20:@53104.4]
  wire  regs_241_reset; // @[RegFile.scala 66:20:@53104.4]
  wire [63:0] regs_241_io_in; // @[RegFile.scala 66:20:@53104.4]
  wire  regs_241_io_reset; // @[RegFile.scala 66:20:@53104.4]
  wire [63:0] regs_241_io_out; // @[RegFile.scala 66:20:@53104.4]
  wire  regs_241_io_enable; // @[RegFile.scala 66:20:@53104.4]
  wire  regs_242_clock; // @[RegFile.scala 66:20:@53118.4]
  wire  regs_242_reset; // @[RegFile.scala 66:20:@53118.4]
  wire [63:0] regs_242_io_in; // @[RegFile.scala 66:20:@53118.4]
  wire  regs_242_io_reset; // @[RegFile.scala 66:20:@53118.4]
  wire [63:0] regs_242_io_out; // @[RegFile.scala 66:20:@53118.4]
  wire  regs_242_io_enable; // @[RegFile.scala 66:20:@53118.4]
  wire  regs_243_clock; // @[RegFile.scala 66:20:@53132.4]
  wire  regs_243_reset; // @[RegFile.scala 66:20:@53132.4]
  wire [63:0] regs_243_io_in; // @[RegFile.scala 66:20:@53132.4]
  wire  regs_243_io_reset; // @[RegFile.scala 66:20:@53132.4]
  wire [63:0] regs_243_io_out; // @[RegFile.scala 66:20:@53132.4]
  wire  regs_243_io_enable; // @[RegFile.scala 66:20:@53132.4]
  wire  regs_244_clock; // @[RegFile.scala 66:20:@53146.4]
  wire  regs_244_reset; // @[RegFile.scala 66:20:@53146.4]
  wire [63:0] regs_244_io_in; // @[RegFile.scala 66:20:@53146.4]
  wire  regs_244_io_reset; // @[RegFile.scala 66:20:@53146.4]
  wire [63:0] regs_244_io_out; // @[RegFile.scala 66:20:@53146.4]
  wire  regs_244_io_enable; // @[RegFile.scala 66:20:@53146.4]
  wire  regs_245_clock; // @[RegFile.scala 66:20:@53160.4]
  wire  regs_245_reset; // @[RegFile.scala 66:20:@53160.4]
  wire [63:0] regs_245_io_in; // @[RegFile.scala 66:20:@53160.4]
  wire  regs_245_io_reset; // @[RegFile.scala 66:20:@53160.4]
  wire [63:0] regs_245_io_out; // @[RegFile.scala 66:20:@53160.4]
  wire  regs_245_io_enable; // @[RegFile.scala 66:20:@53160.4]
  wire  regs_246_clock; // @[RegFile.scala 66:20:@53174.4]
  wire  regs_246_reset; // @[RegFile.scala 66:20:@53174.4]
  wire [63:0] regs_246_io_in; // @[RegFile.scala 66:20:@53174.4]
  wire  regs_246_io_reset; // @[RegFile.scala 66:20:@53174.4]
  wire [63:0] regs_246_io_out; // @[RegFile.scala 66:20:@53174.4]
  wire  regs_246_io_enable; // @[RegFile.scala 66:20:@53174.4]
  wire  regs_247_clock; // @[RegFile.scala 66:20:@53188.4]
  wire  regs_247_reset; // @[RegFile.scala 66:20:@53188.4]
  wire [63:0] regs_247_io_in; // @[RegFile.scala 66:20:@53188.4]
  wire  regs_247_io_reset; // @[RegFile.scala 66:20:@53188.4]
  wire [63:0] regs_247_io_out; // @[RegFile.scala 66:20:@53188.4]
  wire  regs_247_io_enable; // @[RegFile.scala 66:20:@53188.4]
  wire  regs_248_clock; // @[RegFile.scala 66:20:@53202.4]
  wire  regs_248_reset; // @[RegFile.scala 66:20:@53202.4]
  wire [63:0] regs_248_io_in; // @[RegFile.scala 66:20:@53202.4]
  wire  regs_248_io_reset; // @[RegFile.scala 66:20:@53202.4]
  wire [63:0] regs_248_io_out; // @[RegFile.scala 66:20:@53202.4]
  wire  regs_248_io_enable; // @[RegFile.scala 66:20:@53202.4]
  wire  regs_249_clock; // @[RegFile.scala 66:20:@53216.4]
  wire  regs_249_reset; // @[RegFile.scala 66:20:@53216.4]
  wire [63:0] regs_249_io_in; // @[RegFile.scala 66:20:@53216.4]
  wire  regs_249_io_reset; // @[RegFile.scala 66:20:@53216.4]
  wire [63:0] regs_249_io_out; // @[RegFile.scala 66:20:@53216.4]
  wire  regs_249_io_enable; // @[RegFile.scala 66:20:@53216.4]
  wire  regs_250_clock; // @[RegFile.scala 66:20:@53230.4]
  wire  regs_250_reset; // @[RegFile.scala 66:20:@53230.4]
  wire [63:0] regs_250_io_in; // @[RegFile.scala 66:20:@53230.4]
  wire  regs_250_io_reset; // @[RegFile.scala 66:20:@53230.4]
  wire [63:0] regs_250_io_out; // @[RegFile.scala 66:20:@53230.4]
  wire  regs_250_io_enable; // @[RegFile.scala 66:20:@53230.4]
  wire  regs_251_clock; // @[RegFile.scala 66:20:@53244.4]
  wire  regs_251_reset; // @[RegFile.scala 66:20:@53244.4]
  wire [63:0] regs_251_io_in; // @[RegFile.scala 66:20:@53244.4]
  wire  regs_251_io_reset; // @[RegFile.scala 66:20:@53244.4]
  wire [63:0] regs_251_io_out; // @[RegFile.scala 66:20:@53244.4]
  wire  regs_251_io_enable; // @[RegFile.scala 66:20:@53244.4]
  wire  regs_252_clock; // @[RegFile.scala 66:20:@53258.4]
  wire  regs_252_reset; // @[RegFile.scala 66:20:@53258.4]
  wire [63:0] regs_252_io_in; // @[RegFile.scala 66:20:@53258.4]
  wire  regs_252_io_reset; // @[RegFile.scala 66:20:@53258.4]
  wire [63:0] regs_252_io_out; // @[RegFile.scala 66:20:@53258.4]
  wire  regs_252_io_enable; // @[RegFile.scala 66:20:@53258.4]
  wire  regs_253_clock; // @[RegFile.scala 66:20:@53272.4]
  wire  regs_253_reset; // @[RegFile.scala 66:20:@53272.4]
  wire [63:0] regs_253_io_in; // @[RegFile.scala 66:20:@53272.4]
  wire  regs_253_io_reset; // @[RegFile.scala 66:20:@53272.4]
  wire [63:0] regs_253_io_out; // @[RegFile.scala 66:20:@53272.4]
  wire  regs_253_io_enable; // @[RegFile.scala 66:20:@53272.4]
  wire  regs_254_clock; // @[RegFile.scala 66:20:@53286.4]
  wire  regs_254_reset; // @[RegFile.scala 66:20:@53286.4]
  wire [63:0] regs_254_io_in; // @[RegFile.scala 66:20:@53286.4]
  wire  regs_254_io_reset; // @[RegFile.scala 66:20:@53286.4]
  wire [63:0] regs_254_io_out; // @[RegFile.scala 66:20:@53286.4]
  wire  regs_254_io_enable; // @[RegFile.scala 66:20:@53286.4]
  wire  regs_255_clock; // @[RegFile.scala 66:20:@53300.4]
  wire  regs_255_reset; // @[RegFile.scala 66:20:@53300.4]
  wire [63:0] regs_255_io_in; // @[RegFile.scala 66:20:@53300.4]
  wire  regs_255_io_reset; // @[RegFile.scala 66:20:@53300.4]
  wire [63:0] regs_255_io_out; // @[RegFile.scala 66:20:@53300.4]
  wire  regs_255_io_enable; // @[RegFile.scala 66:20:@53300.4]
  wire  regs_256_clock; // @[RegFile.scala 66:20:@53314.4]
  wire  regs_256_reset; // @[RegFile.scala 66:20:@53314.4]
  wire [63:0] regs_256_io_in; // @[RegFile.scala 66:20:@53314.4]
  wire  regs_256_io_reset; // @[RegFile.scala 66:20:@53314.4]
  wire [63:0] regs_256_io_out; // @[RegFile.scala 66:20:@53314.4]
  wire  regs_256_io_enable; // @[RegFile.scala 66:20:@53314.4]
  wire  regs_257_clock; // @[RegFile.scala 66:20:@53328.4]
  wire  regs_257_reset; // @[RegFile.scala 66:20:@53328.4]
  wire [63:0] regs_257_io_in; // @[RegFile.scala 66:20:@53328.4]
  wire  regs_257_io_reset; // @[RegFile.scala 66:20:@53328.4]
  wire [63:0] regs_257_io_out; // @[RegFile.scala 66:20:@53328.4]
  wire  regs_257_io_enable; // @[RegFile.scala 66:20:@53328.4]
  wire  regs_258_clock; // @[RegFile.scala 66:20:@53342.4]
  wire  regs_258_reset; // @[RegFile.scala 66:20:@53342.4]
  wire [63:0] regs_258_io_in; // @[RegFile.scala 66:20:@53342.4]
  wire  regs_258_io_reset; // @[RegFile.scala 66:20:@53342.4]
  wire [63:0] regs_258_io_out; // @[RegFile.scala 66:20:@53342.4]
  wire  regs_258_io_enable; // @[RegFile.scala 66:20:@53342.4]
  wire  regs_259_clock; // @[RegFile.scala 66:20:@53356.4]
  wire  regs_259_reset; // @[RegFile.scala 66:20:@53356.4]
  wire [63:0] regs_259_io_in; // @[RegFile.scala 66:20:@53356.4]
  wire  regs_259_io_reset; // @[RegFile.scala 66:20:@53356.4]
  wire [63:0] regs_259_io_out; // @[RegFile.scala 66:20:@53356.4]
  wire  regs_259_io_enable; // @[RegFile.scala 66:20:@53356.4]
  wire  regs_260_clock; // @[RegFile.scala 66:20:@53370.4]
  wire  regs_260_reset; // @[RegFile.scala 66:20:@53370.4]
  wire [63:0] regs_260_io_in; // @[RegFile.scala 66:20:@53370.4]
  wire  regs_260_io_reset; // @[RegFile.scala 66:20:@53370.4]
  wire [63:0] regs_260_io_out; // @[RegFile.scala 66:20:@53370.4]
  wire  regs_260_io_enable; // @[RegFile.scala 66:20:@53370.4]
  wire  regs_261_clock; // @[RegFile.scala 66:20:@53384.4]
  wire  regs_261_reset; // @[RegFile.scala 66:20:@53384.4]
  wire [63:0] regs_261_io_in; // @[RegFile.scala 66:20:@53384.4]
  wire  regs_261_io_reset; // @[RegFile.scala 66:20:@53384.4]
  wire [63:0] regs_261_io_out; // @[RegFile.scala 66:20:@53384.4]
  wire  regs_261_io_enable; // @[RegFile.scala 66:20:@53384.4]
  wire  regs_262_clock; // @[RegFile.scala 66:20:@53398.4]
  wire  regs_262_reset; // @[RegFile.scala 66:20:@53398.4]
  wire [63:0] regs_262_io_in; // @[RegFile.scala 66:20:@53398.4]
  wire  regs_262_io_reset; // @[RegFile.scala 66:20:@53398.4]
  wire [63:0] regs_262_io_out; // @[RegFile.scala 66:20:@53398.4]
  wire  regs_262_io_enable; // @[RegFile.scala 66:20:@53398.4]
  wire  regs_263_clock; // @[RegFile.scala 66:20:@53412.4]
  wire  regs_263_reset; // @[RegFile.scala 66:20:@53412.4]
  wire [63:0] regs_263_io_in; // @[RegFile.scala 66:20:@53412.4]
  wire  regs_263_io_reset; // @[RegFile.scala 66:20:@53412.4]
  wire [63:0] regs_263_io_out; // @[RegFile.scala 66:20:@53412.4]
  wire  regs_263_io_enable; // @[RegFile.scala 66:20:@53412.4]
  wire  regs_264_clock; // @[RegFile.scala 66:20:@53426.4]
  wire  regs_264_reset; // @[RegFile.scala 66:20:@53426.4]
  wire [63:0] regs_264_io_in; // @[RegFile.scala 66:20:@53426.4]
  wire  regs_264_io_reset; // @[RegFile.scala 66:20:@53426.4]
  wire [63:0] regs_264_io_out; // @[RegFile.scala 66:20:@53426.4]
  wire  regs_264_io_enable; // @[RegFile.scala 66:20:@53426.4]
  wire  regs_265_clock; // @[RegFile.scala 66:20:@53440.4]
  wire  regs_265_reset; // @[RegFile.scala 66:20:@53440.4]
  wire [63:0] regs_265_io_in; // @[RegFile.scala 66:20:@53440.4]
  wire  regs_265_io_reset; // @[RegFile.scala 66:20:@53440.4]
  wire [63:0] regs_265_io_out; // @[RegFile.scala 66:20:@53440.4]
  wire  regs_265_io_enable; // @[RegFile.scala 66:20:@53440.4]
  wire  regs_266_clock; // @[RegFile.scala 66:20:@53454.4]
  wire  regs_266_reset; // @[RegFile.scala 66:20:@53454.4]
  wire [63:0] regs_266_io_in; // @[RegFile.scala 66:20:@53454.4]
  wire  regs_266_io_reset; // @[RegFile.scala 66:20:@53454.4]
  wire [63:0] regs_266_io_out; // @[RegFile.scala 66:20:@53454.4]
  wire  regs_266_io_enable; // @[RegFile.scala 66:20:@53454.4]
  wire  regs_267_clock; // @[RegFile.scala 66:20:@53468.4]
  wire  regs_267_reset; // @[RegFile.scala 66:20:@53468.4]
  wire [63:0] regs_267_io_in; // @[RegFile.scala 66:20:@53468.4]
  wire  regs_267_io_reset; // @[RegFile.scala 66:20:@53468.4]
  wire [63:0] regs_267_io_out; // @[RegFile.scala 66:20:@53468.4]
  wire  regs_267_io_enable; // @[RegFile.scala 66:20:@53468.4]
  wire  regs_268_clock; // @[RegFile.scala 66:20:@53482.4]
  wire  regs_268_reset; // @[RegFile.scala 66:20:@53482.4]
  wire [63:0] regs_268_io_in; // @[RegFile.scala 66:20:@53482.4]
  wire  regs_268_io_reset; // @[RegFile.scala 66:20:@53482.4]
  wire [63:0] regs_268_io_out; // @[RegFile.scala 66:20:@53482.4]
  wire  regs_268_io_enable; // @[RegFile.scala 66:20:@53482.4]
  wire  regs_269_clock; // @[RegFile.scala 66:20:@53496.4]
  wire  regs_269_reset; // @[RegFile.scala 66:20:@53496.4]
  wire [63:0] regs_269_io_in; // @[RegFile.scala 66:20:@53496.4]
  wire  regs_269_io_reset; // @[RegFile.scala 66:20:@53496.4]
  wire [63:0] regs_269_io_out; // @[RegFile.scala 66:20:@53496.4]
  wire  regs_269_io_enable; // @[RegFile.scala 66:20:@53496.4]
  wire  regs_270_clock; // @[RegFile.scala 66:20:@53510.4]
  wire  regs_270_reset; // @[RegFile.scala 66:20:@53510.4]
  wire [63:0] regs_270_io_in; // @[RegFile.scala 66:20:@53510.4]
  wire  regs_270_io_reset; // @[RegFile.scala 66:20:@53510.4]
  wire [63:0] regs_270_io_out; // @[RegFile.scala 66:20:@53510.4]
  wire  regs_270_io_enable; // @[RegFile.scala 66:20:@53510.4]
  wire  regs_271_clock; // @[RegFile.scala 66:20:@53524.4]
  wire  regs_271_reset; // @[RegFile.scala 66:20:@53524.4]
  wire [63:0] regs_271_io_in; // @[RegFile.scala 66:20:@53524.4]
  wire  regs_271_io_reset; // @[RegFile.scala 66:20:@53524.4]
  wire [63:0] regs_271_io_out; // @[RegFile.scala 66:20:@53524.4]
  wire  regs_271_io_enable; // @[RegFile.scala 66:20:@53524.4]
  wire  regs_272_clock; // @[RegFile.scala 66:20:@53538.4]
  wire  regs_272_reset; // @[RegFile.scala 66:20:@53538.4]
  wire [63:0] regs_272_io_in; // @[RegFile.scala 66:20:@53538.4]
  wire  regs_272_io_reset; // @[RegFile.scala 66:20:@53538.4]
  wire [63:0] regs_272_io_out; // @[RegFile.scala 66:20:@53538.4]
  wire  regs_272_io_enable; // @[RegFile.scala 66:20:@53538.4]
  wire  regs_273_clock; // @[RegFile.scala 66:20:@53552.4]
  wire  regs_273_reset; // @[RegFile.scala 66:20:@53552.4]
  wire [63:0] regs_273_io_in; // @[RegFile.scala 66:20:@53552.4]
  wire  regs_273_io_reset; // @[RegFile.scala 66:20:@53552.4]
  wire [63:0] regs_273_io_out; // @[RegFile.scala 66:20:@53552.4]
  wire  regs_273_io_enable; // @[RegFile.scala 66:20:@53552.4]
  wire  regs_274_clock; // @[RegFile.scala 66:20:@53566.4]
  wire  regs_274_reset; // @[RegFile.scala 66:20:@53566.4]
  wire [63:0] regs_274_io_in; // @[RegFile.scala 66:20:@53566.4]
  wire  regs_274_io_reset; // @[RegFile.scala 66:20:@53566.4]
  wire [63:0] regs_274_io_out; // @[RegFile.scala 66:20:@53566.4]
  wire  regs_274_io_enable; // @[RegFile.scala 66:20:@53566.4]
  wire  regs_275_clock; // @[RegFile.scala 66:20:@53580.4]
  wire  regs_275_reset; // @[RegFile.scala 66:20:@53580.4]
  wire [63:0] regs_275_io_in; // @[RegFile.scala 66:20:@53580.4]
  wire  regs_275_io_reset; // @[RegFile.scala 66:20:@53580.4]
  wire [63:0] regs_275_io_out; // @[RegFile.scala 66:20:@53580.4]
  wire  regs_275_io_enable; // @[RegFile.scala 66:20:@53580.4]
  wire  regs_276_clock; // @[RegFile.scala 66:20:@53594.4]
  wire  regs_276_reset; // @[RegFile.scala 66:20:@53594.4]
  wire [63:0] regs_276_io_in; // @[RegFile.scala 66:20:@53594.4]
  wire  regs_276_io_reset; // @[RegFile.scala 66:20:@53594.4]
  wire [63:0] regs_276_io_out; // @[RegFile.scala 66:20:@53594.4]
  wire  regs_276_io_enable; // @[RegFile.scala 66:20:@53594.4]
  wire  regs_277_clock; // @[RegFile.scala 66:20:@53608.4]
  wire  regs_277_reset; // @[RegFile.scala 66:20:@53608.4]
  wire [63:0] regs_277_io_in; // @[RegFile.scala 66:20:@53608.4]
  wire  regs_277_io_reset; // @[RegFile.scala 66:20:@53608.4]
  wire [63:0] regs_277_io_out; // @[RegFile.scala 66:20:@53608.4]
  wire  regs_277_io_enable; // @[RegFile.scala 66:20:@53608.4]
  wire  regs_278_clock; // @[RegFile.scala 66:20:@53622.4]
  wire  regs_278_reset; // @[RegFile.scala 66:20:@53622.4]
  wire [63:0] regs_278_io_in; // @[RegFile.scala 66:20:@53622.4]
  wire  regs_278_io_reset; // @[RegFile.scala 66:20:@53622.4]
  wire [63:0] regs_278_io_out; // @[RegFile.scala 66:20:@53622.4]
  wire  regs_278_io_enable; // @[RegFile.scala 66:20:@53622.4]
  wire  regs_279_clock; // @[RegFile.scala 66:20:@53636.4]
  wire  regs_279_reset; // @[RegFile.scala 66:20:@53636.4]
  wire [63:0] regs_279_io_in; // @[RegFile.scala 66:20:@53636.4]
  wire  regs_279_io_reset; // @[RegFile.scala 66:20:@53636.4]
  wire [63:0] regs_279_io_out; // @[RegFile.scala 66:20:@53636.4]
  wire  regs_279_io_enable; // @[RegFile.scala 66:20:@53636.4]
  wire  regs_280_clock; // @[RegFile.scala 66:20:@53650.4]
  wire  regs_280_reset; // @[RegFile.scala 66:20:@53650.4]
  wire [63:0] regs_280_io_in; // @[RegFile.scala 66:20:@53650.4]
  wire  regs_280_io_reset; // @[RegFile.scala 66:20:@53650.4]
  wire [63:0] regs_280_io_out; // @[RegFile.scala 66:20:@53650.4]
  wire  regs_280_io_enable; // @[RegFile.scala 66:20:@53650.4]
  wire  regs_281_clock; // @[RegFile.scala 66:20:@53664.4]
  wire  regs_281_reset; // @[RegFile.scala 66:20:@53664.4]
  wire [63:0] regs_281_io_in; // @[RegFile.scala 66:20:@53664.4]
  wire  regs_281_io_reset; // @[RegFile.scala 66:20:@53664.4]
  wire [63:0] regs_281_io_out; // @[RegFile.scala 66:20:@53664.4]
  wire  regs_281_io_enable; // @[RegFile.scala 66:20:@53664.4]
  wire  regs_282_clock; // @[RegFile.scala 66:20:@53678.4]
  wire  regs_282_reset; // @[RegFile.scala 66:20:@53678.4]
  wire [63:0] regs_282_io_in; // @[RegFile.scala 66:20:@53678.4]
  wire  regs_282_io_reset; // @[RegFile.scala 66:20:@53678.4]
  wire [63:0] regs_282_io_out; // @[RegFile.scala 66:20:@53678.4]
  wire  regs_282_io_enable; // @[RegFile.scala 66:20:@53678.4]
  wire  regs_283_clock; // @[RegFile.scala 66:20:@53692.4]
  wire  regs_283_reset; // @[RegFile.scala 66:20:@53692.4]
  wire [63:0] regs_283_io_in; // @[RegFile.scala 66:20:@53692.4]
  wire  regs_283_io_reset; // @[RegFile.scala 66:20:@53692.4]
  wire [63:0] regs_283_io_out; // @[RegFile.scala 66:20:@53692.4]
  wire  regs_283_io_enable; // @[RegFile.scala 66:20:@53692.4]
  wire  regs_284_clock; // @[RegFile.scala 66:20:@53706.4]
  wire  regs_284_reset; // @[RegFile.scala 66:20:@53706.4]
  wire [63:0] regs_284_io_in; // @[RegFile.scala 66:20:@53706.4]
  wire  regs_284_io_reset; // @[RegFile.scala 66:20:@53706.4]
  wire [63:0] regs_284_io_out; // @[RegFile.scala 66:20:@53706.4]
  wire  regs_284_io_enable; // @[RegFile.scala 66:20:@53706.4]
  wire  regs_285_clock; // @[RegFile.scala 66:20:@53720.4]
  wire  regs_285_reset; // @[RegFile.scala 66:20:@53720.4]
  wire [63:0] regs_285_io_in; // @[RegFile.scala 66:20:@53720.4]
  wire  regs_285_io_reset; // @[RegFile.scala 66:20:@53720.4]
  wire [63:0] regs_285_io_out; // @[RegFile.scala 66:20:@53720.4]
  wire  regs_285_io_enable; // @[RegFile.scala 66:20:@53720.4]
  wire  regs_286_clock; // @[RegFile.scala 66:20:@53734.4]
  wire  regs_286_reset; // @[RegFile.scala 66:20:@53734.4]
  wire [63:0] regs_286_io_in; // @[RegFile.scala 66:20:@53734.4]
  wire  regs_286_io_reset; // @[RegFile.scala 66:20:@53734.4]
  wire [63:0] regs_286_io_out; // @[RegFile.scala 66:20:@53734.4]
  wire  regs_286_io_enable; // @[RegFile.scala 66:20:@53734.4]
  wire  regs_287_clock; // @[RegFile.scala 66:20:@53748.4]
  wire  regs_287_reset; // @[RegFile.scala 66:20:@53748.4]
  wire [63:0] regs_287_io_in; // @[RegFile.scala 66:20:@53748.4]
  wire  regs_287_io_reset; // @[RegFile.scala 66:20:@53748.4]
  wire [63:0] regs_287_io_out; // @[RegFile.scala 66:20:@53748.4]
  wire  regs_287_io_enable; // @[RegFile.scala 66:20:@53748.4]
  wire  regs_288_clock; // @[RegFile.scala 66:20:@53762.4]
  wire  regs_288_reset; // @[RegFile.scala 66:20:@53762.4]
  wire [63:0] regs_288_io_in; // @[RegFile.scala 66:20:@53762.4]
  wire  regs_288_io_reset; // @[RegFile.scala 66:20:@53762.4]
  wire [63:0] regs_288_io_out; // @[RegFile.scala 66:20:@53762.4]
  wire  regs_288_io_enable; // @[RegFile.scala 66:20:@53762.4]
  wire  regs_289_clock; // @[RegFile.scala 66:20:@53776.4]
  wire  regs_289_reset; // @[RegFile.scala 66:20:@53776.4]
  wire [63:0] regs_289_io_in; // @[RegFile.scala 66:20:@53776.4]
  wire  regs_289_io_reset; // @[RegFile.scala 66:20:@53776.4]
  wire [63:0] regs_289_io_out; // @[RegFile.scala 66:20:@53776.4]
  wire  regs_289_io_enable; // @[RegFile.scala 66:20:@53776.4]
  wire  regs_290_clock; // @[RegFile.scala 66:20:@53790.4]
  wire  regs_290_reset; // @[RegFile.scala 66:20:@53790.4]
  wire [63:0] regs_290_io_in; // @[RegFile.scala 66:20:@53790.4]
  wire  regs_290_io_reset; // @[RegFile.scala 66:20:@53790.4]
  wire [63:0] regs_290_io_out; // @[RegFile.scala 66:20:@53790.4]
  wire  regs_290_io_enable; // @[RegFile.scala 66:20:@53790.4]
  wire  regs_291_clock; // @[RegFile.scala 66:20:@53804.4]
  wire  regs_291_reset; // @[RegFile.scala 66:20:@53804.4]
  wire [63:0] regs_291_io_in; // @[RegFile.scala 66:20:@53804.4]
  wire  regs_291_io_reset; // @[RegFile.scala 66:20:@53804.4]
  wire [63:0] regs_291_io_out; // @[RegFile.scala 66:20:@53804.4]
  wire  regs_291_io_enable; // @[RegFile.scala 66:20:@53804.4]
  wire  regs_292_clock; // @[RegFile.scala 66:20:@53818.4]
  wire  regs_292_reset; // @[RegFile.scala 66:20:@53818.4]
  wire [63:0] regs_292_io_in; // @[RegFile.scala 66:20:@53818.4]
  wire  regs_292_io_reset; // @[RegFile.scala 66:20:@53818.4]
  wire [63:0] regs_292_io_out; // @[RegFile.scala 66:20:@53818.4]
  wire  regs_292_io_enable; // @[RegFile.scala 66:20:@53818.4]
  wire  regs_293_clock; // @[RegFile.scala 66:20:@53832.4]
  wire  regs_293_reset; // @[RegFile.scala 66:20:@53832.4]
  wire [63:0] regs_293_io_in; // @[RegFile.scala 66:20:@53832.4]
  wire  regs_293_io_reset; // @[RegFile.scala 66:20:@53832.4]
  wire [63:0] regs_293_io_out; // @[RegFile.scala 66:20:@53832.4]
  wire  regs_293_io_enable; // @[RegFile.scala 66:20:@53832.4]
  wire  regs_294_clock; // @[RegFile.scala 66:20:@53846.4]
  wire  regs_294_reset; // @[RegFile.scala 66:20:@53846.4]
  wire [63:0] regs_294_io_in; // @[RegFile.scala 66:20:@53846.4]
  wire  regs_294_io_reset; // @[RegFile.scala 66:20:@53846.4]
  wire [63:0] regs_294_io_out; // @[RegFile.scala 66:20:@53846.4]
  wire  regs_294_io_enable; // @[RegFile.scala 66:20:@53846.4]
  wire  regs_295_clock; // @[RegFile.scala 66:20:@53860.4]
  wire  regs_295_reset; // @[RegFile.scala 66:20:@53860.4]
  wire [63:0] regs_295_io_in; // @[RegFile.scala 66:20:@53860.4]
  wire  regs_295_io_reset; // @[RegFile.scala 66:20:@53860.4]
  wire [63:0] regs_295_io_out; // @[RegFile.scala 66:20:@53860.4]
  wire  regs_295_io_enable; // @[RegFile.scala 66:20:@53860.4]
  wire  regs_296_clock; // @[RegFile.scala 66:20:@53874.4]
  wire  regs_296_reset; // @[RegFile.scala 66:20:@53874.4]
  wire [63:0] regs_296_io_in; // @[RegFile.scala 66:20:@53874.4]
  wire  regs_296_io_reset; // @[RegFile.scala 66:20:@53874.4]
  wire [63:0] regs_296_io_out; // @[RegFile.scala 66:20:@53874.4]
  wire  regs_296_io_enable; // @[RegFile.scala 66:20:@53874.4]
  wire  regs_297_clock; // @[RegFile.scala 66:20:@53888.4]
  wire  regs_297_reset; // @[RegFile.scala 66:20:@53888.4]
  wire [63:0] regs_297_io_in; // @[RegFile.scala 66:20:@53888.4]
  wire  regs_297_io_reset; // @[RegFile.scala 66:20:@53888.4]
  wire [63:0] regs_297_io_out; // @[RegFile.scala 66:20:@53888.4]
  wire  regs_297_io_enable; // @[RegFile.scala 66:20:@53888.4]
  wire  regs_298_clock; // @[RegFile.scala 66:20:@53902.4]
  wire  regs_298_reset; // @[RegFile.scala 66:20:@53902.4]
  wire [63:0] regs_298_io_in; // @[RegFile.scala 66:20:@53902.4]
  wire  regs_298_io_reset; // @[RegFile.scala 66:20:@53902.4]
  wire [63:0] regs_298_io_out; // @[RegFile.scala 66:20:@53902.4]
  wire  regs_298_io_enable; // @[RegFile.scala 66:20:@53902.4]
  wire  regs_299_clock; // @[RegFile.scala 66:20:@53916.4]
  wire  regs_299_reset; // @[RegFile.scala 66:20:@53916.4]
  wire [63:0] regs_299_io_in; // @[RegFile.scala 66:20:@53916.4]
  wire  regs_299_io_reset; // @[RegFile.scala 66:20:@53916.4]
  wire [63:0] regs_299_io_out; // @[RegFile.scala 66:20:@53916.4]
  wire  regs_299_io_enable; // @[RegFile.scala 66:20:@53916.4]
  wire  regs_300_clock; // @[RegFile.scala 66:20:@53930.4]
  wire  regs_300_reset; // @[RegFile.scala 66:20:@53930.4]
  wire [63:0] regs_300_io_in; // @[RegFile.scala 66:20:@53930.4]
  wire  regs_300_io_reset; // @[RegFile.scala 66:20:@53930.4]
  wire [63:0] regs_300_io_out; // @[RegFile.scala 66:20:@53930.4]
  wire  regs_300_io_enable; // @[RegFile.scala 66:20:@53930.4]
  wire  regs_301_clock; // @[RegFile.scala 66:20:@53944.4]
  wire  regs_301_reset; // @[RegFile.scala 66:20:@53944.4]
  wire [63:0] regs_301_io_in; // @[RegFile.scala 66:20:@53944.4]
  wire  regs_301_io_reset; // @[RegFile.scala 66:20:@53944.4]
  wire [63:0] regs_301_io_out; // @[RegFile.scala 66:20:@53944.4]
  wire  regs_301_io_enable; // @[RegFile.scala 66:20:@53944.4]
  wire  regs_302_clock; // @[RegFile.scala 66:20:@53958.4]
  wire  regs_302_reset; // @[RegFile.scala 66:20:@53958.4]
  wire [63:0] regs_302_io_in; // @[RegFile.scala 66:20:@53958.4]
  wire  regs_302_io_reset; // @[RegFile.scala 66:20:@53958.4]
  wire [63:0] regs_302_io_out; // @[RegFile.scala 66:20:@53958.4]
  wire  regs_302_io_enable; // @[RegFile.scala 66:20:@53958.4]
  wire  regs_303_clock; // @[RegFile.scala 66:20:@53972.4]
  wire  regs_303_reset; // @[RegFile.scala 66:20:@53972.4]
  wire [63:0] regs_303_io_in; // @[RegFile.scala 66:20:@53972.4]
  wire  regs_303_io_reset; // @[RegFile.scala 66:20:@53972.4]
  wire [63:0] regs_303_io_out; // @[RegFile.scala 66:20:@53972.4]
  wire  regs_303_io_enable; // @[RegFile.scala 66:20:@53972.4]
  wire  regs_304_clock; // @[RegFile.scala 66:20:@53986.4]
  wire  regs_304_reset; // @[RegFile.scala 66:20:@53986.4]
  wire [63:0] regs_304_io_in; // @[RegFile.scala 66:20:@53986.4]
  wire  regs_304_io_reset; // @[RegFile.scala 66:20:@53986.4]
  wire [63:0] regs_304_io_out; // @[RegFile.scala 66:20:@53986.4]
  wire  regs_304_io_enable; // @[RegFile.scala 66:20:@53986.4]
  wire  regs_305_clock; // @[RegFile.scala 66:20:@54000.4]
  wire  regs_305_reset; // @[RegFile.scala 66:20:@54000.4]
  wire [63:0] regs_305_io_in; // @[RegFile.scala 66:20:@54000.4]
  wire  regs_305_io_reset; // @[RegFile.scala 66:20:@54000.4]
  wire [63:0] regs_305_io_out; // @[RegFile.scala 66:20:@54000.4]
  wire  regs_305_io_enable; // @[RegFile.scala 66:20:@54000.4]
  wire  regs_306_clock; // @[RegFile.scala 66:20:@54014.4]
  wire  regs_306_reset; // @[RegFile.scala 66:20:@54014.4]
  wire [63:0] regs_306_io_in; // @[RegFile.scala 66:20:@54014.4]
  wire  regs_306_io_reset; // @[RegFile.scala 66:20:@54014.4]
  wire [63:0] regs_306_io_out; // @[RegFile.scala 66:20:@54014.4]
  wire  regs_306_io_enable; // @[RegFile.scala 66:20:@54014.4]
  wire  regs_307_clock; // @[RegFile.scala 66:20:@54028.4]
  wire  regs_307_reset; // @[RegFile.scala 66:20:@54028.4]
  wire [63:0] regs_307_io_in; // @[RegFile.scala 66:20:@54028.4]
  wire  regs_307_io_reset; // @[RegFile.scala 66:20:@54028.4]
  wire [63:0] regs_307_io_out; // @[RegFile.scala 66:20:@54028.4]
  wire  regs_307_io_enable; // @[RegFile.scala 66:20:@54028.4]
  wire  regs_308_clock; // @[RegFile.scala 66:20:@54042.4]
  wire  regs_308_reset; // @[RegFile.scala 66:20:@54042.4]
  wire [63:0] regs_308_io_in; // @[RegFile.scala 66:20:@54042.4]
  wire  regs_308_io_reset; // @[RegFile.scala 66:20:@54042.4]
  wire [63:0] regs_308_io_out; // @[RegFile.scala 66:20:@54042.4]
  wire  regs_308_io_enable; // @[RegFile.scala 66:20:@54042.4]
  wire  regs_309_clock; // @[RegFile.scala 66:20:@54056.4]
  wire  regs_309_reset; // @[RegFile.scala 66:20:@54056.4]
  wire [63:0] regs_309_io_in; // @[RegFile.scala 66:20:@54056.4]
  wire  regs_309_io_reset; // @[RegFile.scala 66:20:@54056.4]
  wire [63:0] regs_309_io_out; // @[RegFile.scala 66:20:@54056.4]
  wire  regs_309_io_enable; // @[RegFile.scala 66:20:@54056.4]
  wire  regs_310_clock; // @[RegFile.scala 66:20:@54070.4]
  wire  regs_310_reset; // @[RegFile.scala 66:20:@54070.4]
  wire [63:0] regs_310_io_in; // @[RegFile.scala 66:20:@54070.4]
  wire  regs_310_io_reset; // @[RegFile.scala 66:20:@54070.4]
  wire [63:0] regs_310_io_out; // @[RegFile.scala 66:20:@54070.4]
  wire  regs_310_io_enable; // @[RegFile.scala 66:20:@54070.4]
  wire  regs_311_clock; // @[RegFile.scala 66:20:@54084.4]
  wire  regs_311_reset; // @[RegFile.scala 66:20:@54084.4]
  wire [63:0] regs_311_io_in; // @[RegFile.scala 66:20:@54084.4]
  wire  regs_311_io_reset; // @[RegFile.scala 66:20:@54084.4]
  wire [63:0] regs_311_io_out; // @[RegFile.scala 66:20:@54084.4]
  wire  regs_311_io_enable; // @[RegFile.scala 66:20:@54084.4]
  wire  regs_312_clock; // @[RegFile.scala 66:20:@54098.4]
  wire  regs_312_reset; // @[RegFile.scala 66:20:@54098.4]
  wire [63:0] regs_312_io_in; // @[RegFile.scala 66:20:@54098.4]
  wire  regs_312_io_reset; // @[RegFile.scala 66:20:@54098.4]
  wire [63:0] regs_312_io_out; // @[RegFile.scala 66:20:@54098.4]
  wire  regs_312_io_enable; // @[RegFile.scala 66:20:@54098.4]
  wire  regs_313_clock; // @[RegFile.scala 66:20:@54112.4]
  wire  regs_313_reset; // @[RegFile.scala 66:20:@54112.4]
  wire [63:0] regs_313_io_in; // @[RegFile.scala 66:20:@54112.4]
  wire  regs_313_io_reset; // @[RegFile.scala 66:20:@54112.4]
  wire [63:0] regs_313_io_out; // @[RegFile.scala 66:20:@54112.4]
  wire  regs_313_io_enable; // @[RegFile.scala 66:20:@54112.4]
  wire  regs_314_clock; // @[RegFile.scala 66:20:@54126.4]
  wire  regs_314_reset; // @[RegFile.scala 66:20:@54126.4]
  wire [63:0] regs_314_io_in; // @[RegFile.scala 66:20:@54126.4]
  wire  regs_314_io_reset; // @[RegFile.scala 66:20:@54126.4]
  wire [63:0] regs_314_io_out; // @[RegFile.scala 66:20:@54126.4]
  wire  regs_314_io_enable; // @[RegFile.scala 66:20:@54126.4]
  wire  regs_315_clock; // @[RegFile.scala 66:20:@54140.4]
  wire  regs_315_reset; // @[RegFile.scala 66:20:@54140.4]
  wire [63:0] regs_315_io_in; // @[RegFile.scala 66:20:@54140.4]
  wire  regs_315_io_reset; // @[RegFile.scala 66:20:@54140.4]
  wire [63:0] regs_315_io_out; // @[RegFile.scala 66:20:@54140.4]
  wire  regs_315_io_enable; // @[RegFile.scala 66:20:@54140.4]
  wire  regs_316_clock; // @[RegFile.scala 66:20:@54154.4]
  wire  regs_316_reset; // @[RegFile.scala 66:20:@54154.4]
  wire [63:0] regs_316_io_in; // @[RegFile.scala 66:20:@54154.4]
  wire  regs_316_io_reset; // @[RegFile.scala 66:20:@54154.4]
  wire [63:0] regs_316_io_out; // @[RegFile.scala 66:20:@54154.4]
  wire  regs_316_io_enable; // @[RegFile.scala 66:20:@54154.4]
  wire  regs_317_clock; // @[RegFile.scala 66:20:@54168.4]
  wire  regs_317_reset; // @[RegFile.scala 66:20:@54168.4]
  wire [63:0] regs_317_io_in; // @[RegFile.scala 66:20:@54168.4]
  wire  regs_317_io_reset; // @[RegFile.scala 66:20:@54168.4]
  wire [63:0] regs_317_io_out; // @[RegFile.scala 66:20:@54168.4]
  wire  regs_317_io_enable; // @[RegFile.scala 66:20:@54168.4]
  wire  regs_318_clock; // @[RegFile.scala 66:20:@54182.4]
  wire  regs_318_reset; // @[RegFile.scala 66:20:@54182.4]
  wire [63:0] regs_318_io_in; // @[RegFile.scala 66:20:@54182.4]
  wire  regs_318_io_reset; // @[RegFile.scala 66:20:@54182.4]
  wire [63:0] regs_318_io_out; // @[RegFile.scala 66:20:@54182.4]
  wire  regs_318_io_enable; // @[RegFile.scala 66:20:@54182.4]
  wire  regs_319_clock; // @[RegFile.scala 66:20:@54196.4]
  wire  regs_319_reset; // @[RegFile.scala 66:20:@54196.4]
  wire [63:0] regs_319_io_in; // @[RegFile.scala 66:20:@54196.4]
  wire  regs_319_io_reset; // @[RegFile.scala 66:20:@54196.4]
  wire [63:0] regs_319_io_out; // @[RegFile.scala 66:20:@54196.4]
  wire  regs_319_io_enable; // @[RegFile.scala 66:20:@54196.4]
  wire  regs_320_clock; // @[RegFile.scala 66:20:@54210.4]
  wire  regs_320_reset; // @[RegFile.scala 66:20:@54210.4]
  wire [63:0] regs_320_io_in; // @[RegFile.scala 66:20:@54210.4]
  wire  regs_320_io_reset; // @[RegFile.scala 66:20:@54210.4]
  wire [63:0] regs_320_io_out; // @[RegFile.scala 66:20:@54210.4]
  wire  regs_320_io_enable; // @[RegFile.scala 66:20:@54210.4]
  wire  regs_321_clock; // @[RegFile.scala 66:20:@54224.4]
  wire  regs_321_reset; // @[RegFile.scala 66:20:@54224.4]
  wire [63:0] regs_321_io_in; // @[RegFile.scala 66:20:@54224.4]
  wire  regs_321_io_reset; // @[RegFile.scala 66:20:@54224.4]
  wire [63:0] regs_321_io_out; // @[RegFile.scala 66:20:@54224.4]
  wire  regs_321_io_enable; // @[RegFile.scala 66:20:@54224.4]
  wire  regs_322_clock; // @[RegFile.scala 66:20:@54238.4]
  wire  regs_322_reset; // @[RegFile.scala 66:20:@54238.4]
  wire [63:0] regs_322_io_in; // @[RegFile.scala 66:20:@54238.4]
  wire  regs_322_io_reset; // @[RegFile.scala 66:20:@54238.4]
  wire [63:0] regs_322_io_out; // @[RegFile.scala 66:20:@54238.4]
  wire  regs_322_io_enable; // @[RegFile.scala 66:20:@54238.4]
  wire  regs_323_clock; // @[RegFile.scala 66:20:@54252.4]
  wire  regs_323_reset; // @[RegFile.scala 66:20:@54252.4]
  wire [63:0] regs_323_io_in; // @[RegFile.scala 66:20:@54252.4]
  wire  regs_323_io_reset; // @[RegFile.scala 66:20:@54252.4]
  wire [63:0] regs_323_io_out; // @[RegFile.scala 66:20:@54252.4]
  wire  regs_323_io_enable; // @[RegFile.scala 66:20:@54252.4]
  wire  regs_324_clock; // @[RegFile.scala 66:20:@54266.4]
  wire  regs_324_reset; // @[RegFile.scala 66:20:@54266.4]
  wire [63:0] regs_324_io_in; // @[RegFile.scala 66:20:@54266.4]
  wire  regs_324_io_reset; // @[RegFile.scala 66:20:@54266.4]
  wire [63:0] regs_324_io_out; // @[RegFile.scala 66:20:@54266.4]
  wire  regs_324_io_enable; // @[RegFile.scala 66:20:@54266.4]
  wire  regs_325_clock; // @[RegFile.scala 66:20:@54280.4]
  wire  regs_325_reset; // @[RegFile.scala 66:20:@54280.4]
  wire [63:0] regs_325_io_in; // @[RegFile.scala 66:20:@54280.4]
  wire  regs_325_io_reset; // @[RegFile.scala 66:20:@54280.4]
  wire [63:0] regs_325_io_out; // @[RegFile.scala 66:20:@54280.4]
  wire  regs_325_io_enable; // @[RegFile.scala 66:20:@54280.4]
  wire  regs_326_clock; // @[RegFile.scala 66:20:@54294.4]
  wire  regs_326_reset; // @[RegFile.scala 66:20:@54294.4]
  wire [63:0] regs_326_io_in; // @[RegFile.scala 66:20:@54294.4]
  wire  regs_326_io_reset; // @[RegFile.scala 66:20:@54294.4]
  wire [63:0] regs_326_io_out; // @[RegFile.scala 66:20:@54294.4]
  wire  regs_326_io_enable; // @[RegFile.scala 66:20:@54294.4]
  wire  regs_327_clock; // @[RegFile.scala 66:20:@54308.4]
  wire  regs_327_reset; // @[RegFile.scala 66:20:@54308.4]
  wire [63:0] regs_327_io_in; // @[RegFile.scala 66:20:@54308.4]
  wire  regs_327_io_reset; // @[RegFile.scala 66:20:@54308.4]
  wire [63:0] regs_327_io_out; // @[RegFile.scala 66:20:@54308.4]
  wire  regs_327_io_enable; // @[RegFile.scala 66:20:@54308.4]
  wire  regs_328_clock; // @[RegFile.scala 66:20:@54322.4]
  wire  regs_328_reset; // @[RegFile.scala 66:20:@54322.4]
  wire [63:0] regs_328_io_in; // @[RegFile.scala 66:20:@54322.4]
  wire  regs_328_io_reset; // @[RegFile.scala 66:20:@54322.4]
  wire [63:0] regs_328_io_out; // @[RegFile.scala 66:20:@54322.4]
  wire  regs_328_io_enable; // @[RegFile.scala 66:20:@54322.4]
  wire  regs_329_clock; // @[RegFile.scala 66:20:@54336.4]
  wire  regs_329_reset; // @[RegFile.scala 66:20:@54336.4]
  wire [63:0] regs_329_io_in; // @[RegFile.scala 66:20:@54336.4]
  wire  regs_329_io_reset; // @[RegFile.scala 66:20:@54336.4]
  wire [63:0] regs_329_io_out; // @[RegFile.scala 66:20:@54336.4]
  wire  regs_329_io_enable; // @[RegFile.scala 66:20:@54336.4]
  wire  regs_330_clock; // @[RegFile.scala 66:20:@54350.4]
  wire  regs_330_reset; // @[RegFile.scala 66:20:@54350.4]
  wire [63:0] regs_330_io_in; // @[RegFile.scala 66:20:@54350.4]
  wire  regs_330_io_reset; // @[RegFile.scala 66:20:@54350.4]
  wire [63:0] regs_330_io_out; // @[RegFile.scala 66:20:@54350.4]
  wire  regs_330_io_enable; // @[RegFile.scala 66:20:@54350.4]
  wire  regs_331_clock; // @[RegFile.scala 66:20:@54364.4]
  wire  regs_331_reset; // @[RegFile.scala 66:20:@54364.4]
  wire [63:0] regs_331_io_in; // @[RegFile.scala 66:20:@54364.4]
  wire  regs_331_io_reset; // @[RegFile.scala 66:20:@54364.4]
  wire [63:0] regs_331_io_out; // @[RegFile.scala 66:20:@54364.4]
  wire  regs_331_io_enable; // @[RegFile.scala 66:20:@54364.4]
  wire  regs_332_clock; // @[RegFile.scala 66:20:@54378.4]
  wire  regs_332_reset; // @[RegFile.scala 66:20:@54378.4]
  wire [63:0] regs_332_io_in; // @[RegFile.scala 66:20:@54378.4]
  wire  regs_332_io_reset; // @[RegFile.scala 66:20:@54378.4]
  wire [63:0] regs_332_io_out; // @[RegFile.scala 66:20:@54378.4]
  wire  regs_332_io_enable; // @[RegFile.scala 66:20:@54378.4]
  wire  regs_333_clock; // @[RegFile.scala 66:20:@54392.4]
  wire  regs_333_reset; // @[RegFile.scala 66:20:@54392.4]
  wire [63:0] regs_333_io_in; // @[RegFile.scala 66:20:@54392.4]
  wire  regs_333_io_reset; // @[RegFile.scala 66:20:@54392.4]
  wire [63:0] regs_333_io_out; // @[RegFile.scala 66:20:@54392.4]
  wire  regs_333_io_enable; // @[RegFile.scala 66:20:@54392.4]
  wire  regs_334_clock; // @[RegFile.scala 66:20:@54406.4]
  wire  regs_334_reset; // @[RegFile.scala 66:20:@54406.4]
  wire [63:0] regs_334_io_in; // @[RegFile.scala 66:20:@54406.4]
  wire  regs_334_io_reset; // @[RegFile.scala 66:20:@54406.4]
  wire [63:0] regs_334_io_out; // @[RegFile.scala 66:20:@54406.4]
  wire  regs_334_io_enable; // @[RegFile.scala 66:20:@54406.4]
  wire  regs_335_clock; // @[RegFile.scala 66:20:@54420.4]
  wire  regs_335_reset; // @[RegFile.scala 66:20:@54420.4]
  wire [63:0] regs_335_io_in; // @[RegFile.scala 66:20:@54420.4]
  wire  regs_335_io_reset; // @[RegFile.scala 66:20:@54420.4]
  wire [63:0] regs_335_io_out; // @[RegFile.scala 66:20:@54420.4]
  wire  regs_335_io_enable; // @[RegFile.scala 66:20:@54420.4]
  wire  regs_336_clock; // @[RegFile.scala 66:20:@54434.4]
  wire  regs_336_reset; // @[RegFile.scala 66:20:@54434.4]
  wire [63:0] regs_336_io_in; // @[RegFile.scala 66:20:@54434.4]
  wire  regs_336_io_reset; // @[RegFile.scala 66:20:@54434.4]
  wire [63:0] regs_336_io_out; // @[RegFile.scala 66:20:@54434.4]
  wire  regs_336_io_enable; // @[RegFile.scala 66:20:@54434.4]
  wire  regs_337_clock; // @[RegFile.scala 66:20:@54448.4]
  wire  regs_337_reset; // @[RegFile.scala 66:20:@54448.4]
  wire [63:0] regs_337_io_in; // @[RegFile.scala 66:20:@54448.4]
  wire  regs_337_io_reset; // @[RegFile.scala 66:20:@54448.4]
  wire [63:0] regs_337_io_out; // @[RegFile.scala 66:20:@54448.4]
  wire  regs_337_io_enable; // @[RegFile.scala 66:20:@54448.4]
  wire  regs_338_clock; // @[RegFile.scala 66:20:@54462.4]
  wire  regs_338_reset; // @[RegFile.scala 66:20:@54462.4]
  wire [63:0] regs_338_io_in; // @[RegFile.scala 66:20:@54462.4]
  wire  regs_338_io_reset; // @[RegFile.scala 66:20:@54462.4]
  wire [63:0] regs_338_io_out; // @[RegFile.scala 66:20:@54462.4]
  wire  regs_338_io_enable; // @[RegFile.scala 66:20:@54462.4]
  wire  regs_339_clock; // @[RegFile.scala 66:20:@54476.4]
  wire  regs_339_reset; // @[RegFile.scala 66:20:@54476.4]
  wire [63:0] regs_339_io_in; // @[RegFile.scala 66:20:@54476.4]
  wire  regs_339_io_reset; // @[RegFile.scala 66:20:@54476.4]
  wire [63:0] regs_339_io_out; // @[RegFile.scala 66:20:@54476.4]
  wire  regs_339_io_enable; // @[RegFile.scala 66:20:@54476.4]
  wire  regs_340_clock; // @[RegFile.scala 66:20:@54490.4]
  wire  regs_340_reset; // @[RegFile.scala 66:20:@54490.4]
  wire [63:0] regs_340_io_in; // @[RegFile.scala 66:20:@54490.4]
  wire  regs_340_io_reset; // @[RegFile.scala 66:20:@54490.4]
  wire [63:0] regs_340_io_out; // @[RegFile.scala 66:20:@54490.4]
  wire  regs_340_io_enable; // @[RegFile.scala 66:20:@54490.4]
  wire  regs_341_clock; // @[RegFile.scala 66:20:@54504.4]
  wire  regs_341_reset; // @[RegFile.scala 66:20:@54504.4]
  wire [63:0] regs_341_io_in; // @[RegFile.scala 66:20:@54504.4]
  wire  regs_341_io_reset; // @[RegFile.scala 66:20:@54504.4]
  wire [63:0] regs_341_io_out; // @[RegFile.scala 66:20:@54504.4]
  wire  regs_341_io_enable; // @[RegFile.scala 66:20:@54504.4]
  wire  regs_342_clock; // @[RegFile.scala 66:20:@54518.4]
  wire  regs_342_reset; // @[RegFile.scala 66:20:@54518.4]
  wire [63:0] regs_342_io_in; // @[RegFile.scala 66:20:@54518.4]
  wire  regs_342_io_reset; // @[RegFile.scala 66:20:@54518.4]
  wire [63:0] regs_342_io_out; // @[RegFile.scala 66:20:@54518.4]
  wire  regs_342_io_enable; // @[RegFile.scala 66:20:@54518.4]
  wire  regs_343_clock; // @[RegFile.scala 66:20:@54532.4]
  wire  regs_343_reset; // @[RegFile.scala 66:20:@54532.4]
  wire [63:0] regs_343_io_in; // @[RegFile.scala 66:20:@54532.4]
  wire  regs_343_io_reset; // @[RegFile.scala 66:20:@54532.4]
  wire [63:0] regs_343_io_out; // @[RegFile.scala 66:20:@54532.4]
  wire  regs_343_io_enable; // @[RegFile.scala 66:20:@54532.4]
  wire  regs_344_clock; // @[RegFile.scala 66:20:@54546.4]
  wire  regs_344_reset; // @[RegFile.scala 66:20:@54546.4]
  wire [63:0] regs_344_io_in; // @[RegFile.scala 66:20:@54546.4]
  wire  regs_344_io_reset; // @[RegFile.scala 66:20:@54546.4]
  wire [63:0] regs_344_io_out; // @[RegFile.scala 66:20:@54546.4]
  wire  regs_344_io_enable; // @[RegFile.scala 66:20:@54546.4]
  wire  regs_345_clock; // @[RegFile.scala 66:20:@54560.4]
  wire  regs_345_reset; // @[RegFile.scala 66:20:@54560.4]
  wire [63:0] regs_345_io_in; // @[RegFile.scala 66:20:@54560.4]
  wire  regs_345_io_reset; // @[RegFile.scala 66:20:@54560.4]
  wire [63:0] regs_345_io_out; // @[RegFile.scala 66:20:@54560.4]
  wire  regs_345_io_enable; // @[RegFile.scala 66:20:@54560.4]
  wire  regs_346_clock; // @[RegFile.scala 66:20:@54574.4]
  wire  regs_346_reset; // @[RegFile.scala 66:20:@54574.4]
  wire [63:0] regs_346_io_in; // @[RegFile.scala 66:20:@54574.4]
  wire  regs_346_io_reset; // @[RegFile.scala 66:20:@54574.4]
  wire [63:0] regs_346_io_out; // @[RegFile.scala 66:20:@54574.4]
  wire  regs_346_io_enable; // @[RegFile.scala 66:20:@54574.4]
  wire  regs_347_clock; // @[RegFile.scala 66:20:@54588.4]
  wire  regs_347_reset; // @[RegFile.scala 66:20:@54588.4]
  wire [63:0] regs_347_io_in; // @[RegFile.scala 66:20:@54588.4]
  wire  regs_347_io_reset; // @[RegFile.scala 66:20:@54588.4]
  wire [63:0] regs_347_io_out; // @[RegFile.scala 66:20:@54588.4]
  wire  regs_347_io_enable; // @[RegFile.scala 66:20:@54588.4]
  wire  regs_348_clock; // @[RegFile.scala 66:20:@54602.4]
  wire  regs_348_reset; // @[RegFile.scala 66:20:@54602.4]
  wire [63:0] regs_348_io_in; // @[RegFile.scala 66:20:@54602.4]
  wire  regs_348_io_reset; // @[RegFile.scala 66:20:@54602.4]
  wire [63:0] regs_348_io_out; // @[RegFile.scala 66:20:@54602.4]
  wire  regs_348_io_enable; // @[RegFile.scala 66:20:@54602.4]
  wire  regs_349_clock; // @[RegFile.scala 66:20:@54616.4]
  wire  regs_349_reset; // @[RegFile.scala 66:20:@54616.4]
  wire [63:0] regs_349_io_in; // @[RegFile.scala 66:20:@54616.4]
  wire  regs_349_io_reset; // @[RegFile.scala 66:20:@54616.4]
  wire [63:0] regs_349_io_out; // @[RegFile.scala 66:20:@54616.4]
  wire  regs_349_io_enable; // @[RegFile.scala 66:20:@54616.4]
  wire  regs_350_clock; // @[RegFile.scala 66:20:@54630.4]
  wire  regs_350_reset; // @[RegFile.scala 66:20:@54630.4]
  wire [63:0] regs_350_io_in; // @[RegFile.scala 66:20:@54630.4]
  wire  regs_350_io_reset; // @[RegFile.scala 66:20:@54630.4]
  wire [63:0] regs_350_io_out; // @[RegFile.scala 66:20:@54630.4]
  wire  regs_350_io_enable; // @[RegFile.scala 66:20:@54630.4]
  wire  regs_351_clock; // @[RegFile.scala 66:20:@54644.4]
  wire  regs_351_reset; // @[RegFile.scala 66:20:@54644.4]
  wire [63:0] regs_351_io_in; // @[RegFile.scala 66:20:@54644.4]
  wire  regs_351_io_reset; // @[RegFile.scala 66:20:@54644.4]
  wire [63:0] regs_351_io_out; // @[RegFile.scala 66:20:@54644.4]
  wire  regs_351_io_enable; // @[RegFile.scala 66:20:@54644.4]
  wire  regs_352_clock; // @[RegFile.scala 66:20:@54658.4]
  wire  regs_352_reset; // @[RegFile.scala 66:20:@54658.4]
  wire [63:0] regs_352_io_in; // @[RegFile.scala 66:20:@54658.4]
  wire  regs_352_io_reset; // @[RegFile.scala 66:20:@54658.4]
  wire [63:0] regs_352_io_out; // @[RegFile.scala 66:20:@54658.4]
  wire  regs_352_io_enable; // @[RegFile.scala 66:20:@54658.4]
  wire  regs_353_clock; // @[RegFile.scala 66:20:@54672.4]
  wire  regs_353_reset; // @[RegFile.scala 66:20:@54672.4]
  wire [63:0] regs_353_io_in; // @[RegFile.scala 66:20:@54672.4]
  wire  regs_353_io_reset; // @[RegFile.scala 66:20:@54672.4]
  wire [63:0] regs_353_io_out; // @[RegFile.scala 66:20:@54672.4]
  wire  regs_353_io_enable; // @[RegFile.scala 66:20:@54672.4]
  wire  regs_354_clock; // @[RegFile.scala 66:20:@54686.4]
  wire  regs_354_reset; // @[RegFile.scala 66:20:@54686.4]
  wire [63:0] regs_354_io_in; // @[RegFile.scala 66:20:@54686.4]
  wire  regs_354_io_reset; // @[RegFile.scala 66:20:@54686.4]
  wire [63:0] regs_354_io_out; // @[RegFile.scala 66:20:@54686.4]
  wire  regs_354_io_enable; // @[RegFile.scala 66:20:@54686.4]
  wire  regs_355_clock; // @[RegFile.scala 66:20:@54700.4]
  wire  regs_355_reset; // @[RegFile.scala 66:20:@54700.4]
  wire [63:0] regs_355_io_in; // @[RegFile.scala 66:20:@54700.4]
  wire  regs_355_io_reset; // @[RegFile.scala 66:20:@54700.4]
  wire [63:0] regs_355_io_out; // @[RegFile.scala 66:20:@54700.4]
  wire  regs_355_io_enable; // @[RegFile.scala 66:20:@54700.4]
  wire  regs_356_clock; // @[RegFile.scala 66:20:@54714.4]
  wire  regs_356_reset; // @[RegFile.scala 66:20:@54714.4]
  wire [63:0] regs_356_io_in; // @[RegFile.scala 66:20:@54714.4]
  wire  regs_356_io_reset; // @[RegFile.scala 66:20:@54714.4]
  wire [63:0] regs_356_io_out; // @[RegFile.scala 66:20:@54714.4]
  wire  regs_356_io_enable; // @[RegFile.scala 66:20:@54714.4]
  wire  regs_357_clock; // @[RegFile.scala 66:20:@54728.4]
  wire  regs_357_reset; // @[RegFile.scala 66:20:@54728.4]
  wire [63:0] regs_357_io_in; // @[RegFile.scala 66:20:@54728.4]
  wire  regs_357_io_reset; // @[RegFile.scala 66:20:@54728.4]
  wire [63:0] regs_357_io_out; // @[RegFile.scala 66:20:@54728.4]
  wire  regs_357_io_enable; // @[RegFile.scala 66:20:@54728.4]
  wire  regs_358_clock; // @[RegFile.scala 66:20:@54742.4]
  wire  regs_358_reset; // @[RegFile.scala 66:20:@54742.4]
  wire [63:0] regs_358_io_in; // @[RegFile.scala 66:20:@54742.4]
  wire  regs_358_io_reset; // @[RegFile.scala 66:20:@54742.4]
  wire [63:0] regs_358_io_out; // @[RegFile.scala 66:20:@54742.4]
  wire  regs_358_io_enable; // @[RegFile.scala 66:20:@54742.4]
  wire  regs_359_clock; // @[RegFile.scala 66:20:@54756.4]
  wire  regs_359_reset; // @[RegFile.scala 66:20:@54756.4]
  wire [63:0] regs_359_io_in; // @[RegFile.scala 66:20:@54756.4]
  wire  regs_359_io_reset; // @[RegFile.scala 66:20:@54756.4]
  wire [63:0] regs_359_io_out; // @[RegFile.scala 66:20:@54756.4]
  wire  regs_359_io_enable; // @[RegFile.scala 66:20:@54756.4]
  wire  regs_360_clock; // @[RegFile.scala 66:20:@54770.4]
  wire  regs_360_reset; // @[RegFile.scala 66:20:@54770.4]
  wire [63:0] regs_360_io_in; // @[RegFile.scala 66:20:@54770.4]
  wire  regs_360_io_reset; // @[RegFile.scala 66:20:@54770.4]
  wire [63:0] regs_360_io_out; // @[RegFile.scala 66:20:@54770.4]
  wire  regs_360_io_enable; // @[RegFile.scala 66:20:@54770.4]
  wire  regs_361_clock; // @[RegFile.scala 66:20:@54784.4]
  wire  regs_361_reset; // @[RegFile.scala 66:20:@54784.4]
  wire [63:0] regs_361_io_in; // @[RegFile.scala 66:20:@54784.4]
  wire  regs_361_io_reset; // @[RegFile.scala 66:20:@54784.4]
  wire [63:0] regs_361_io_out; // @[RegFile.scala 66:20:@54784.4]
  wire  regs_361_io_enable; // @[RegFile.scala 66:20:@54784.4]
  wire  regs_362_clock; // @[RegFile.scala 66:20:@54798.4]
  wire  regs_362_reset; // @[RegFile.scala 66:20:@54798.4]
  wire [63:0] regs_362_io_in; // @[RegFile.scala 66:20:@54798.4]
  wire  regs_362_io_reset; // @[RegFile.scala 66:20:@54798.4]
  wire [63:0] regs_362_io_out; // @[RegFile.scala 66:20:@54798.4]
  wire  regs_362_io_enable; // @[RegFile.scala 66:20:@54798.4]
  wire  regs_363_clock; // @[RegFile.scala 66:20:@54812.4]
  wire  regs_363_reset; // @[RegFile.scala 66:20:@54812.4]
  wire [63:0] regs_363_io_in; // @[RegFile.scala 66:20:@54812.4]
  wire  regs_363_io_reset; // @[RegFile.scala 66:20:@54812.4]
  wire [63:0] regs_363_io_out; // @[RegFile.scala 66:20:@54812.4]
  wire  regs_363_io_enable; // @[RegFile.scala 66:20:@54812.4]
  wire  regs_364_clock; // @[RegFile.scala 66:20:@54826.4]
  wire  regs_364_reset; // @[RegFile.scala 66:20:@54826.4]
  wire [63:0] regs_364_io_in; // @[RegFile.scala 66:20:@54826.4]
  wire  regs_364_io_reset; // @[RegFile.scala 66:20:@54826.4]
  wire [63:0] regs_364_io_out; // @[RegFile.scala 66:20:@54826.4]
  wire  regs_364_io_enable; // @[RegFile.scala 66:20:@54826.4]
  wire  regs_365_clock; // @[RegFile.scala 66:20:@54840.4]
  wire  regs_365_reset; // @[RegFile.scala 66:20:@54840.4]
  wire [63:0] regs_365_io_in; // @[RegFile.scala 66:20:@54840.4]
  wire  regs_365_io_reset; // @[RegFile.scala 66:20:@54840.4]
  wire [63:0] regs_365_io_out; // @[RegFile.scala 66:20:@54840.4]
  wire  regs_365_io_enable; // @[RegFile.scala 66:20:@54840.4]
  wire  regs_366_clock; // @[RegFile.scala 66:20:@54854.4]
  wire  regs_366_reset; // @[RegFile.scala 66:20:@54854.4]
  wire [63:0] regs_366_io_in; // @[RegFile.scala 66:20:@54854.4]
  wire  regs_366_io_reset; // @[RegFile.scala 66:20:@54854.4]
  wire [63:0] regs_366_io_out; // @[RegFile.scala 66:20:@54854.4]
  wire  regs_366_io_enable; // @[RegFile.scala 66:20:@54854.4]
  wire  regs_367_clock; // @[RegFile.scala 66:20:@54868.4]
  wire  regs_367_reset; // @[RegFile.scala 66:20:@54868.4]
  wire [63:0] regs_367_io_in; // @[RegFile.scala 66:20:@54868.4]
  wire  regs_367_io_reset; // @[RegFile.scala 66:20:@54868.4]
  wire [63:0] regs_367_io_out; // @[RegFile.scala 66:20:@54868.4]
  wire  regs_367_io_enable; // @[RegFile.scala 66:20:@54868.4]
  wire  regs_368_clock; // @[RegFile.scala 66:20:@54882.4]
  wire  regs_368_reset; // @[RegFile.scala 66:20:@54882.4]
  wire [63:0] regs_368_io_in; // @[RegFile.scala 66:20:@54882.4]
  wire  regs_368_io_reset; // @[RegFile.scala 66:20:@54882.4]
  wire [63:0] regs_368_io_out; // @[RegFile.scala 66:20:@54882.4]
  wire  regs_368_io_enable; // @[RegFile.scala 66:20:@54882.4]
  wire  regs_369_clock; // @[RegFile.scala 66:20:@54896.4]
  wire  regs_369_reset; // @[RegFile.scala 66:20:@54896.4]
  wire [63:0] regs_369_io_in; // @[RegFile.scala 66:20:@54896.4]
  wire  regs_369_io_reset; // @[RegFile.scala 66:20:@54896.4]
  wire [63:0] regs_369_io_out; // @[RegFile.scala 66:20:@54896.4]
  wire  regs_369_io_enable; // @[RegFile.scala 66:20:@54896.4]
  wire  regs_370_clock; // @[RegFile.scala 66:20:@54910.4]
  wire  regs_370_reset; // @[RegFile.scala 66:20:@54910.4]
  wire [63:0] regs_370_io_in; // @[RegFile.scala 66:20:@54910.4]
  wire  regs_370_io_reset; // @[RegFile.scala 66:20:@54910.4]
  wire [63:0] regs_370_io_out; // @[RegFile.scala 66:20:@54910.4]
  wire  regs_370_io_enable; // @[RegFile.scala 66:20:@54910.4]
  wire  regs_371_clock; // @[RegFile.scala 66:20:@54924.4]
  wire  regs_371_reset; // @[RegFile.scala 66:20:@54924.4]
  wire [63:0] regs_371_io_in; // @[RegFile.scala 66:20:@54924.4]
  wire  regs_371_io_reset; // @[RegFile.scala 66:20:@54924.4]
  wire [63:0] regs_371_io_out; // @[RegFile.scala 66:20:@54924.4]
  wire  regs_371_io_enable; // @[RegFile.scala 66:20:@54924.4]
  wire  regs_372_clock; // @[RegFile.scala 66:20:@54938.4]
  wire  regs_372_reset; // @[RegFile.scala 66:20:@54938.4]
  wire [63:0] regs_372_io_in; // @[RegFile.scala 66:20:@54938.4]
  wire  regs_372_io_reset; // @[RegFile.scala 66:20:@54938.4]
  wire [63:0] regs_372_io_out; // @[RegFile.scala 66:20:@54938.4]
  wire  regs_372_io_enable; // @[RegFile.scala 66:20:@54938.4]
  wire  regs_373_clock; // @[RegFile.scala 66:20:@54952.4]
  wire  regs_373_reset; // @[RegFile.scala 66:20:@54952.4]
  wire [63:0] regs_373_io_in; // @[RegFile.scala 66:20:@54952.4]
  wire  regs_373_io_reset; // @[RegFile.scala 66:20:@54952.4]
  wire [63:0] regs_373_io_out; // @[RegFile.scala 66:20:@54952.4]
  wire  regs_373_io_enable; // @[RegFile.scala 66:20:@54952.4]
  wire  regs_374_clock; // @[RegFile.scala 66:20:@54966.4]
  wire  regs_374_reset; // @[RegFile.scala 66:20:@54966.4]
  wire [63:0] regs_374_io_in; // @[RegFile.scala 66:20:@54966.4]
  wire  regs_374_io_reset; // @[RegFile.scala 66:20:@54966.4]
  wire [63:0] regs_374_io_out; // @[RegFile.scala 66:20:@54966.4]
  wire  regs_374_io_enable; // @[RegFile.scala 66:20:@54966.4]
  wire  regs_375_clock; // @[RegFile.scala 66:20:@54980.4]
  wire  regs_375_reset; // @[RegFile.scala 66:20:@54980.4]
  wire [63:0] regs_375_io_in; // @[RegFile.scala 66:20:@54980.4]
  wire  regs_375_io_reset; // @[RegFile.scala 66:20:@54980.4]
  wire [63:0] regs_375_io_out; // @[RegFile.scala 66:20:@54980.4]
  wire  regs_375_io_enable; // @[RegFile.scala 66:20:@54980.4]
  wire  regs_376_clock; // @[RegFile.scala 66:20:@54994.4]
  wire  regs_376_reset; // @[RegFile.scala 66:20:@54994.4]
  wire [63:0] regs_376_io_in; // @[RegFile.scala 66:20:@54994.4]
  wire  regs_376_io_reset; // @[RegFile.scala 66:20:@54994.4]
  wire [63:0] regs_376_io_out; // @[RegFile.scala 66:20:@54994.4]
  wire  regs_376_io_enable; // @[RegFile.scala 66:20:@54994.4]
  wire  regs_377_clock; // @[RegFile.scala 66:20:@55008.4]
  wire  regs_377_reset; // @[RegFile.scala 66:20:@55008.4]
  wire [63:0] regs_377_io_in; // @[RegFile.scala 66:20:@55008.4]
  wire  regs_377_io_reset; // @[RegFile.scala 66:20:@55008.4]
  wire [63:0] regs_377_io_out; // @[RegFile.scala 66:20:@55008.4]
  wire  regs_377_io_enable; // @[RegFile.scala 66:20:@55008.4]
  wire  regs_378_clock; // @[RegFile.scala 66:20:@55022.4]
  wire  regs_378_reset; // @[RegFile.scala 66:20:@55022.4]
  wire [63:0] regs_378_io_in; // @[RegFile.scala 66:20:@55022.4]
  wire  regs_378_io_reset; // @[RegFile.scala 66:20:@55022.4]
  wire [63:0] regs_378_io_out; // @[RegFile.scala 66:20:@55022.4]
  wire  regs_378_io_enable; // @[RegFile.scala 66:20:@55022.4]
  wire  regs_379_clock; // @[RegFile.scala 66:20:@55036.4]
  wire  regs_379_reset; // @[RegFile.scala 66:20:@55036.4]
  wire [63:0] regs_379_io_in; // @[RegFile.scala 66:20:@55036.4]
  wire  regs_379_io_reset; // @[RegFile.scala 66:20:@55036.4]
  wire [63:0] regs_379_io_out; // @[RegFile.scala 66:20:@55036.4]
  wire  regs_379_io_enable; // @[RegFile.scala 66:20:@55036.4]
  wire  regs_380_clock; // @[RegFile.scala 66:20:@55050.4]
  wire  regs_380_reset; // @[RegFile.scala 66:20:@55050.4]
  wire [63:0] regs_380_io_in; // @[RegFile.scala 66:20:@55050.4]
  wire  regs_380_io_reset; // @[RegFile.scala 66:20:@55050.4]
  wire [63:0] regs_380_io_out; // @[RegFile.scala 66:20:@55050.4]
  wire  regs_380_io_enable; // @[RegFile.scala 66:20:@55050.4]
  wire  regs_381_clock; // @[RegFile.scala 66:20:@55064.4]
  wire  regs_381_reset; // @[RegFile.scala 66:20:@55064.4]
  wire [63:0] regs_381_io_in; // @[RegFile.scala 66:20:@55064.4]
  wire  regs_381_io_reset; // @[RegFile.scala 66:20:@55064.4]
  wire [63:0] regs_381_io_out; // @[RegFile.scala 66:20:@55064.4]
  wire  regs_381_io_enable; // @[RegFile.scala 66:20:@55064.4]
  wire  regs_382_clock; // @[RegFile.scala 66:20:@55078.4]
  wire  regs_382_reset; // @[RegFile.scala 66:20:@55078.4]
  wire [63:0] regs_382_io_in; // @[RegFile.scala 66:20:@55078.4]
  wire  regs_382_io_reset; // @[RegFile.scala 66:20:@55078.4]
  wire [63:0] regs_382_io_out; // @[RegFile.scala 66:20:@55078.4]
  wire  regs_382_io_enable; // @[RegFile.scala 66:20:@55078.4]
  wire  regs_383_clock; // @[RegFile.scala 66:20:@55092.4]
  wire  regs_383_reset; // @[RegFile.scala 66:20:@55092.4]
  wire [63:0] regs_383_io_in; // @[RegFile.scala 66:20:@55092.4]
  wire  regs_383_io_reset; // @[RegFile.scala 66:20:@55092.4]
  wire [63:0] regs_383_io_out; // @[RegFile.scala 66:20:@55092.4]
  wire  regs_383_io_enable; // @[RegFile.scala 66:20:@55092.4]
  wire  regs_384_clock; // @[RegFile.scala 66:20:@55106.4]
  wire  regs_384_reset; // @[RegFile.scala 66:20:@55106.4]
  wire [63:0] regs_384_io_in; // @[RegFile.scala 66:20:@55106.4]
  wire  regs_384_io_reset; // @[RegFile.scala 66:20:@55106.4]
  wire [63:0] regs_384_io_out; // @[RegFile.scala 66:20:@55106.4]
  wire  regs_384_io_enable; // @[RegFile.scala 66:20:@55106.4]
  wire  regs_385_clock; // @[RegFile.scala 66:20:@55120.4]
  wire  regs_385_reset; // @[RegFile.scala 66:20:@55120.4]
  wire [63:0] regs_385_io_in; // @[RegFile.scala 66:20:@55120.4]
  wire  regs_385_io_reset; // @[RegFile.scala 66:20:@55120.4]
  wire [63:0] regs_385_io_out; // @[RegFile.scala 66:20:@55120.4]
  wire  regs_385_io_enable; // @[RegFile.scala 66:20:@55120.4]
  wire  regs_386_clock; // @[RegFile.scala 66:20:@55134.4]
  wire  regs_386_reset; // @[RegFile.scala 66:20:@55134.4]
  wire [63:0] regs_386_io_in; // @[RegFile.scala 66:20:@55134.4]
  wire  regs_386_io_reset; // @[RegFile.scala 66:20:@55134.4]
  wire [63:0] regs_386_io_out; // @[RegFile.scala 66:20:@55134.4]
  wire  regs_386_io_enable; // @[RegFile.scala 66:20:@55134.4]
  wire  regs_387_clock; // @[RegFile.scala 66:20:@55148.4]
  wire  regs_387_reset; // @[RegFile.scala 66:20:@55148.4]
  wire [63:0] regs_387_io_in; // @[RegFile.scala 66:20:@55148.4]
  wire  regs_387_io_reset; // @[RegFile.scala 66:20:@55148.4]
  wire [63:0] regs_387_io_out; // @[RegFile.scala 66:20:@55148.4]
  wire  regs_387_io_enable; // @[RegFile.scala 66:20:@55148.4]
  wire  regs_388_clock; // @[RegFile.scala 66:20:@55162.4]
  wire  regs_388_reset; // @[RegFile.scala 66:20:@55162.4]
  wire [63:0] regs_388_io_in; // @[RegFile.scala 66:20:@55162.4]
  wire  regs_388_io_reset; // @[RegFile.scala 66:20:@55162.4]
  wire [63:0] regs_388_io_out; // @[RegFile.scala 66:20:@55162.4]
  wire  regs_388_io_enable; // @[RegFile.scala 66:20:@55162.4]
  wire  regs_389_clock; // @[RegFile.scala 66:20:@55176.4]
  wire  regs_389_reset; // @[RegFile.scala 66:20:@55176.4]
  wire [63:0] regs_389_io_in; // @[RegFile.scala 66:20:@55176.4]
  wire  regs_389_io_reset; // @[RegFile.scala 66:20:@55176.4]
  wire [63:0] regs_389_io_out; // @[RegFile.scala 66:20:@55176.4]
  wire  regs_389_io_enable; // @[RegFile.scala 66:20:@55176.4]
  wire  regs_390_clock; // @[RegFile.scala 66:20:@55190.4]
  wire  regs_390_reset; // @[RegFile.scala 66:20:@55190.4]
  wire [63:0] regs_390_io_in; // @[RegFile.scala 66:20:@55190.4]
  wire  regs_390_io_reset; // @[RegFile.scala 66:20:@55190.4]
  wire [63:0] regs_390_io_out; // @[RegFile.scala 66:20:@55190.4]
  wire  regs_390_io_enable; // @[RegFile.scala 66:20:@55190.4]
  wire  regs_391_clock; // @[RegFile.scala 66:20:@55204.4]
  wire  regs_391_reset; // @[RegFile.scala 66:20:@55204.4]
  wire [63:0] regs_391_io_in; // @[RegFile.scala 66:20:@55204.4]
  wire  regs_391_io_reset; // @[RegFile.scala 66:20:@55204.4]
  wire [63:0] regs_391_io_out; // @[RegFile.scala 66:20:@55204.4]
  wire  regs_391_io_enable; // @[RegFile.scala 66:20:@55204.4]
  wire  regs_392_clock; // @[RegFile.scala 66:20:@55218.4]
  wire  regs_392_reset; // @[RegFile.scala 66:20:@55218.4]
  wire [63:0] regs_392_io_in; // @[RegFile.scala 66:20:@55218.4]
  wire  regs_392_io_reset; // @[RegFile.scala 66:20:@55218.4]
  wire [63:0] regs_392_io_out; // @[RegFile.scala 66:20:@55218.4]
  wire  regs_392_io_enable; // @[RegFile.scala 66:20:@55218.4]
  wire  regs_393_clock; // @[RegFile.scala 66:20:@55232.4]
  wire  regs_393_reset; // @[RegFile.scala 66:20:@55232.4]
  wire [63:0] regs_393_io_in; // @[RegFile.scala 66:20:@55232.4]
  wire  regs_393_io_reset; // @[RegFile.scala 66:20:@55232.4]
  wire [63:0] regs_393_io_out; // @[RegFile.scala 66:20:@55232.4]
  wire  regs_393_io_enable; // @[RegFile.scala 66:20:@55232.4]
  wire  regs_394_clock; // @[RegFile.scala 66:20:@55246.4]
  wire  regs_394_reset; // @[RegFile.scala 66:20:@55246.4]
  wire [63:0] regs_394_io_in; // @[RegFile.scala 66:20:@55246.4]
  wire  regs_394_io_reset; // @[RegFile.scala 66:20:@55246.4]
  wire [63:0] regs_394_io_out; // @[RegFile.scala 66:20:@55246.4]
  wire  regs_394_io_enable; // @[RegFile.scala 66:20:@55246.4]
  wire  regs_395_clock; // @[RegFile.scala 66:20:@55260.4]
  wire  regs_395_reset; // @[RegFile.scala 66:20:@55260.4]
  wire [63:0] regs_395_io_in; // @[RegFile.scala 66:20:@55260.4]
  wire  regs_395_io_reset; // @[RegFile.scala 66:20:@55260.4]
  wire [63:0] regs_395_io_out; // @[RegFile.scala 66:20:@55260.4]
  wire  regs_395_io_enable; // @[RegFile.scala 66:20:@55260.4]
  wire  regs_396_clock; // @[RegFile.scala 66:20:@55274.4]
  wire  regs_396_reset; // @[RegFile.scala 66:20:@55274.4]
  wire [63:0] regs_396_io_in; // @[RegFile.scala 66:20:@55274.4]
  wire  regs_396_io_reset; // @[RegFile.scala 66:20:@55274.4]
  wire [63:0] regs_396_io_out; // @[RegFile.scala 66:20:@55274.4]
  wire  regs_396_io_enable; // @[RegFile.scala 66:20:@55274.4]
  wire  regs_397_clock; // @[RegFile.scala 66:20:@55288.4]
  wire  regs_397_reset; // @[RegFile.scala 66:20:@55288.4]
  wire [63:0] regs_397_io_in; // @[RegFile.scala 66:20:@55288.4]
  wire  regs_397_io_reset; // @[RegFile.scala 66:20:@55288.4]
  wire [63:0] regs_397_io_out; // @[RegFile.scala 66:20:@55288.4]
  wire  regs_397_io_enable; // @[RegFile.scala 66:20:@55288.4]
  wire  regs_398_clock; // @[RegFile.scala 66:20:@55302.4]
  wire  regs_398_reset; // @[RegFile.scala 66:20:@55302.4]
  wire [63:0] regs_398_io_in; // @[RegFile.scala 66:20:@55302.4]
  wire  regs_398_io_reset; // @[RegFile.scala 66:20:@55302.4]
  wire [63:0] regs_398_io_out; // @[RegFile.scala 66:20:@55302.4]
  wire  regs_398_io_enable; // @[RegFile.scala 66:20:@55302.4]
  wire  regs_399_clock; // @[RegFile.scala 66:20:@55316.4]
  wire  regs_399_reset; // @[RegFile.scala 66:20:@55316.4]
  wire [63:0] regs_399_io_in; // @[RegFile.scala 66:20:@55316.4]
  wire  regs_399_io_reset; // @[RegFile.scala 66:20:@55316.4]
  wire [63:0] regs_399_io_out; // @[RegFile.scala 66:20:@55316.4]
  wire  regs_399_io_enable; // @[RegFile.scala 66:20:@55316.4]
  wire  regs_400_clock; // @[RegFile.scala 66:20:@55330.4]
  wire  regs_400_reset; // @[RegFile.scala 66:20:@55330.4]
  wire [63:0] regs_400_io_in; // @[RegFile.scala 66:20:@55330.4]
  wire  regs_400_io_reset; // @[RegFile.scala 66:20:@55330.4]
  wire [63:0] regs_400_io_out; // @[RegFile.scala 66:20:@55330.4]
  wire  regs_400_io_enable; // @[RegFile.scala 66:20:@55330.4]
  wire  regs_401_clock; // @[RegFile.scala 66:20:@55344.4]
  wire  regs_401_reset; // @[RegFile.scala 66:20:@55344.4]
  wire [63:0] regs_401_io_in; // @[RegFile.scala 66:20:@55344.4]
  wire  regs_401_io_reset; // @[RegFile.scala 66:20:@55344.4]
  wire [63:0] regs_401_io_out; // @[RegFile.scala 66:20:@55344.4]
  wire  regs_401_io_enable; // @[RegFile.scala 66:20:@55344.4]
  wire  regs_402_clock; // @[RegFile.scala 66:20:@55358.4]
  wire  regs_402_reset; // @[RegFile.scala 66:20:@55358.4]
  wire [63:0] regs_402_io_in; // @[RegFile.scala 66:20:@55358.4]
  wire  regs_402_io_reset; // @[RegFile.scala 66:20:@55358.4]
  wire [63:0] regs_402_io_out; // @[RegFile.scala 66:20:@55358.4]
  wire  regs_402_io_enable; // @[RegFile.scala 66:20:@55358.4]
  wire  regs_403_clock; // @[RegFile.scala 66:20:@55372.4]
  wire  regs_403_reset; // @[RegFile.scala 66:20:@55372.4]
  wire [63:0] regs_403_io_in; // @[RegFile.scala 66:20:@55372.4]
  wire  regs_403_io_reset; // @[RegFile.scala 66:20:@55372.4]
  wire [63:0] regs_403_io_out; // @[RegFile.scala 66:20:@55372.4]
  wire  regs_403_io_enable; // @[RegFile.scala 66:20:@55372.4]
  wire  regs_404_clock; // @[RegFile.scala 66:20:@55386.4]
  wire  regs_404_reset; // @[RegFile.scala 66:20:@55386.4]
  wire [63:0] regs_404_io_in; // @[RegFile.scala 66:20:@55386.4]
  wire  regs_404_io_reset; // @[RegFile.scala 66:20:@55386.4]
  wire [63:0] regs_404_io_out; // @[RegFile.scala 66:20:@55386.4]
  wire  regs_404_io_enable; // @[RegFile.scala 66:20:@55386.4]
  wire  regs_405_clock; // @[RegFile.scala 66:20:@55400.4]
  wire  regs_405_reset; // @[RegFile.scala 66:20:@55400.4]
  wire [63:0] regs_405_io_in; // @[RegFile.scala 66:20:@55400.4]
  wire  regs_405_io_reset; // @[RegFile.scala 66:20:@55400.4]
  wire [63:0] regs_405_io_out; // @[RegFile.scala 66:20:@55400.4]
  wire  regs_405_io_enable; // @[RegFile.scala 66:20:@55400.4]
  wire  regs_406_clock; // @[RegFile.scala 66:20:@55414.4]
  wire  regs_406_reset; // @[RegFile.scala 66:20:@55414.4]
  wire [63:0] regs_406_io_in; // @[RegFile.scala 66:20:@55414.4]
  wire  regs_406_io_reset; // @[RegFile.scala 66:20:@55414.4]
  wire [63:0] regs_406_io_out; // @[RegFile.scala 66:20:@55414.4]
  wire  regs_406_io_enable; // @[RegFile.scala 66:20:@55414.4]
  wire  regs_407_clock; // @[RegFile.scala 66:20:@55428.4]
  wire  regs_407_reset; // @[RegFile.scala 66:20:@55428.4]
  wire [63:0] regs_407_io_in; // @[RegFile.scala 66:20:@55428.4]
  wire  regs_407_io_reset; // @[RegFile.scala 66:20:@55428.4]
  wire [63:0] regs_407_io_out; // @[RegFile.scala 66:20:@55428.4]
  wire  regs_407_io_enable; // @[RegFile.scala 66:20:@55428.4]
  wire  regs_408_clock; // @[RegFile.scala 66:20:@55442.4]
  wire  regs_408_reset; // @[RegFile.scala 66:20:@55442.4]
  wire [63:0] regs_408_io_in; // @[RegFile.scala 66:20:@55442.4]
  wire  regs_408_io_reset; // @[RegFile.scala 66:20:@55442.4]
  wire [63:0] regs_408_io_out; // @[RegFile.scala 66:20:@55442.4]
  wire  regs_408_io_enable; // @[RegFile.scala 66:20:@55442.4]
  wire  regs_409_clock; // @[RegFile.scala 66:20:@55456.4]
  wire  regs_409_reset; // @[RegFile.scala 66:20:@55456.4]
  wire [63:0] regs_409_io_in; // @[RegFile.scala 66:20:@55456.4]
  wire  regs_409_io_reset; // @[RegFile.scala 66:20:@55456.4]
  wire [63:0] regs_409_io_out; // @[RegFile.scala 66:20:@55456.4]
  wire  regs_409_io_enable; // @[RegFile.scala 66:20:@55456.4]
  wire  regs_410_clock; // @[RegFile.scala 66:20:@55470.4]
  wire  regs_410_reset; // @[RegFile.scala 66:20:@55470.4]
  wire [63:0] regs_410_io_in; // @[RegFile.scala 66:20:@55470.4]
  wire  regs_410_io_reset; // @[RegFile.scala 66:20:@55470.4]
  wire [63:0] regs_410_io_out; // @[RegFile.scala 66:20:@55470.4]
  wire  regs_410_io_enable; // @[RegFile.scala 66:20:@55470.4]
  wire  regs_411_clock; // @[RegFile.scala 66:20:@55484.4]
  wire  regs_411_reset; // @[RegFile.scala 66:20:@55484.4]
  wire [63:0] regs_411_io_in; // @[RegFile.scala 66:20:@55484.4]
  wire  regs_411_io_reset; // @[RegFile.scala 66:20:@55484.4]
  wire [63:0] regs_411_io_out; // @[RegFile.scala 66:20:@55484.4]
  wire  regs_411_io_enable; // @[RegFile.scala 66:20:@55484.4]
  wire  regs_412_clock; // @[RegFile.scala 66:20:@55498.4]
  wire  regs_412_reset; // @[RegFile.scala 66:20:@55498.4]
  wire [63:0] regs_412_io_in; // @[RegFile.scala 66:20:@55498.4]
  wire  regs_412_io_reset; // @[RegFile.scala 66:20:@55498.4]
  wire [63:0] regs_412_io_out; // @[RegFile.scala 66:20:@55498.4]
  wire  regs_412_io_enable; // @[RegFile.scala 66:20:@55498.4]
  wire  regs_413_clock; // @[RegFile.scala 66:20:@55512.4]
  wire  regs_413_reset; // @[RegFile.scala 66:20:@55512.4]
  wire [63:0] regs_413_io_in; // @[RegFile.scala 66:20:@55512.4]
  wire  regs_413_io_reset; // @[RegFile.scala 66:20:@55512.4]
  wire [63:0] regs_413_io_out; // @[RegFile.scala 66:20:@55512.4]
  wire  regs_413_io_enable; // @[RegFile.scala 66:20:@55512.4]
  wire  regs_414_clock; // @[RegFile.scala 66:20:@55526.4]
  wire  regs_414_reset; // @[RegFile.scala 66:20:@55526.4]
  wire [63:0] regs_414_io_in; // @[RegFile.scala 66:20:@55526.4]
  wire  regs_414_io_reset; // @[RegFile.scala 66:20:@55526.4]
  wire [63:0] regs_414_io_out; // @[RegFile.scala 66:20:@55526.4]
  wire  regs_414_io_enable; // @[RegFile.scala 66:20:@55526.4]
  wire  regs_415_clock; // @[RegFile.scala 66:20:@55540.4]
  wire  regs_415_reset; // @[RegFile.scala 66:20:@55540.4]
  wire [63:0] regs_415_io_in; // @[RegFile.scala 66:20:@55540.4]
  wire  regs_415_io_reset; // @[RegFile.scala 66:20:@55540.4]
  wire [63:0] regs_415_io_out; // @[RegFile.scala 66:20:@55540.4]
  wire  regs_415_io_enable; // @[RegFile.scala 66:20:@55540.4]
  wire  regs_416_clock; // @[RegFile.scala 66:20:@55554.4]
  wire  regs_416_reset; // @[RegFile.scala 66:20:@55554.4]
  wire [63:0] regs_416_io_in; // @[RegFile.scala 66:20:@55554.4]
  wire  regs_416_io_reset; // @[RegFile.scala 66:20:@55554.4]
  wire [63:0] regs_416_io_out; // @[RegFile.scala 66:20:@55554.4]
  wire  regs_416_io_enable; // @[RegFile.scala 66:20:@55554.4]
  wire  regs_417_clock; // @[RegFile.scala 66:20:@55568.4]
  wire  regs_417_reset; // @[RegFile.scala 66:20:@55568.4]
  wire [63:0] regs_417_io_in; // @[RegFile.scala 66:20:@55568.4]
  wire  regs_417_io_reset; // @[RegFile.scala 66:20:@55568.4]
  wire [63:0] regs_417_io_out; // @[RegFile.scala 66:20:@55568.4]
  wire  regs_417_io_enable; // @[RegFile.scala 66:20:@55568.4]
  wire  regs_418_clock; // @[RegFile.scala 66:20:@55582.4]
  wire  regs_418_reset; // @[RegFile.scala 66:20:@55582.4]
  wire [63:0] regs_418_io_in; // @[RegFile.scala 66:20:@55582.4]
  wire  regs_418_io_reset; // @[RegFile.scala 66:20:@55582.4]
  wire [63:0] regs_418_io_out; // @[RegFile.scala 66:20:@55582.4]
  wire  regs_418_io_enable; // @[RegFile.scala 66:20:@55582.4]
  wire  regs_419_clock; // @[RegFile.scala 66:20:@55596.4]
  wire  regs_419_reset; // @[RegFile.scala 66:20:@55596.4]
  wire [63:0] regs_419_io_in; // @[RegFile.scala 66:20:@55596.4]
  wire  regs_419_io_reset; // @[RegFile.scala 66:20:@55596.4]
  wire [63:0] regs_419_io_out; // @[RegFile.scala 66:20:@55596.4]
  wire  regs_419_io_enable; // @[RegFile.scala 66:20:@55596.4]
  wire  regs_420_clock; // @[RegFile.scala 66:20:@55610.4]
  wire  regs_420_reset; // @[RegFile.scala 66:20:@55610.4]
  wire [63:0] regs_420_io_in; // @[RegFile.scala 66:20:@55610.4]
  wire  regs_420_io_reset; // @[RegFile.scala 66:20:@55610.4]
  wire [63:0] regs_420_io_out; // @[RegFile.scala 66:20:@55610.4]
  wire  regs_420_io_enable; // @[RegFile.scala 66:20:@55610.4]
  wire  regs_421_clock; // @[RegFile.scala 66:20:@55624.4]
  wire  regs_421_reset; // @[RegFile.scala 66:20:@55624.4]
  wire [63:0] regs_421_io_in; // @[RegFile.scala 66:20:@55624.4]
  wire  regs_421_io_reset; // @[RegFile.scala 66:20:@55624.4]
  wire [63:0] regs_421_io_out; // @[RegFile.scala 66:20:@55624.4]
  wire  regs_421_io_enable; // @[RegFile.scala 66:20:@55624.4]
  wire  regs_422_clock; // @[RegFile.scala 66:20:@55638.4]
  wire  regs_422_reset; // @[RegFile.scala 66:20:@55638.4]
  wire [63:0] regs_422_io_in; // @[RegFile.scala 66:20:@55638.4]
  wire  regs_422_io_reset; // @[RegFile.scala 66:20:@55638.4]
  wire [63:0] regs_422_io_out; // @[RegFile.scala 66:20:@55638.4]
  wire  regs_422_io_enable; // @[RegFile.scala 66:20:@55638.4]
  wire  regs_423_clock; // @[RegFile.scala 66:20:@55652.4]
  wire  regs_423_reset; // @[RegFile.scala 66:20:@55652.4]
  wire [63:0] regs_423_io_in; // @[RegFile.scala 66:20:@55652.4]
  wire  regs_423_io_reset; // @[RegFile.scala 66:20:@55652.4]
  wire [63:0] regs_423_io_out; // @[RegFile.scala 66:20:@55652.4]
  wire  regs_423_io_enable; // @[RegFile.scala 66:20:@55652.4]
  wire  regs_424_clock; // @[RegFile.scala 66:20:@55666.4]
  wire  regs_424_reset; // @[RegFile.scala 66:20:@55666.4]
  wire [63:0] regs_424_io_in; // @[RegFile.scala 66:20:@55666.4]
  wire  regs_424_io_reset; // @[RegFile.scala 66:20:@55666.4]
  wire [63:0] regs_424_io_out; // @[RegFile.scala 66:20:@55666.4]
  wire  regs_424_io_enable; // @[RegFile.scala 66:20:@55666.4]
  wire  regs_425_clock; // @[RegFile.scala 66:20:@55680.4]
  wire  regs_425_reset; // @[RegFile.scala 66:20:@55680.4]
  wire [63:0] regs_425_io_in; // @[RegFile.scala 66:20:@55680.4]
  wire  regs_425_io_reset; // @[RegFile.scala 66:20:@55680.4]
  wire [63:0] regs_425_io_out; // @[RegFile.scala 66:20:@55680.4]
  wire  regs_425_io_enable; // @[RegFile.scala 66:20:@55680.4]
  wire  regs_426_clock; // @[RegFile.scala 66:20:@55694.4]
  wire  regs_426_reset; // @[RegFile.scala 66:20:@55694.4]
  wire [63:0] regs_426_io_in; // @[RegFile.scala 66:20:@55694.4]
  wire  regs_426_io_reset; // @[RegFile.scala 66:20:@55694.4]
  wire [63:0] regs_426_io_out; // @[RegFile.scala 66:20:@55694.4]
  wire  regs_426_io_enable; // @[RegFile.scala 66:20:@55694.4]
  wire  regs_427_clock; // @[RegFile.scala 66:20:@55708.4]
  wire  regs_427_reset; // @[RegFile.scala 66:20:@55708.4]
  wire [63:0] regs_427_io_in; // @[RegFile.scala 66:20:@55708.4]
  wire  regs_427_io_reset; // @[RegFile.scala 66:20:@55708.4]
  wire [63:0] regs_427_io_out; // @[RegFile.scala 66:20:@55708.4]
  wire  regs_427_io_enable; // @[RegFile.scala 66:20:@55708.4]
  wire  regs_428_clock; // @[RegFile.scala 66:20:@55722.4]
  wire  regs_428_reset; // @[RegFile.scala 66:20:@55722.4]
  wire [63:0] regs_428_io_in; // @[RegFile.scala 66:20:@55722.4]
  wire  regs_428_io_reset; // @[RegFile.scala 66:20:@55722.4]
  wire [63:0] regs_428_io_out; // @[RegFile.scala 66:20:@55722.4]
  wire  regs_428_io_enable; // @[RegFile.scala 66:20:@55722.4]
  wire  regs_429_clock; // @[RegFile.scala 66:20:@55736.4]
  wire  regs_429_reset; // @[RegFile.scala 66:20:@55736.4]
  wire [63:0] regs_429_io_in; // @[RegFile.scala 66:20:@55736.4]
  wire  regs_429_io_reset; // @[RegFile.scala 66:20:@55736.4]
  wire [63:0] regs_429_io_out; // @[RegFile.scala 66:20:@55736.4]
  wire  regs_429_io_enable; // @[RegFile.scala 66:20:@55736.4]
  wire  regs_430_clock; // @[RegFile.scala 66:20:@55750.4]
  wire  regs_430_reset; // @[RegFile.scala 66:20:@55750.4]
  wire [63:0] regs_430_io_in; // @[RegFile.scala 66:20:@55750.4]
  wire  regs_430_io_reset; // @[RegFile.scala 66:20:@55750.4]
  wire [63:0] regs_430_io_out; // @[RegFile.scala 66:20:@55750.4]
  wire  regs_430_io_enable; // @[RegFile.scala 66:20:@55750.4]
  wire  regs_431_clock; // @[RegFile.scala 66:20:@55764.4]
  wire  regs_431_reset; // @[RegFile.scala 66:20:@55764.4]
  wire [63:0] regs_431_io_in; // @[RegFile.scala 66:20:@55764.4]
  wire  regs_431_io_reset; // @[RegFile.scala 66:20:@55764.4]
  wire [63:0] regs_431_io_out; // @[RegFile.scala 66:20:@55764.4]
  wire  regs_431_io_enable; // @[RegFile.scala 66:20:@55764.4]
  wire  regs_432_clock; // @[RegFile.scala 66:20:@55778.4]
  wire  regs_432_reset; // @[RegFile.scala 66:20:@55778.4]
  wire [63:0] regs_432_io_in; // @[RegFile.scala 66:20:@55778.4]
  wire  regs_432_io_reset; // @[RegFile.scala 66:20:@55778.4]
  wire [63:0] regs_432_io_out; // @[RegFile.scala 66:20:@55778.4]
  wire  regs_432_io_enable; // @[RegFile.scala 66:20:@55778.4]
  wire  regs_433_clock; // @[RegFile.scala 66:20:@55792.4]
  wire  regs_433_reset; // @[RegFile.scala 66:20:@55792.4]
  wire [63:0] regs_433_io_in; // @[RegFile.scala 66:20:@55792.4]
  wire  regs_433_io_reset; // @[RegFile.scala 66:20:@55792.4]
  wire [63:0] regs_433_io_out; // @[RegFile.scala 66:20:@55792.4]
  wire  regs_433_io_enable; // @[RegFile.scala 66:20:@55792.4]
  wire  regs_434_clock; // @[RegFile.scala 66:20:@55806.4]
  wire  regs_434_reset; // @[RegFile.scala 66:20:@55806.4]
  wire [63:0] regs_434_io_in; // @[RegFile.scala 66:20:@55806.4]
  wire  regs_434_io_reset; // @[RegFile.scala 66:20:@55806.4]
  wire [63:0] regs_434_io_out; // @[RegFile.scala 66:20:@55806.4]
  wire  regs_434_io_enable; // @[RegFile.scala 66:20:@55806.4]
  wire  regs_435_clock; // @[RegFile.scala 66:20:@55820.4]
  wire  regs_435_reset; // @[RegFile.scala 66:20:@55820.4]
  wire [63:0] regs_435_io_in; // @[RegFile.scala 66:20:@55820.4]
  wire  regs_435_io_reset; // @[RegFile.scala 66:20:@55820.4]
  wire [63:0] regs_435_io_out; // @[RegFile.scala 66:20:@55820.4]
  wire  regs_435_io_enable; // @[RegFile.scala 66:20:@55820.4]
  wire  regs_436_clock; // @[RegFile.scala 66:20:@55834.4]
  wire  regs_436_reset; // @[RegFile.scala 66:20:@55834.4]
  wire [63:0] regs_436_io_in; // @[RegFile.scala 66:20:@55834.4]
  wire  regs_436_io_reset; // @[RegFile.scala 66:20:@55834.4]
  wire [63:0] regs_436_io_out; // @[RegFile.scala 66:20:@55834.4]
  wire  regs_436_io_enable; // @[RegFile.scala 66:20:@55834.4]
  wire  regs_437_clock; // @[RegFile.scala 66:20:@55848.4]
  wire  regs_437_reset; // @[RegFile.scala 66:20:@55848.4]
  wire [63:0] regs_437_io_in; // @[RegFile.scala 66:20:@55848.4]
  wire  regs_437_io_reset; // @[RegFile.scala 66:20:@55848.4]
  wire [63:0] regs_437_io_out; // @[RegFile.scala 66:20:@55848.4]
  wire  regs_437_io_enable; // @[RegFile.scala 66:20:@55848.4]
  wire  regs_438_clock; // @[RegFile.scala 66:20:@55862.4]
  wire  regs_438_reset; // @[RegFile.scala 66:20:@55862.4]
  wire [63:0] regs_438_io_in; // @[RegFile.scala 66:20:@55862.4]
  wire  regs_438_io_reset; // @[RegFile.scala 66:20:@55862.4]
  wire [63:0] regs_438_io_out; // @[RegFile.scala 66:20:@55862.4]
  wire  regs_438_io_enable; // @[RegFile.scala 66:20:@55862.4]
  wire  regs_439_clock; // @[RegFile.scala 66:20:@55876.4]
  wire  regs_439_reset; // @[RegFile.scala 66:20:@55876.4]
  wire [63:0] regs_439_io_in; // @[RegFile.scala 66:20:@55876.4]
  wire  regs_439_io_reset; // @[RegFile.scala 66:20:@55876.4]
  wire [63:0] regs_439_io_out; // @[RegFile.scala 66:20:@55876.4]
  wire  regs_439_io_enable; // @[RegFile.scala 66:20:@55876.4]
  wire  regs_440_clock; // @[RegFile.scala 66:20:@55890.4]
  wire  regs_440_reset; // @[RegFile.scala 66:20:@55890.4]
  wire [63:0] regs_440_io_in; // @[RegFile.scala 66:20:@55890.4]
  wire  regs_440_io_reset; // @[RegFile.scala 66:20:@55890.4]
  wire [63:0] regs_440_io_out; // @[RegFile.scala 66:20:@55890.4]
  wire  regs_440_io_enable; // @[RegFile.scala 66:20:@55890.4]
  wire  regs_441_clock; // @[RegFile.scala 66:20:@55904.4]
  wire  regs_441_reset; // @[RegFile.scala 66:20:@55904.4]
  wire [63:0] regs_441_io_in; // @[RegFile.scala 66:20:@55904.4]
  wire  regs_441_io_reset; // @[RegFile.scala 66:20:@55904.4]
  wire [63:0] regs_441_io_out; // @[RegFile.scala 66:20:@55904.4]
  wire  regs_441_io_enable; // @[RegFile.scala 66:20:@55904.4]
  wire  regs_442_clock; // @[RegFile.scala 66:20:@55918.4]
  wire  regs_442_reset; // @[RegFile.scala 66:20:@55918.4]
  wire [63:0] regs_442_io_in; // @[RegFile.scala 66:20:@55918.4]
  wire  regs_442_io_reset; // @[RegFile.scala 66:20:@55918.4]
  wire [63:0] regs_442_io_out; // @[RegFile.scala 66:20:@55918.4]
  wire  regs_442_io_enable; // @[RegFile.scala 66:20:@55918.4]
  wire  regs_443_clock; // @[RegFile.scala 66:20:@55932.4]
  wire  regs_443_reset; // @[RegFile.scala 66:20:@55932.4]
  wire [63:0] regs_443_io_in; // @[RegFile.scala 66:20:@55932.4]
  wire  regs_443_io_reset; // @[RegFile.scala 66:20:@55932.4]
  wire [63:0] regs_443_io_out; // @[RegFile.scala 66:20:@55932.4]
  wire  regs_443_io_enable; // @[RegFile.scala 66:20:@55932.4]
  wire  regs_444_clock; // @[RegFile.scala 66:20:@55946.4]
  wire  regs_444_reset; // @[RegFile.scala 66:20:@55946.4]
  wire [63:0] regs_444_io_in; // @[RegFile.scala 66:20:@55946.4]
  wire  regs_444_io_reset; // @[RegFile.scala 66:20:@55946.4]
  wire [63:0] regs_444_io_out; // @[RegFile.scala 66:20:@55946.4]
  wire  regs_444_io_enable; // @[RegFile.scala 66:20:@55946.4]
  wire  regs_445_clock; // @[RegFile.scala 66:20:@55960.4]
  wire  regs_445_reset; // @[RegFile.scala 66:20:@55960.4]
  wire [63:0] regs_445_io_in; // @[RegFile.scala 66:20:@55960.4]
  wire  regs_445_io_reset; // @[RegFile.scala 66:20:@55960.4]
  wire [63:0] regs_445_io_out; // @[RegFile.scala 66:20:@55960.4]
  wire  regs_445_io_enable; // @[RegFile.scala 66:20:@55960.4]
  wire  regs_446_clock; // @[RegFile.scala 66:20:@55974.4]
  wire  regs_446_reset; // @[RegFile.scala 66:20:@55974.4]
  wire [63:0] regs_446_io_in; // @[RegFile.scala 66:20:@55974.4]
  wire  regs_446_io_reset; // @[RegFile.scala 66:20:@55974.4]
  wire [63:0] regs_446_io_out; // @[RegFile.scala 66:20:@55974.4]
  wire  regs_446_io_enable; // @[RegFile.scala 66:20:@55974.4]
  wire  regs_447_clock; // @[RegFile.scala 66:20:@55988.4]
  wire  regs_447_reset; // @[RegFile.scala 66:20:@55988.4]
  wire [63:0] regs_447_io_in; // @[RegFile.scala 66:20:@55988.4]
  wire  regs_447_io_reset; // @[RegFile.scala 66:20:@55988.4]
  wire [63:0] regs_447_io_out; // @[RegFile.scala 66:20:@55988.4]
  wire  regs_447_io_enable; // @[RegFile.scala 66:20:@55988.4]
  wire  regs_448_clock; // @[RegFile.scala 66:20:@56002.4]
  wire  regs_448_reset; // @[RegFile.scala 66:20:@56002.4]
  wire [63:0] regs_448_io_in; // @[RegFile.scala 66:20:@56002.4]
  wire  regs_448_io_reset; // @[RegFile.scala 66:20:@56002.4]
  wire [63:0] regs_448_io_out; // @[RegFile.scala 66:20:@56002.4]
  wire  regs_448_io_enable; // @[RegFile.scala 66:20:@56002.4]
  wire  regs_449_clock; // @[RegFile.scala 66:20:@56016.4]
  wire  regs_449_reset; // @[RegFile.scala 66:20:@56016.4]
  wire [63:0] regs_449_io_in; // @[RegFile.scala 66:20:@56016.4]
  wire  regs_449_io_reset; // @[RegFile.scala 66:20:@56016.4]
  wire [63:0] regs_449_io_out; // @[RegFile.scala 66:20:@56016.4]
  wire  regs_449_io_enable; // @[RegFile.scala 66:20:@56016.4]
  wire  regs_450_clock; // @[RegFile.scala 66:20:@56030.4]
  wire  regs_450_reset; // @[RegFile.scala 66:20:@56030.4]
  wire [63:0] regs_450_io_in; // @[RegFile.scala 66:20:@56030.4]
  wire  regs_450_io_reset; // @[RegFile.scala 66:20:@56030.4]
  wire [63:0] regs_450_io_out; // @[RegFile.scala 66:20:@56030.4]
  wire  regs_450_io_enable; // @[RegFile.scala 66:20:@56030.4]
  wire  regs_451_clock; // @[RegFile.scala 66:20:@56044.4]
  wire  regs_451_reset; // @[RegFile.scala 66:20:@56044.4]
  wire [63:0] regs_451_io_in; // @[RegFile.scala 66:20:@56044.4]
  wire  regs_451_io_reset; // @[RegFile.scala 66:20:@56044.4]
  wire [63:0] regs_451_io_out; // @[RegFile.scala 66:20:@56044.4]
  wire  regs_451_io_enable; // @[RegFile.scala 66:20:@56044.4]
  wire  regs_452_clock; // @[RegFile.scala 66:20:@56058.4]
  wire  regs_452_reset; // @[RegFile.scala 66:20:@56058.4]
  wire [63:0] regs_452_io_in; // @[RegFile.scala 66:20:@56058.4]
  wire  regs_452_io_reset; // @[RegFile.scala 66:20:@56058.4]
  wire [63:0] regs_452_io_out; // @[RegFile.scala 66:20:@56058.4]
  wire  regs_452_io_enable; // @[RegFile.scala 66:20:@56058.4]
  wire  regs_453_clock; // @[RegFile.scala 66:20:@56072.4]
  wire  regs_453_reset; // @[RegFile.scala 66:20:@56072.4]
  wire [63:0] regs_453_io_in; // @[RegFile.scala 66:20:@56072.4]
  wire  regs_453_io_reset; // @[RegFile.scala 66:20:@56072.4]
  wire [63:0] regs_453_io_out; // @[RegFile.scala 66:20:@56072.4]
  wire  regs_453_io_enable; // @[RegFile.scala 66:20:@56072.4]
  wire  regs_454_clock; // @[RegFile.scala 66:20:@56086.4]
  wire  regs_454_reset; // @[RegFile.scala 66:20:@56086.4]
  wire [63:0] regs_454_io_in; // @[RegFile.scala 66:20:@56086.4]
  wire  regs_454_io_reset; // @[RegFile.scala 66:20:@56086.4]
  wire [63:0] regs_454_io_out; // @[RegFile.scala 66:20:@56086.4]
  wire  regs_454_io_enable; // @[RegFile.scala 66:20:@56086.4]
  wire  regs_455_clock; // @[RegFile.scala 66:20:@56100.4]
  wire  regs_455_reset; // @[RegFile.scala 66:20:@56100.4]
  wire [63:0] regs_455_io_in; // @[RegFile.scala 66:20:@56100.4]
  wire  regs_455_io_reset; // @[RegFile.scala 66:20:@56100.4]
  wire [63:0] regs_455_io_out; // @[RegFile.scala 66:20:@56100.4]
  wire  regs_455_io_enable; // @[RegFile.scala 66:20:@56100.4]
  wire  regs_456_clock; // @[RegFile.scala 66:20:@56114.4]
  wire  regs_456_reset; // @[RegFile.scala 66:20:@56114.4]
  wire [63:0] regs_456_io_in; // @[RegFile.scala 66:20:@56114.4]
  wire  regs_456_io_reset; // @[RegFile.scala 66:20:@56114.4]
  wire [63:0] regs_456_io_out; // @[RegFile.scala 66:20:@56114.4]
  wire  regs_456_io_enable; // @[RegFile.scala 66:20:@56114.4]
  wire  regs_457_clock; // @[RegFile.scala 66:20:@56128.4]
  wire  regs_457_reset; // @[RegFile.scala 66:20:@56128.4]
  wire [63:0] regs_457_io_in; // @[RegFile.scala 66:20:@56128.4]
  wire  regs_457_io_reset; // @[RegFile.scala 66:20:@56128.4]
  wire [63:0] regs_457_io_out; // @[RegFile.scala 66:20:@56128.4]
  wire  regs_457_io_enable; // @[RegFile.scala 66:20:@56128.4]
  wire  regs_458_clock; // @[RegFile.scala 66:20:@56142.4]
  wire  regs_458_reset; // @[RegFile.scala 66:20:@56142.4]
  wire [63:0] regs_458_io_in; // @[RegFile.scala 66:20:@56142.4]
  wire  regs_458_io_reset; // @[RegFile.scala 66:20:@56142.4]
  wire [63:0] regs_458_io_out; // @[RegFile.scala 66:20:@56142.4]
  wire  regs_458_io_enable; // @[RegFile.scala 66:20:@56142.4]
  wire  regs_459_clock; // @[RegFile.scala 66:20:@56156.4]
  wire  regs_459_reset; // @[RegFile.scala 66:20:@56156.4]
  wire [63:0] regs_459_io_in; // @[RegFile.scala 66:20:@56156.4]
  wire  regs_459_io_reset; // @[RegFile.scala 66:20:@56156.4]
  wire [63:0] regs_459_io_out; // @[RegFile.scala 66:20:@56156.4]
  wire  regs_459_io_enable; // @[RegFile.scala 66:20:@56156.4]
  wire  regs_460_clock; // @[RegFile.scala 66:20:@56170.4]
  wire  regs_460_reset; // @[RegFile.scala 66:20:@56170.4]
  wire [63:0] regs_460_io_in; // @[RegFile.scala 66:20:@56170.4]
  wire  regs_460_io_reset; // @[RegFile.scala 66:20:@56170.4]
  wire [63:0] regs_460_io_out; // @[RegFile.scala 66:20:@56170.4]
  wire  regs_460_io_enable; // @[RegFile.scala 66:20:@56170.4]
  wire  regs_461_clock; // @[RegFile.scala 66:20:@56184.4]
  wire  regs_461_reset; // @[RegFile.scala 66:20:@56184.4]
  wire [63:0] regs_461_io_in; // @[RegFile.scala 66:20:@56184.4]
  wire  regs_461_io_reset; // @[RegFile.scala 66:20:@56184.4]
  wire [63:0] regs_461_io_out; // @[RegFile.scala 66:20:@56184.4]
  wire  regs_461_io_enable; // @[RegFile.scala 66:20:@56184.4]
  wire  regs_462_clock; // @[RegFile.scala 66:20:@56198.4]
  wire  regs_462_reset; // @[RegFile.scala 66:20:@56198.4]
  wire [63:0] regs_462_io_in; // @[RegFile.scala 66:20:@56198.4]
  wire  regs_462_io_reset; // @[RegFile.scala 66:20:@56198.4]
  wire [63:0] regs_462_io_out; // @[RegFile.scala 66:20:@56198.4]
  wire  regs_462_io_enable; // @[RegFile.scala 66:20:@56198.4]
  wire  regs_463_clock; // @[RegFile.scala 66:20:@56212.4]
  wire  regs_463_reset; // @[RegFile.scala 66:20:@56212.4]
  wire [63:0] regs_463_io_in; // @[RegFile.scala 66:20:@56212.4]
  wire  regs_463_io_reset; // @[RegFile.scala 66:20:@56212.4]
  wire [63:0] regs_463_io_out; // @[RegFile.scala 66:20:@56212.4]
  wire  regs_463_io_enable; // @[RegFile.scala 66:20:@56212.4]
  wire  regs_464_clock; // @[RegFile.scala 66:20:@56226.4]
  wire  regs_464_reset; // @[RegFile.scala 66:20:@56226.4]
  wire [63:0] regs_464_io_in; // @[RegFile.scala 66:20:@56226.4]
  wire  regs_464_io_reset; // @[RegFile.scala 66:20:@56226.4]
  wire [63:0] regs_464_io_out; // @[RegFile.scala 66:20:@56226.4]
  wire  regs_464_io_enable; // @[RegFile.scala 66:20:@56226.4]
  wire  regs_465_clock; // @[RegFile.scala 66:20:@56240.4]
  wire  regs_465_reset; // @[RegFile.scala 66:20:@56240.4]
  wire [63:0] regs_465_io_in; // @[RegFile.scala 66:20:@56240.4]
  wire  regs_465_io_reset; // @[RegFile.scala 66:20:@56240.4]
  wire [63:0] regs_465_io_out; // @[RegFile.scala 66:20:@56240.4]
  wire  regs_465_io_enable; // @[RegFile.scala 66:20:@56240.4]
  wire  regs_466_clock; // @[RegFile.scala 66:20:@56254.4]
  wire  regs_466_reset; // @[RegFile.scala 66:20:@56254.4]
  wire [63:0] regs_466_io_in; // @[RegFile.scala 66:20:@56254.4]
  wire  regs_466_io_reset; // @[RegFile.scala 66:20:@56254.4]
  wire [63:0] regs_466_io_out; // @[RegFile.scala 66:20:@56254.4]
  wire  regs_466_io_enable; // @[RegFile.scala 66:20:@56254.4]
  wire  regs_467_clock; // @[RegFile.scala 66:20:@56268.4]
  wire  regs_467_reset; // @[RegFile.scala 66:20:@56268.4]
  wire [63:0] regs_467_io_in; // @[RegFile.scala 66:20:@56268.4]
  wire  regs_467_io_reset; // @[RegFile.scala 66:20:@56268.4]
  wire [63:0] regs_467_io_out; // @[RegFile.scala 66:20:@56268.4]
  wire  regs_467_io_enable; // @[RegFile.scala 66:20:@56268.4]
  wire  regs_468_clock; // @[RegFile.scala 66:20:@56282.4]
  wire  regs_468_reset; // @[RegFile.scala 66:20:@56282.4]
  wire [63:0] regs_468_io_in; // @[RegFile.scala 66:20:@56282.4]
  wire  regs_468_io_reset; // @[RegFile.scala 66:20:@56282.4]
  wire [63:0] regs_468_io_out; // @[RegFile.scala 66:20:@56282.4]
  wire  regs_468_io_enable; // @[RegFile.scala 66:20:@56282.4]
  wire  regs_469_clock; // @[RegFile.scala 66:20:@56296.4]
  wire  regs_469_reset; // @[RegFile.scala 66:20:@56296.4]
  wire [63:0] regs_469_io_in; // @[RegFile.scala 66:20:@56296.4]
  wire  regs_469_io_reset; // @[RegFile.scala 66:20:@56296.4]
  wire [63:0] regs_469_io_out; // @[RegFile.scala 66:20:@56296.4]
  wire  regs_469_io_enable; // @[RegFile.scala 66:20:@56296.4]
  wire  regs_470_clock; // @[RegFile.scala 66:20:@56310.4]
  wire  regs_470_reset; // @[RegFile.scala 66:20:@56310.4]
  wire [63:0] regs_470_io_in; // @[RegFile.scala 66:20:@56310.4]
  wire  regs_470_io_reset; // @[RegFile.scala 66:20:@56310.4]
  wire [63:0] regs_470_io_out; // @[RegFile.scala 66:20:@56310.4]
  wire  regs_470_io_enable; // @[RegFile.scala 66:20:@56310.4]
  wire  regs_471_clock; // @[RegFile.scala 66:20:@56324.4]
  wire  regs_471_reset; // @[RegFile.scala 66:20:@56324.4]
  wire [63:0] regs_471_io_in; // @[RegFile.scala 66:20:@56324.4]
  wire  regs_471_io_reset; // @[RegFile.scala 66:20:@56324.4]
  wire [63:0] regs_471_io_out; // @[RegFile.scala 66:20:@56324.4]
  wire  regs_471_io_enable; // @[RegFile.scala 66:20:@56324.4]
  wire  regs_472_clock; // @[RegFile.scala 66:20:@56338.4]
  wire  regs_472_reset; // @[RegFile.scala 66:20:@56338.4]
  wire [63:0] regs_472_io_in; // @[RegFile.scala 66:20:@56338.4]
  wire  regs_472_io_reset; // @[RegFile.scala 66:20:@56338.4]
  wire [63:0] regs_472_io_out; // @[RegFile.scala 66:20:@56338.4]
  wire  regs_472_io_enable; // @[RegFile.scala 66:20:@56338.4]
  wire  regs_473_clock; // @[RegFile.scala 66:20:@56352.4]
  wire  regs_473_reset; // @[RegFile.scala 66:20:@56352.4]
  wire [63:0] regs_473_io_in; // @[RegFile.scala 66:20:@56352.4]
  wire  regs_473_io_reset; // @[RegFile.scala 66:20:@56352.4]
  wire [63:0] regs_473_io_out; // @[RegFile.scala 66:20:@56352.4]
  wire  regs_473_io_enable; // @[RegFile.scala 66:20:@56352.4]
  wire  regs_474_clock; // @[RegFile.scala 66:20:@56366.4]
  wire  regs_474_reset; // @[RegFile.scala 66:20:@56366.4]
  wire [63:0] regs_474_io_in; // @[RegFile.scala 66:20:@56366.4]
  wire  regs_474_io_reset; // @[RegFile.scala 66:20:@56366.4]
  wire [63:0] regs_474_io_out; // @[RegFile.scala 66:20:@56366.4]
  wire  regs_474_io_enable; // @[RegFile.scala 66:20:@56366.4]
  wire  regs_475_clock; // @[RegFile.scala 66:20:@56380.4]
  wire  regs_475_reset; // @[RegFile.scala 66:20:@56380.4]
  wire [63:0] regs_475_io_in; // @[RegFile.scala 66:20:@56380.4]
  wire  regs_475_io_reset; // @[RegFile.scala 66:20:@56380.4]
  wire [63:0] regs_475_io_out; // @[RegFile.scala 66:20:@56380.4]
  wire  regs_475_io_enable; // @[RegFile.scala 66:20:@56380.4]
  wire  regs_476_clock; // @[RegFile.scala 66:20:@56394.4]
  wire  regs_476_reset; // @[RegFile.scala 66:20:@56394.4]
  wire [63:0] regs_476_io_in; // @[RegFile.scala 66:20:@56394.4]
  wire  regs_476_io_reset; // @[RegFile.scala 66:20:@56394.4]
  wire [63:0] regs_476_io_out; // @[RegFile.scala 66:20:@56394.4]
  wire  regs_476_io_enable; // @[RegFile.scala 66:20:@56394.4]
  wire  regs_477_clock; // @[RegFile.scala 66:20:@56408.4]
  wire  regs_477_reset; // @[RegFile.scala 66:20:@56408.4]
  wire [63:0] regs_477_io_in; // @[RegFile.scala 66:20:@56408.4]
  wire  regs_477_io_reset; // @[RegFile.scala 66:20:@56408.4]
  wire [63:0] regs_477_io_out; // @[RegFile.scala 66:20:@56408.4]
  wire  regs_477_io_enable; // @[RegFile.scala 66:20:@56408.4]
  wire  regs_478_clock; // @[RegFile.scala 66:20:@56422.4]
  wire  regs_478_reset; // @[RegFile.scala 66:20:@56422.4]
  wire [63:0] regs_478_io_in; // @[RegFile.scala 66:20:@56422.4]
  wire  regs_478_io_reset; // @[RegFile.scala 66:20:@56422.4]
  wire [63:0] regs_478_io_out; // @[RegFile.scala 66:20:@56422.4]
  wire  regs_478_io_enable; // @[RegFile.scala 66:20:@56422.4]
  wire  regs_479_clock; // @[RegFile.scala 66:20:@56436.4]
  wire  regs_479_reset; // @[RegFile.scala 66:20:@56436.4]
  wire [63:0] regs_479_io_in; // @[RegFile.scala 66:20:@56436.4]
  wire  regs_479_io_reset; // @[RegFile.scala 66:20:@56436.4]
  wire [63:0] regs_479_io_out; // @[RegFile.scala 66:20:@56436.4]
  wire  regs_479_io_enable; // @[RegFile.scala 66:20:@56436.4]
  wire  regs_480_clock; // @[RegFile.scala 66:20:@56450.4]
  wire  regs_480_reset; // @[RegFile.scala 66:20:@56450.4]
  wire [63:0] regs_480_io_in; // @[RegFile.scala 66:20:@56450.4]
  wire  regs_480_io_reset; // @[RegFile.scala 66:20:@56450.4]
  wire [63:0] regs_480_io_out; // @[RegFile.scala 66:20:@56450.4]
  wire  regs_480_io_enable; // @[RegFile.scala 66:20:@56450.4]
  wire  regs_481_clock; // @[RegFile.scala 66:20:@56464.4]
  wire  regs_481_reset; // @[RegFile.scala 66:20:@56464.4]
  wire [63:0] regs_481_io_in; // @[RegFile.scala 66:20:@56464.4]
  wire  regs_481_io_reset; // @[RegFile.scala 66:20:@56464.4]
  wire [63:0] regs_481_io_out; // @[RegFile.scala 66:20:@56464.4]
  wire  regs_481_io_enable; // @[RegFile.scala 66:20:@56464.4]
  wire  regs_482_clock; // @[RegFile.scala 66:20:@56478.4]
  wire  regs_482_reset; // @[RegFile.scala 66:20:@56478.4]
  wire [63:0] regs_482_io_in; // @[RegFile.scala 66:20:@56478.4]
  wire  regs_482_io_reset; // @[RegFile.scala 66:20:@56478.4]
  wire [63:0] regs_482_io_out; // @[RegFile.scala 66:20:@56478.4]
  wire  regs_482_io_enable; // @[RegFile.scala 66:20:@56478.4]
  wire  regs_483_clock; // @[RegFile.scala 66:20:@56492.4]
  wire  regs_483_reset; // @[RegFile.scala 66:20:@56492.4]
  wire [63:0] regs_483_io_in; // @[RegFile.scala 66:20:@56492.4]
  wire  regs_483_io_reset; // @[RegFile.scala 66:20:@56492.4]
  wire [63:0] regs_483_io_out; // @[RegFile.scala 66:20:@56492.4]
  wire  regs_483_io_enable; // @[RegFile.scala 66:20:@56492.4]
  wire  regs_484_clock; // @[RegFile.scala 66:20:@56506.4]
  wire  regs_484_reset; // @[RegFile.scala 66:20:@56506.4]
  wire [63:0] regs_484_io_in; // @[RegFile.scala 66:20:@56506.4]
  wire  regs_484_io_reset; // @[RegFile.scala 66:20:@56506.4]
  wire [63:0] regs_484_io_out; // @[RegFile.scala 66:20:@56506.4]
  wire  regs_484_io_enable; // @[RegFile.scala 66:20:@56506.4]
  wire  regs_485_clock; // @[RegFile.scala 66:20:@56520.4]
  wire  regs_485_reset; // @[RegFile.scala 66:20:@56520.4]
  wire [63:0] regs_485_io_in; // @[RegFile.scala 66:20:@56520.4]
  wire  regs_485_io_reset; // @[RegFile.scala 66:20:@56520.4]
  wire [63:0] regs_485_io_out; // @[RegFile.scala 66:20:@56520.4]
  wire  regs_485_io_enable; // @[RegFile.scala 66:20:@56520.4]
  wire  regs_486_clock; // @[RegFile.scala 66:20:@56534.4]
  wire  regs_486_reset; // @[RegFile.scala 66:20:@56534.4]
  wire [63:0] regs_486_io_in; // @[RegFile.scala 66:20:@56534.4]
  wire  regs_486_io_reset; // @[RegFile.scala 66:20:@56534.4]
  wire [63:0] regs_486_io_out; // @[RegFile.scala 66:20:@56534.4]
  wire  regs_486_io_enable; // @[RegFile.scala 66:20:@56534.4]
  wire  regs_487_clock; // @[RegFile.scala 66:20:@56548.4]
  wire  regs_487_reset; // @[RegFile.scala 66:20:@56548.4]
  wire [63:0] regs_487_io_in; // @[RegFile.scala 66:20:@56548.4]
  wire  regs_487_io_reset; // @[RegFile.scala 66:20:@56548.4]
  wire [63:0] regs_487_io_out; // @[RegFile.scala 66:20:@56548.4]
  wire  regs_487_io_enable; // @[RegFile.scala 66:20:@56548.4]
  wire  regs_488_clock; // @[RegFile.scala 66:20:@56562.4]
  wire  regs_488_reset; // @[RegFile.scala 66:20:@56562.4]
  wire [63:0] regs_488_io_in; // @[RegFile.scala 66:20:@56562.4]
  wire  regs_488_io_reset; // @[RegFile.scala 66:20:@56562.4]
  wire [63:0] regs_488_io_out; // @[RegFile.scala 66:20:@56562.4]
  wire  regs_488_io_enable; // @[RegFile.scala 66:20:@56562.4]
  wire  regs_489_clock; // @[RegFile.scala 66:20:@56576.4]
  wire  regs_489_reset; // @[RegFile.scala 66:20:@56576.4]
  wire [63:0] regs_489_io_in; // @[RegFile.scala 66:20:@56576.4]
  wire  regs_489_io_reset; // @[RegFile.scala 66:20:@56576.4]
  wire [63:0] regs_489_io_out; // @[RegFile.scala 66:20:@56576.4]
  wire  regs_489_io_enable; // @[RegFile.scala 66:20:@56576.4]
  wire  regs_490_clock; // @[RegFile.scala 66:20:@56590.4]
  wire  regs_490_reset; // @[RegFile.scala 66:20:@56590.4]
  wire [63:0] regs_490_io_in; // @[RegFile.scala 66:20:@56590.4]
  wire  regs_490_io_reset; // @[RegFile.scala 66:20:@56590.4]
  wire [63:0] regs_490_io_out; // @[RegFile.scala 66:20:@56590.4]
  wire  regs_490_io_enable; // @[RegFile.scala 66:20:@56590.4]
  wire  regs_491_clock; // @[RegFile.scala 66:20:@56604.4]
  wire  regs_491_reset; // @[RegFile.scala 66:20:@56604.4]
  wire [63:0] regs_491_io_in; // @[RegFile.scala 66:20:@56604.4]
  wire  regs_491_io_reset; // @[RegFile.scala 66:20:@56604.4]
  wire [63:0] regs_491_io_out; // @[RegFile.scala 66:20:@56604.4]
  wire  regs_491_io_enable; // @[RegFile.scala 66:20:@56604.4]
  wire  regs_492_clock; // @[RegFile.scala 66:20:@56618.4]
  wire  regs_492_reset; // @[RegFile.scala 66:20:@56618.4]
  wire [63:0] regs_492_io_in; // @[RegFile.scala 66:20:@56618.4]
  wire  regs_492_io_reset; // @[RegFile.scala 66:20:@56618.4]
  wire [63:0] regs_492_io_out; // @[RegFile.scala 66:20:@56618.4]
  wire  regs_492_io_enable; // @[RegFile.scala 66:20:@56618.4]
  wire  regs_493_clock; // @[RegFile.scala 66:20:@56632.4]
  wire  regs_493_reset; // @[RegFile.scala 66:20:@56632.4]
  wire [63:0] regs_493_io_in; // @[RegFile.scala 66:20:@56632.4]
  wire  regs_493_io_reset; // @[RegFile.scala 66:20:@56632.4]
  wire [63:0] regs_493_io_out; // @[RegFile.scala 66:20:@56632.4]
  wire  regs_493_io_enable; // @[RegFile.scala 66:20:@56632.4]
  wire  regs_494_clock; // @[RegFile.scala 66:20:@56646.4]
  wire  regs_494_reset; // @[RegFile.scala 66:20:@56646.4]
  wire [63:0] regs_494_io_in; // @[RegFile.scala 66:20:@56646.4]
  wire  regs_494_io_reset; // @[RegFile.scala 66:20:@56646.4]
  wire [63:0] regs_494_io_out; // @[RegFile.scala 66:20:@56646.4]
  wire  regs_494_io_enable; // @[RegFile.scala 66:20:@56646.4]
  wire  regs_495_clock; // @[RegFile.scala 66:20:@56660.4]
  wire  regs_495_reset; // @[RegFile.scala 66:20:@56660.4]
  wire [63:0] regs_495_io_in; // @[RegFile.scala 66:20:@56660.4]
  wire  regs_495_io_reset; // @[RegFile.scala 66:20:@56660.4]
  wire [63:0] regs_495_io_out; // @[RegFile.scala 66:20:@56660.4]
  wire  regs_495_io_enable; // @[RegFile.scala 66:20:@56660.4]
  wire  regs_496_clock; // @[RegFile.scala 66:20:@56674.4]
  wire  regs_496_reset; // @[RegFile.scala 66:20:@56674.4]
  wire [63:0] regs_496_io_in; // @[RegFile.scala 66:20:@56674.4]
  wire  regs_496_io_reset; // @[RegFile.scala 66:20:@56674.4]
  wire [63:0] regs_496_io_out; // @[RegFile.scala 66:20:@56674.4]
  wire  regs_496_io_enable; // @[RegFile.scala 66:20:@56674.4]
  wire  regs_497_clock; // @[RegFile.scala 66:20:@56688.4]
  wire  regs_497_reset; // @[RegFile.scala 66:20:@56688.4]
  wire [63:0] regs_497_io_in; // @[RegFile.scala 66:20:@56688.4]
  wire  regs_497_io_reset; // @[RegFile.scala 66:20:@56688.4]
  wire [63:0] regs_497_io_out; // @[RegFile.scala 66:20:@56688.4]
  wire  regs_497_io_enable; // @[RegFile.scala 66:20:@56688.4]
  wire  regs_498_clock; // @[RegFile.scala 66:20:@56702.4]
  wire  regs_498_reset; // @[RegFile.scala 66:20:@56702.4]
  wire [63:0] regs_498_io_in; // @[RegFile.scala 66:20:@56702.4]
  wire  regs_498_io_reset; // @[RegFile.scala 66:20:@56702.4]
  wire [63:0] regs_498_io_out; // @[RegFile.scala 66:20:@56702.4]
  wire  regs_498_io_enable; // @[RegFile.scala 66:20:@56702.4]
  wire  regs_499_clock; // @[RegFile.scala 66:20:@56716.4]
  wire  regs_499_reset; // @[RegFile.scala 66:20:@56716.4]
  wire [63:0] regs_499_io_in; // @[RegFile.scala 66:20:@56716.4]
  wire  regs_499_io_reset; // @[RegFile.scala 66:20:@56716.4]
  wire [63:0] regs_499_io_out; // @[RegFile.scala 66:20:@56716.4]
  wire  regs_499_io_enable; // @[RegFile.scala 66:20:@56716.4]
  wire  regs_500_clock; // @[RegFile.scala 66:20:@56730.4]
  wire  regs_500_reset; // @[RegFile.scala 66:20:@56730.4]
  wire [63:0] regs_500_io_in; // @[RegFile.scala 66:20:@56730.4]
  wire  regs_500_io_reset; // @[RegFile.scala 66:20:@56730.4]
  wire [63:0] regs_500_io_out; // @[RegFile.scala 66:20:@56730.4]
  wire  regs_500_io_enable; // @[RegFile.scala 66:20:@56730.4]
  wire  regs_501_clock; // @[RegFile.scala 66:20:@56744.4]
  wire  regs_501_reset; // @[RegFile.scala 66:20:@56744.4]
  wire [63:0] regs_501_io_in; // @[RegFile.scala 66:20:@56744.4]
  wire  regs_501_io_reset; // @[RegFile.scala 66:20:@56744.4]
  wire [63:0] regs_501_io_out; // @[RegFile.scala 66:20:@56744.4]
  wire  regs_501_io_enable; // @[RegFile.scala 66:20:@56744.4]
  wire  regs_502_clock; // @[RegFile.scala 66:20:@56758.4]
  wire  regs_502_reset; // @[RegFile.scala 66:20:@56758.4]
  wire [63:0] regs_502_io_in; // @[RegFile.scala 66:20:@56758.4]
  wire  regs_502_io_reset; // @[RegFile.scala 66:20:@56758.4]
  wire [63:0] regs_502_io_out; // @[RegFile.scala 66:20:@56758.4]
  wire  regs_502_io_enable; // @[RegFile.scala 66:20:@56758.4]
  wire  regs_503_clock; // @[RegFile.scala 66:20:@56772.4]
  wire  regs_503_reset; // @[RegFile.scala 66:20:@56772.4]
  wire [63:0] regs_503_io_in; // @[RegFile.scala 66:20:@56772.4]
  wire  regs_503_io_reset; // @[RegFile.scala 66:20:@56772.4]
  wire [63:0] regs_503_io_out; // @[RegFile.scala 66:20:@56772.4]
  wire  regs_503_io_enable; // @[RegFile.scala 66:20:@56772.4]
  wire  regs_504_clock; // @[RegFile.scala 66:20:@56786.4]
  wire  regs_504_reset; // @[RegFile.scala 66:20:@56786.4]
  wire [63:0] regs_504_io_in; // @[RegFile.scala 66:20:@56786.4]
  wire  regs_504_io_reset; // @[RegFile.scala 66:20:@56786.4]
  wire [63:0] regs_504_io_out; // @[RegFile.scala 66:20:@56786.4]
  wire  regs_504_io_enable; // @[RegFile.scala 66:20:@56786.4]
  wire  regs_505_clock; // @[RegFile.scala 66:20:@56800.4]
  wire  regs_505_reset; // @[RegFile.scala 66:20:@56800.4]
  wire [63:0] regs_505_io_in; // @[RegFile.scala 66:20:@56800.4]
  wire  regs_505_io_reset; // @[RegFile.scala 66:20:@56800.4]
  wire [63:0] regs_505_io_out; // @[RegFile.scala 66:20:@56800.4]
  wire  regs_505_io_enable; // @[RegFile.scala 66:20:@56800.4]
  wire  regs_506_clock; // @[RegFile.scala 66:20:@56814.4]
  wire  regs_506_reset; // @[RegFile.scala 66:20:@56814.4]
  wire [63:0] regs_506_io_in; // @[RegFile.scala 66:20:@56814.4]
  wire  regs_506_io_reset; // @[RegFile.scala 66:20:@56814.4]
  wire [63:0] regs_506_io_out; // @[RegFile.scala 66:20:@56814.4]
  wire  regs_506_io_enable; // @[RegFile.scala 66:20:@56814.4]
  wire  regs_507_clock; // @[RegFile.scala 66:20:@56828.4]
  wire  regs_507_reset; // @[RegFile.scala 66:20:@56828.4]
  wire [63:0] regs_507_io_in; // @[RegFile.scala 66:20:@56828.4]
  wire  regs_507_io_reset; // @[RegFile.scala 66:20:@56828.4]
  wire [63:0] regs_507_io_out; // @[RegFile.scala 66:20:@56828.4]
  wire  regs_507_io_enable; // @[RegFile.scala 66:20:@56828.4]
  wire  regs_508_clock; // @[RegFile.scala 66:20:@56842.4]
  wire  regs_508_reset; // @[RegFile.scala 66:20:@56842.4]
  wire [63:0] regs_508_io_in; // @[RegFile.scala 66:20:@56842.4]
  wire  regs_508_io_reset; // @[RegFile.scala 66:20:@56842.4]
  wire [63:0] regs_508_io_out; // @[RegFile.scala 66:20:@56842.4]
  wire  regs_508_io_enable; // @[RegFile.scala 66:20:@56842.4]
  wire  regs_509_clock; // @[RegFile.scala 66:20:@56856.4]
  wire  regs_509_reset; // @[RegFile.scala 66:20:@56856.4]
  wire [63:0] regs_509_io_in; // @[RegFile.scala 66:20:@56856.4]
  wire  regs_509_io_reset; // @[RegFile.scala 66:20:@56856.4]
  wire [63:0] regs_509_io_out; // @[RegFile.scala 66:20:@56856.4]
  wire  regs_509_io_enable; // @[RegFile.scala 66:20:@56856.4]
  wire  regs_510_clock; // @[RegFile.scala 66:20:@56870.4]
  wire  regs_510_reset; // @[RegFile.scala 66:20:@56870.4]
  wire [63:0] regs_510_io_in; // @[RegFile.scala 66:20:@56870.4]
  wire  regs_510_io_reset; // @[RegFile.scala 66:20:@56870.4]
  wire [63:0] regs_510_io_out; // @[RegFile.scala 66:20:@56870.4]
  wire  regs_510_io_enable; // @[RegFile.scala 66:20:@56870.4]
  wire  regs_511_clock; // @[RegFile.scala 66:20:@56884.4]
  wire  regs_511_reset; // @[RegFile.scala 66:20:@56884.4]
  wire [63:0] regs_511_io_in; // @[RegFile.scala 66:20:@56884.4]
  wire  regs_511_io_reset; // @[RegFile.scala 66:20:@56884.4]
  wire [63:0] regs_511_io_out; // @[RegFile.scala 66:20:@56884.4]
  wire  regs_511_io_enable; // @[RegFile.scala 66:20:@56884.4]
  wire  regs_512_clock; // @[RegFile.scala 66:20:@56898.4]
  wire  regs_512_reset; // @[RegFile.scala 66:20:@56898.4]
  wire [63:0] regs_512_io_in; // @[RegFile.scala 66:20:@56898.4]
  wire  regs_512_io_reset; // @[RegFile.scala 66:20:@56898.4]
  wire [63:0] regs_512_io_out; // @[RegFile.scala 66:20:@56898.4]
  wire  regs_512_io_enable; // @[RegFile.scala 66:20:@56898.4]
  wire  regs_513_clock; // @[RegFile.scala 66:20:@56912.4]
  wire  regs_513_reset; // @[RegFile.scala 66:20:@56912.4]
  wire [63:0] regs_513_io_in; // @[RegFile.scala 66:20:@56912.4]
  wire  regs_513_io_reset; // @[RegFile.scala 66:20:@56912.4]
  wire [63:0] regs_513_io_out; // @[RegFile.scala 66:20:@56912.4]
  wire  regs_513_io_enable; // @[RegFile.scala 66:20:@56912.4]
  wire  regs_514_clock; // @[RegFile.scala 66:20:@56926.4]
  wire  regs_514_reset; // @[RegFile.scala 66:20:@56926.4]
  wire [63:0] regs_514_io_in; // @[RegFile.scala 66:20:@56926.4]
  wire  regs_514_io_reset; // @[RegFile.scala 66:20:@56926.4]
  wire [63:0] regs_514_io_out; // @[RegFile.scala 66:20:@56926.4]
  wire  regs_514_io_enable; // @[RegFile.scala 66:20:@56926.4]
  wire  regs_515_clock; // @[RegFile.scala 66:20:@56940.4]
  wire  regs_515_reset; // @[RegFile.scala 66:20:@56940.4]
  wire [63:0] regs_515_io_in; // @[RegFile.scala 66:20:@56940.4]
  wire  regs_515_io_reset; // @[RegFile.scala 66:20:@56940.4]
  wire [63:0] regs_515_io_out; // @[RegFile.scala 66:20:@56940.4]
  wire  regs_515_io_enable; // @[RegFile.scala 66:20:@56940.4]
  wire  regs_516_clock; // @[RegFile.scala 66:20:@56954.4]
  wire  regs_516_reset; // @[RegFile.scala 66:20:@56954.4]
  wire [63:0] regs_516_io_in; // @[RegFile.scala 66:20:@56954.4]
  wire  regs_516_io_reset; // @[RegFile.scala 66:20:@56954.4]
  wire [63:0] regs_516_io_out; // @[RegFile.scala 66:20:@56954.4]
  wire  regs_516_io_enable; // @[RegFile.scala 66:20:@56954.4]
  wire  regs_517_clock; // @[RegFile.scala 66:20:@56968.4]
  wire  regs_517_reset; // @[RegFile.scala 66:20:@56968.4]
  wire [63:0] regs_517_io_in; // @[RegFile.scala 66:20:@56968.4]
  wire  regs_517_io_reset; // @[RegFile.scala 66:20:@56968.4]
  wire [63:0] regs_517_io_out; // @[RegFile.scala 66:20:@56968.4]
  wire  regs_517_io_enable; // @[RegFile.scala 66:20:@56968.4]
  wire [63:0] rport_io_ins_0; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_1; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_2; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_3; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_4; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_5; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_6; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_7; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_8; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_9; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_10; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_11; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_12; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_13; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_14; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_15; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_16; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_17; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_18; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_19; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_20; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_21; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_22; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_23; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_24; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_25; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_26; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_27; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_28; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_29; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_30; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_31; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_32; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_33; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_34; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_35; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_36; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_37; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_38; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_39; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_40; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_41; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_42; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_43; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_44; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_45; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_46; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_47; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_48; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_49; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_50; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_51; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_52; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_53; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_54; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_55; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_56; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_57; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_58; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_59; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_60; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_61; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_62; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_63; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_64; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_65; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_66; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_67; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_68; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_69; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_70; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_71; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_72; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_73; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_74; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_75; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_76; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_77; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_78; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_79; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_80; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_81; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_82; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_83; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_84; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_85; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_86; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_87; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_88; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_89; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_90; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_91; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_92; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_93; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_94; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_95; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_96; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_97; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_98; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_99; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_100; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_101; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_102; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_103; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_104; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_105; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_106; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_107; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_108; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_109; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_110; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_111; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_112; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_113; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_114; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_115; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_116; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_117; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_118; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_119; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_120; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_121; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_122; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_123; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_124; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_125; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_126; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_127; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_128; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_129; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_130; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_131; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_132; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_133; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_134; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_135; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_136; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_137; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_138; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_139; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_140; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_141; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_142; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_143; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_144; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_145; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_146; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_147; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_148; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_149; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_150; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_151; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_152; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_153; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_154; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_155; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_156; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_157; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_158; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_159; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_160; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_161; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_162; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_163; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_164; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_165; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_166; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_167; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_168; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_169; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_170; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_171; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_172; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_173; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_174; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_175; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_176; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_177; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_178; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_179; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_180; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_181; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_182; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_183; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_184; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_185; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_186; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_187; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_188; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_189; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_190; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_191; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_192; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_193; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_194; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_195; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_196; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_197; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_198; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_199; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_200; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_201; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_202; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_203; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_204; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_205; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_206; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_207; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_208; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_209; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_210; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_211; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_212; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_213; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_214; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_215; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_216; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_217; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_218; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_219; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_220; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_221; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_222; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_223; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_224; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_225; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_226; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_227; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_228; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_229; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_230; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_231; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_232; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_233; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_234; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_235; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_236; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_237; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_238; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_239; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_240; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_241; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_242; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_243; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_244; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_245; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_246; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_247; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_248; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_249; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_250; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_251; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_252; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_253; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_254; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_255; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_256; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_257; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_258; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_259; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_260; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_261; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_262; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_263; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_264; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_265; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_266; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_267; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_268; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_269; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_270; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_271; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_272; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_273; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_274; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_275; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_276; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_277; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_278; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_279; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_280; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_281; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_282; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_283; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_284; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_285; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_286; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_287; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_288; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_289; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_290; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_291; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_292; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_293; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_294; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_295; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_296; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_297; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_298; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_299; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_300; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_301; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_302; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_303; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_304; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_305; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_306; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_307; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_308; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_309; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_310; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_311; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_312; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_313; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_314; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_315; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_316; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_317; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_318; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_319; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_320; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_321; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_322; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_323; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_324; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_325; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_326; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_327; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_328; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_329; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_330; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_331; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_332; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_333; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_334; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_335; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_336; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_337; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_338; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_339; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_340; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_341; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_342; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_343; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_344; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_345; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_346; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_347; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_348; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_349; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_350; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_351; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_352; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_353; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_354; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_355; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_356; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_357; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_358; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_359; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_360; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_361; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_362; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_363; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_364; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_365; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_366; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_367; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_368; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_369; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_370; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_371; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_372; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_373; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_374; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_375; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_376; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_377; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_378; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_379; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_380; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_381; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_382; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_383; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_384; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_385; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_386; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_387; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_388; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_389; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_390; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_391; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_392; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_393; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_394; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_395; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_396; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_397; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_398; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_399; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_400; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_401; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_402; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_403; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_404; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_405; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_406; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_407; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_408; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_409; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_410; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_411; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_412; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_413; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_414; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_415; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_416; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_417; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_418; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_419; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_420; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_421; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_422; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_423; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_424; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_425; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_426; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_427; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_428; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_429; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_430; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_431; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_432; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_433; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_434; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_435; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_436; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_437; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_438; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_439; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_440; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_441; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_442; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_443; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_444; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_445; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_446; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_447; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_448; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_449; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_450; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_451; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_452; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_453; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_454; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_455; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_456; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_457; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_458; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_459; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_460; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_461; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_462; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_463; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_464; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_465; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_466; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_467; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_468; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_469; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_470; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_471; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_472; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_473; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_474; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_475; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_476; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_477; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_478; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_479; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_480; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_481; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_482; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_483; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_484; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_485; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_486; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_487; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_488; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_489; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_490; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_491; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_492; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_493; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_494; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_495; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_496; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_497; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_498; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_499; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_500; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_501; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_502; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_503; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_504; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_505; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_506; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_507; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_508; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_509; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_510; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_511; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_512; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_513; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_514; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_515; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_516; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_ins_517; // @[RegFile.scala 95:21:@56982.4]
  wire [9:0] rport_io_sel; // @[RegFile.scala 95:21:@56982.4]
  wire [63:0] rport_io_out; // @[RegFile.scala 95:21:@56982.4]
  wire  _T_3166; // @[RegFile.scala 80:42:@49732.4]
  wire  _T_3172; // @[RegFile.scala 68:46:@49744.4]
  wire  _T_3173; // @[RegFile.scala 68:34:@49745.4]
  wire  _T_3186; // @[RegFile.scala 80:42:@49763.4]
  wire  _T_3192; // @[RegFile.scala 74:80:@49775.4]
  wire  _T_3193; // @[RegFile.scala 74:68:@49776.4]
  wire  _T_3199; // @[RegFile.scala 74:80:@49789.4]
  wire  _T_3200; // @[RegFile.scala 74:68:@49790.4]
  wire  _T_3206; // @[RegFile.scala 74:80:@49803.4]
  wire  _T_3207; // @[RegFile.scala 74:68:@49804.4]
  wire  _T_3213; // @[RegFile.scala 74:80:@49817.4]
  wire  _T_3214; // @[RegFile.scala 74:68:@49818.4]
  wire  _T_3220; // @[RegFile.scala 74:80:@49831.4]
  wire  _T_3221; // @[RegFile.scala 74:68:@49832.4]
  wire  _T_3227; // @[RegFile.scala 74:80:@49845.4]
  wire  _T_3228; // @[RegFile.scala 74:68:@49846.4]
  wire  _T_3234; // @[RegFile.scala 74:80:@49859.4]
  wire  _T_3235; // @[RegFile.scala 74:68:@49860.4]
  wire  _T_3241; // @[RegFile.scala 74:80:@49873.4]
  wire  _T_3242; // @[RegFile.scala 74:68:@49874.4]
  wire  _T_3248; // @[RegFile.scala 74:80:@49887.4]
  wire  _T_3249; // @[RegFile.scala 74:68:@49888.4]
  wire  _T_3255; // @[RegFile.scala 74:80:@49901.4]
  wire  _T_3256; // @[RegFile.scala 74:68:@49902.4]
  wire  _T_3262; // @[RegFile.scala 74:80:@49915.4]
  wire  _T_3263; // @[RegFile.scala 74:68:@49916.4]
  wire  _T_3269; // @[RegFile.scala 74:80:@49929.4]
  wire  _T_3270; // @[RegFile.scala 74:68:@49930.4]
  wire  _T_3276; // @[RegFile.scala 74:80:@49943.4]
  wire  _T_3277; // @[RegFile.scala 74:68:@49944.4]
  wire  _T_3283; // @[RegFile.scala 74:80:@49957.4]
  wire  _T_3284; // @[RegFile.scala 74:68:@49958.4]
  wire  _T_3290; // @[RegFile.scala 74:80:@49971.4]
  wire  _T_3291; // @[RegFile.scala 74:68:@49972.4]
  wire  _T_3297; // @[RegFile.scala 74:80:@49985.4]
  wire  _T_3298; // @[RegFile.scala 74:68:@49986.4]
  FringeFF regs_0 ( // @[RegFile.scala 66:20:@49729.4]
    .clock(regs_0_clock),
    .reset(regs_0_reset),
    .io_in(regs_0_io_in),
    .io_reset(regs_0_io_reset),
    .io_out(regs_0_io_out),
    .io_enable(regs_0_io_enable)
  );
  FringeFF regs_1 ( // @[RegFile.scala 66:20:@49741.4]
    .clock(regs_1_clock),
    .reset(regs_1_reset),
    .io_in(regs_1_io_in),
    .io_reset(regs_1_io_reset),
    .io_out(regs_1_io_out),
    .io_enable(regs_1_io_enable)
  );
  FringeFF regs_2 ( // @[RegFile.scala 66:20:@49760.4]
    .clock(regs_2_clock),
    .reset(regs_2_reset),
    .io_in(regs_2_io_in),
    .io_reset(regs_2_io_reset),
    .io_out(regs_2_io_out),
    .io_enable(regs_2_io_enable)
  );
  FringeFF regs_3 ( // @[RegFile.scala 66:20:@49772.4]
    .clock(regs_3_clock),
    .reset(regs_3_reset),
    .io_in(regs_3_io_in),
    .io_reset(regs_3_io_reset),
    .io_out(regs_3_io_out),
    .io_enable(regs_3_io_enable)
  );
  FringeFF regs_4 ( // @[RegFile.scala 66:20:@49786.4]
    .clock(regs_4_clock),
    .reset(regs_4_reset),
    .io_in(regs_4_io_in),
    .io_reset(regs_4_io_reset),
    .io_out(regs_4_io_out),
    .io_enable(regs_4_io_enable)
  );
  FringeFF regs_5 ( // @[RegFile.scala 66:20:@49800.4]
    .clock(regs_5_clock),
    .reset(regs_5_reset),
    .io_in(regs_5_io_in),
    .io_reset(regs_5_io_reset),
    .io_out(regs_5_io_out),
    .io_enable(regs_5_io_enable)
  );
  FringeFF regs_6 ( // @[RegFile.scala 66:20:@49814.4]
    .clock(regs_6_clock),
    .reset(regs_6_reset),
    .io_in(regs_6_io_in),
    .io_reset(regs_6_io_reset),
    .io_out(regs_6_io_out),
    .io_enable(regs_6_io_enable)
  );
  FringeFF regs_7 ( // @[RegFile.scala 66:20:@49828.4]
    .clock(regs_7_clock),
    .reset(regs_7_reset),
    .io_in(regs_7_io_in),
    .io_reset(regs_7_io_reset),
    .io_out(regs_7_io_out),
    .io_enable(regs_7_io_enable)
  );
  FringeFF regs_8 ( // @[RegFile.scala 66:20:@49842.4]
    .clock(regs_8_clock),
    .reset(regs_8_reset),
    .io_in(regs_8_io_in),
    .io_reset(regs_8_io_reset),
    .io_out(regs_8_io_out),
    .io_enable(regs_8_io_enable)
  );
  FringeFF regs_9 ( // @[RegFile.scala 66:20:@49856.4]
    .clock(regs_9_clock),
    .reset(regs_9_reset),
    .io_in(regs_9_io_in),
    .io_reset(regs_9_io_reset),
    .io_out(regs_9_io_out),
    .io_enable(regs_9_io_enable)
  );
  FringeFF regs_10 ( // @[RegFile.scala 66:20:@49870.4]
    .clock(regs_10_clock),
    .reset(regs_10_reset),
    .io_in(regs_10_io_in),
    .io_reset(regs_10_io_reset),
    .io_out(regs_10_io_out),
    .io_enable(regs_10_io_enable)
  );
  FringeFF regs_11 ( // @[RegFile.scala 66:20:@49884.4]
    .clock(regs_11_clock),
    .reset(regs_11_reset),
    .io_in(regs_11_io_in),
    .io_reset(regs_11_io_reset),
    .io_out(regs_11_io_out),
    .io_enable(regs_11_io_enable)
  );
  FringeFF regs_12 ( // @[RegFile.scala 66:20:@49898.4]
    .clock(regs_12_clock),
    .reset(regs_12_reset),
    .io_in(regs_12_io_in),
    .io_reset(regs_12_io_reset),
    .io_out(regs_12_io_out),
    .io_enable(regs_12_io_enable)
  );
  FringeFF regs_13 ( // @[RegFile.scala 66:20:@49912.4]
    .clock(regs_13_clock),
    .reset(regs_13_reset),
    .io_in(regs_13_io_in),
    .io_reset(regs_13_io_reset),
    .io_out(regs_13_io_out),
    .io_enable(regs_13_io_enable)
  );
  FringeFF regs_14 ( // @[RegFile.scala 66:20:@49926.4]
    .clock(regs_14_clock),
    .reset(regs_14_reset),
    .io_in(regs_14_io_in),
    .io_reset(regs_14_io_reset),
    .io_out(regs_14_io_out),
    .io_enable(regs_14_io_enable)
  );
  FringeFF regs_15 ( // @[RegFile.scala 66:20:@49940.4]
    .clock(regs_15_clock),
    .reset(regs_15_reset),
    .io_in(regs_15_io_in),
    .io_reset(regs_15_io_reset),
    .io_out(regs_15_io_out),
    .io_enable(regs_15_io_enable)
  );
  FringeFF regs_16 ( // @[RegFile.scala 66:20:@49954.4]
    .clock(regs_16_clock),
    .reset(regs_16_reset),
    .io_in(regs_16_io_in),
    .io_reset(regs_16_io_reset),
    .io_out(regs_16_io_out),
    .io_enable(regs_16_io_enable)
  );
  FringeFF regs_17 ( // @[RegFile.scala 66:20:@49968.4]
    .clock(regs_17_clock),
    .reset(regs_17_reset),
    .io_in(regs_17_io_in),
    .io_reset(regs_17_io_reset),
    .io_out(regs_17_io_out),
    .io_enable(regs_17_io_enable)
  );
  FringeFF regs_18 ( // @[RegFile.scala 66:20:@49982.4]
    .clock(regs_18_clock),
    .reset(regs_18_reset),
    .io_in(regs_18_io_in),
    .io_reset(regs_18_io_reset),
    .io_out(regs_18_io_out),
    .io_enable(regs_18_io_enable)
  );
  FringeFF regs_19 ( // @[RegFile.scala 66:20:@49996.4]
    .clock(regs_19_clock),
    .reset(regs_19_reset),
    .io_in(regs_19_io_in),
    .io_reset(regs_19_io_reset),
    .io_out(regs_19_io_out),
    .io_enable(regs_19_io_enable)
  );
  FringeFF regs_20 ( // @[RegFile.scala 66:20:@50010.4]
    .clock(regs_20_clock),
    .reset(regs_20_reset),
    .io_in(regs_20_io_in),
    .io_reset(regs_20_io_reset),
    .io_out(regs_20_io_out),
    .io_enable(regs_20_io_enable)
  );
  FringeFF regs_21 ( // @[RegFile.scala 66:20:@50024.4]
    .clock(regs_21_clock),
    .reset(regs_21_reset),
    .io_in(regs_21_io_in),
    .io_reset(regs_21_io_reset),
    .io_out(regs_21_io_out),
    .io_enable(regs_21_io_enable)
  );
  FringeFF regs_22 ( // @[RegFile.scala 66:20:@50038.4]
    .clock(regs_22_clock),
    .reset(regs_22_reset),
    .io_in(regs_22_io_in),
    .io_reset(regs_22_io_reset),
    .io_out(regs_22_io_out),
    .io_enable(regs_22_io_enable)
  );
  FringeFF regs_23 ( // @[RegFile.scala 66:20:@50052.4]
    .clock(regs_23_clock),
    .reset(regs_23_reset),
    .io_in(regs_23_io_in),
    .io_reset(regs_23_io_reset),
    .io_out(regs_23_io_out),
    .io_enable(regs_23_io_enable)
  );
  FringeFF regs_24 ( // @[RegFile.scala 66:20:@50066.4]
    .clock(regs_24_clock),
    .reset(regs_24_reset),
    .io_in(regs_24_io_in),
    .io_reset(regs_24_io_reset),
    .io_out(regs_24_io_out),
    .io_enable(regs_24_io_enable)
  );
  FringeFF regs_25 ( // @[RegFile.scala 66:20:@50080.4]
    .clock(regs_25_clock),
    .reset(regs_25_reset),
    .io_in(regs_25_io_in),
    .io_reset(regs_25_io_reset),
    .io_out(regs_25_io_out),
    .io_enable(regs_25_io_enable)
  );
  FringeFF regs_26 ( // @[RegFile.scala 66:20:@50094.4]
    .clock(regs_26_clock),
    .reset(regs_26_reset),
    .io_in(regs_26_io_in),
    .io_reset(regs_26_io_reset),
    .io_out(regs_26_io_out),
    .io_enable(regs_26_io_enable)
  );
  FringeFF regs_27 ( // @[RegFile.scala 66:20:@50108.4]
    .clock(regs_27_clock),
    .reset(regs_27_reset),
    .io_in(regs_27_io_in),
    .io_reset(regs_27_io_reset),
    .io_out(regs_27_io_out),
    .io_enable(regs_27_io_enable)
  );
  FringeFF regs_28 ( // @[RegFile.scala 66:20:@50122.4]
    .clock(regs_28_clock),
    .reset(regs_28_reset),
    .io_in(regs_28_io_in),
    .io_reset(regs_28_io_reset),
    .io_out(regs_28_io_out),
    .io_enable(regs_28_io_enable)
  );
  FringeFF regs_29 ( // @[RegFile.scala 66:20:@50136.4]
    .clock(regs_29_clock),
    .reset(regs_29_reset),
    .io_in(regs_29_io_in),
    .io_reset(regs_29_io_reset),
    .io_out(regs_29_io_out),
    .io_enable(regs_29_io_enable)
  );
  FringeFF regs_30 ( // @[RegFile.scala 66:20:@50150.4]
    .clock(regs_30_clock),
    .reset(regs_30_reset),
    .io_in(regs_30_io_in),
    .io_reset(regs_30_io_reset),
    .io_out(regs_30_io_out),
    .io_enable(regs_30_io_enable)
  );
  FringeFF regs_31 ( // @[RegFile.scala 66:20:@50164.4]
    .clock(regs_31_clock),
    .reset(regs_31_reset),
    .io_in(regs_31_io_in),
    .io_reset(regs_31_io_reset),
    .io_out(regs_31_io_out),
    .io_enable(regs_31_io_enable)
  );
  FringeFF regs_32 ( // @[RegFile.scala 66:20:@50178.4]
    .clock(regs_32_clock),
    .reset(regs_32_reset),
    .io_in(regs_32_io_in),
    .io_reset(regs_32_io_reset),
    .io_out(regs_32_io_out),
    .io_enable(regs_32_io_enable)
  );
  FringeFF regs_33 ( // @[RegFile.scala 66:20:@50192.4]
    .clock(regs_33_clock),
    .reset(regs_33_reset),
    .io_in(regs_33_io_in),
    .io_reset(regs_33_io_reset),
    .io_out(regs_33_io_out),
    .io_enable(regs_33_io_enable)
  );
  FringeFF regs_34 ( // @[RegFile.scala 66:20:@50206.4]
    .clock(regs_34_clock),
    .reset(regs_34_reset),
    .io_in(regs_34_io_in),
    .io_reset(regs_34_io_reset),
    .io_out(regs_34_io_out),
    .io_enable(regs_34_io_enable)
  );
  FringeFF regs_35 ( // @[RegFile.scala 66:20:@50220.4]
    .clock(regs_35_clock),
    .reset(regs_35_reset),
    .io_in(regs_35_io_in),
    .io_reset(regs_35_io_reset),
    .io_out(regs_35_io_out),
    .io_enable(regs_35_io_enable)
  );
  FringeFF regs_36 ( // @[RegFile.scala 66:20:@50234.4]
    .clock(regs_36_clock),
    .reset(regs_36_reset),
    .io_in(regs_36_io_in),
    .io_reset(regs_36_io_reset),
    .io_out(regs_36_io_out),
    .io_enable(regs_36_io_enable)
  );
  FringeFF regs_37 ( // @[RegFile.scala 66:20:@50248.4]
    .clock(regs_37_clock),
    .reset(regs_37_reset),
    .io_in(regs_37_io_in),
    .io_reset(regs_37_io_reset),
    .io_out(regs_37_io_out),
    .io_enable(regs_37_io_enable)
  );
  FringeFF regs_38 ( // @[RegFile.scala 66:20:@50262.4]
    .clock(regs_38_clock),
    .reset(regs_38_reset),
    .io_in(regs_38_io_in),
    .io_reset(regs_38_io_reset),
    .io_out(regs_38_io_out),
    .io_enable(regs_38_io_enable)
  );
  FringeFF regs_39 ( // @[RegFile.scala 66:20:@50276.4]
    .clock(regs_39_clock),
    .reset(regs_39_reset),
    .io_in(regs_39_io_in),
    .io_reset(regs_39_io_reset),
    .io_out(regs_39_io_out),
    .io_enable(regs_39_io_enable)
  );
  FringeFF regs_40 ( // @[RegFile.scala 66:20:@50290.4]
    .clock(regs_40_clock),
    .reset(regs_40_reset),
    .io_in(regs_40_io_in),
    .io_reset(regs_40_io_reset),
    .io_out(regs_40_io_out),
    .io_enable(regs_40_io_enable)
  );
  FringeFF regs_41 ( // @[RegFile.scala 66:20:@50304.4]
    .clock(regs_41_clock),
    .reset(regs_41_reset),
    .io_in(regs_41_io_in),
    .io_reset(regs_41_io_reset),
    .io_out(regs_41_io_out),
    .io_enable(regs_41_io_enable)
  );
  FringeFF regs_42 ( // @[RegFile.scala 66:20:@50318.4]
    .clock(regs_42_clock),
    .reset(regs_42_reset),
    .io_in(regs_42_io_in),
    .io_reset(regs_42_io_reset),
    .io_out(regs_42_io_out),
    .io_enable(regs_42_io_enable)
  );
  FringeFF regs_43 ( // @[RegFile.scala 66:20:@50332.4]
    .clock(regs_43_clock),
    .reset(regs_43_reset),
    .io_in(regs_43_io_in),
    .io_reset(regs_43_io_reset),
    .io_out(regs_43_io_out),
    .io_enable(regs_43_io_enable)
  );
  FringeFF regs_44 ( // @[RegFile.scala 66:20:@50346.4]
    .clock(regs_44_clock),
    .reset(regs_44_reset),
    .io_in(regs_44_io_in),
    .io_reset(regs_44_io_reset),
    .io_out(regs_44_io_out),
    .io_enable(regs_44_io_enable)
  );
  FringeFF regs_45 ( // @[RegFile.scala 66:20:@50360.4]
    .clock(regs_45_clock),
    .reset(regs_45_reset),
    .io_in(regs_45_io_in),
    .io_reset(regs_45_io_reset),
    .io_out(regs_45_io_out),
    .io_enable(regs_45_io_enable)
  );
  FringeFF regs_46 ( // @[RegFile.scala 66:20:@50374.4]
    .clock(regs_46_clock),
    .reset(regs_46_reset),
    .io_in(regs_46_io_in),
    .io_reset(regs_46_io_reset),
    .io_out(regs_46_io_out),
    .io_enable(regs_46_io_enable)
  );
  FringeFF regs_47 ( // @[RegFile.scala 66:20:@50388.4]
    .clock(regs_47_clock),
    .reset(regs_47_reset),
    .io_in(regs_47_io_in),
    .io_reset(regs_47_io_reset),
    .io_out(regs_47_io_out),
    .io_enable(regs_47_io_enable)
  );
  FringeFF regs_48 ( // @[RegFile.scala 66:20:@50402.4]
    .clock(regs_48_clock),
    .reset(regs_48_reset),
    .io_in(regs_48_io_in),
    .io_reset(regs_48_io_reset),
    .io_out(regs_48_io_out),
    .io_enable(regs_48_io_enable)
  );
  FringeFF regs_49 ( // @[RegFile.scala 66:20:@50416.4]
    .clock(regs_49_clock),
    .reset(regs_49_reset),
    .io_in(regs_49_io_in),
    .io_reset(regs_49_io_reset),
    .io_out(regs_49_io_out),
    .io_enable(regs_49_io_enable)
  );
  FringeFF regs_50 ( // @[RegFile.scala 66:20:@50430.4]
    .clock(regs_50_clock),
    .reset(regs_50_reset),
    .io_in(regs_50_io_in),
    .io_reset(regs_50_io_reset),
    .io_out(regs_50_io_out),
    .io_enable(regs_50_io_enable)
  );
  FringeFF regs_51 ( // @[RegFile.scala 66:20:@50444.4]
    .clock(regs_51_clock),
    .reset(regs_51_reset),
    .io_in(regs_51_io_in),
    .io_reset(regs_51_io_reset),
    .io_out(regs_51_io_out),
    .io_enable(regs_51_io_enable)
  );
  FringeFF regs_52 ( // @[RegFile.scala 66:20:@50458.4]
    .clock(regs_52_clock),
    .reset(regs_52_reset),
    .io_in(regs_52_io_in),
    .io_reset(regs_52_io_reset),
    .io_out(regs_52_io_out),
    .io_enable(regs_52_io_enable)
  );
  FringeFF regs_53 ( // @[RegFile.scala 66:20:@50472.4]
    .clock(regs_53_clock),
    .reset(regs_53_reset),
    .io_in(regs_53_io_in),
    .io_reset(regs_53_io_reset),
    .io_out(regs_53_io_out),
    .io_enable(regs_53_io_enable)
  );
  FringeFF regs_54 ( // @[RegFile.scala 66:20:@50486.4]
    .clock(regs_54_clock),
    .reset(regs_54_reset),
    .io_in(regs_54_io_in),
    .io_reset(regs_54_io_reset),
    .io_out(regs_54_io_out),
    .io_enable(regs_54_io_enable)
  );
  FringeFF regs_55 ( // @[RegFile.scala 66:20:@50500.4]
    .clock(regs_55_clock),
    .reset(regs_55_reset),
    .io_in(regs_55_io_in),
    .io_reset(regs_55_io_reset),
    .io_out(regs_55_io_out),
    .io_enable(regs_55_io_enable)
  );
  FringeFF regs_56 ( // @[RegFile.scala 66:20:@50514.4]
    .clock(regs_56_clock),
    .reset(regs_56_reset),
    .io_in(regs_56_io_in),
    .io_reset(regs_56_io_reset),
    .io_out(regs_56_io_out),
    .io_enable(regs_56_io_enable)
  );
  FringeFF regs_57 ( // @[RegFile.scala 66:20:@50528.4]
    .clock(regs_57_clock),
    .reset(regs_57_reset),
    .io_in(regs_57_io_in),
    .io_reset(regs_57_io_reset),
    .io_out(regs_57_io_out),
    .io_enable(regs_57_io_enable)
  );
  FringeFF regs_58 ( // @[RegFile.scala 66:20:@50542.4]
    .clock(regs_58_clock),
    .reset(regs_58_reset),
    .io_in(regs_58_io_in),
    .io_reset(regs_58_io_reset),
    .io_out(regs_58_io_out),
    .io_enable(regs_58_io_enable)
  );
  FringeFF regs_59 ( // @[RegFile.scala 66:20:@50556.4]
    .clock(regs_59_clock),
    .reset(regs_59_reset),
    .io_in(regs_59_io_in),
    .io_reset(regs_59_io_reset),
    .io_out(regs_59_io_out),
    .io_enable(regs_59_io_enable)
  );
  FringeFF regs_60 ( // @[RegFile.scala 66:20:@50570.4]
    .clock(regs_60_clock),
    .reset(regs_60_reset),
    .io_in(regs_60_io_in),
    .io_reset(regs_60_io_reset),
    .io_out(regs_60_io_out),
    .io_enable(regs_60_io_enable)
  );
  FringeFF regs_61 ( // @[RegFile.scala 66:20:@50584.4]
    .clock(regs_61_clock),
    .reset(regs_61_reset),
    .io_in(regs_61_io_in),
    .io_reset(regs_61_io_reset),
    .io_out(regs_61_io_out),
    .io_enable(regs_61_io_enable)
  );
  FringeFF regs_62 ( // @[RegFile.scala 66:20:@50598.4]
    .clock(regs_62_clock),
    .reset(regs_62_reset),
    .io_in(regs_62_io_in),
    .io_reset(regs_62_io_reset),
    .io_out(regs_62_io_out),
    .io_enable(regs_62_io_enable)
  );
  FringeFF regs_63 ( // @[RegFile.scala 66:20:@50612.4]
    .clock(regs_63_clock),
    .reset(regs_63_reset),
    .io_in(regs_63_io_in),
    .io_reset(regs_63_io_reset),
    .io_out(regs_63_io_out),
    .io_enable(regs_63_io_enable)
  );
  FringeFF regs_64 ( // @[RegFile.scala 66:20:@50626.4]
    .clock(regs_64_clock),
    .reset(regs_64_reset),
    .io_in(regs_64_io_in),
    .io_reset(regs_64_io_reset),
    .io_out(regs_64_io_out),
    .io_enable(regs_64_io_enable)
  );
  FringeFF regs_65 ( // @[RegFile.scala 66:20:@50640.4]
    .clock(regs_65_clock),
    .reset(regs_65_reset),
    .io_in(regs_65_io_in),
    .io_reset(regs_65_io_reset),
    .io_out(regs_65_io_out),
    .io_enable(regs_65_io_enable)
  );
  FringeFF regs_66 ( // @[RegFile.scala 66:20:@50654.4]
    .clock(regs_66_clock),
    .reset(regs_66_reset),
    .io_in(regs_66_io_in),
    .io_reset(regs_66_io_reset),
    .io_out(regs_66_io_out),
    .io_enable(regs_66_io_enable)
  );
  FringeFF regs_67 ( // @[RegFile.scala 66:20:@50668.4]
    .clock(regs_67_clock),
    .reset(regs_67_reset),
    .io_in(regs_67_io_in),
    .io_reset(regs_67_io_reset),
    .io_out(regs_67_io_out),
    .io_enable(regs_67_io_enable)
  );
  FringeFF regs_68 ( // @[RegFile.scala 66:20:@50682.4]
    .clock(regs_68_clock),
    .reset(regs_68_reset),
    .io_in(regs_68_io_in),
    .io_reset(regs_68_io_reset),
    .io_out(regs_68_io_out),
    .io_enable(regs_68_io_enable)
  );
  FringeFF regs_69 ( // @[RegFile.scala 66:20:@50696.4]
    .clock(regs_69_clock),
    .reset(regs_69_reset),
    .io_in(regs_69_io_in),
    .io_reset(regs_69_io_reset),
    .io_out(regs_69_io_out),
    .io_enable(regs_69_io_enable)
  );
  FringeFF regs_70 ( // @[RegFile.scala 66:20:@50710.4]
    .clock(regs_70_clock),
    .reset(regs_70_reset),
    .io_in(regs_70_io_in),
    .io_reset(regs_70_io_reset),
    .io_out(regs_70_io_out),
    .io_enable(regs_70_io_enable)
  );
  FringeFF regs_71 ( // @[RegFile.scala 66:20:@50724.4]
    .clock(regs_71_clock),
    .reset(regs_71_reset),
    .io_in(regs_71_io_in),
    .io_reset(regs_71_io_reset),
    .io_out(regs_71_io_out),
    .io_enable(regs_71_io_enable)
  );
  FringeFF regs_72 ( // @[RegFile.scala 66:20:@50738.4]
    .clock(regs_72_clock),
    .reset(regs_72_reset),
    .io_in(regs_72_io_in),
    .io_reset(regs_72_io_reset),
    .io_out(regs_72_io_out),
    .io_enable(regs_72_io_enable)
  );
  FringeFF regs_73 ( // @[RegFile.scala 66:20:@50752.4]
    .clock(regs_73_clock),
    .reset(regs_73_reset),
    .io_in(regs_73_io_in),
    .io_reset(regs_73_io_reset),
    .io_out(regs_73_io_out),
    .io_enable(regs_73_io_enable)
  );
  FringeFF regs_74 ( // @[RegFile.scala 66:20:@50766.4]
    .clock(regs_74_clock),
    .reset(regs_74_reset),
    .io_in(regs_74_io_in),
    .io_reset(regs_74_io_reset),
    .io_out(regs_74_io_out),
    .io_enable(regs_74_io_enable)
  );
  FringeFF regs_75 ( // @[RegFile.scala 66:20:@50780.4]
    .clock(regs_75_clock),
    .reset(regs_75_reset),
    .io_in(regs_75_io_in),
    .io_reset(regs_75_io_reset),
    .io_out(regs_75_io_out),
    .io_enable(regs_75_io_enable)
  );
  FringeFF regs_76 ( // @[RegFile.scala 66:20:@50794.4]
    .clock(regs_76_clock),
    .reset(regs_76_reset),
    .io_in(regs_76_io_in),
    .io_reset(regs_76_io_reset),
    .io_out(regs_76_io_out),
    .io_enable(regs_76_io_enable)
  );
  FringeFF regs_77 ( // @[RegFile.scala 66:20:@50808.4]
    .clock(regs_77_clock),
    .reset(regs_77_reset),
    .io_in(regs_77_io_in),
    .io_reset(regs_77_io_reset),
    .io_out(regs_77_io_out),
    .io_enable(regs_77_io_enable)
  );
  FringeFF regs_78 ( // @[RegFile.scala 66:20:@50822.4]
    .clock(regs_78_clock),
    .reset(regs_78_reset),
    .io_in(regs_78_io_in),
    .io_reset(regs_78_io_reset),
    .io_out(regs_78_io_out),
    .io_enable(regs_78_io_enable)
  );
  FringeFF regs_79 ( // @[RegFile.scala 66:20:@50836.4]
    .clock(regs_79_clock),
    .reset(regs_79_reset),
    .io_in(regs_79_io_in),
    .io_reset(regs_79_io_reset),
    .io_out(regs_79_io_out),
    .io_enable(regs_79_io_enable)
  );
  FringeFF regs_80 ( // @[RegFile.scala 66:20:@50850.4]
    .clock(regs_80_clock),
    .reset(regs_80_reset),
    .io_in(regs_80_io_in),
    .io_reset(regs_80_io_reset),
    .io_out(regs_80_io_out),
    .io_enable(regs_80_io_enable)
  );
  FringeFF regs_81 ( // @[RegFile.scala 66:20:@50864.4]
    .clock(regs_81_clock),
    .reset(regs_81_reset),
    .io_in(regs_81_io_in),
    .io_reset(regs_81_io_reset),
    .io_out(regs_81_io_out),
    .io_enable(regs_81_io_enable)
  );
  FringeFF regs_82 ( // @[RegFile.scala 66:20:@50878.4]
    .clock(regs_82_clock),
    .reset(regs_82_reset),
    .io_in(regs_82_io_in),
    .io_reset(regs_82_io_reset),
    .io_out(regs_82_io_out),
    .io_enable(regs_82_io_enable)
  );
  FringeFF regs_83 ( // @[RegFile.scala 66:20:@50892.4]
    .clock(regs_83_clock),
    .reset(regs_83_reset),
    .io_in(regs_83_io_in),
    .io_reset(regs_83_io_reset),
    .io_out(regs_83_io_out),
    .io_enable(regs_83_io_enable)
  );
  FringeFF regs_84 ( // @[RegFile.scala 66:20:@50906.4]
    .clock(regs_84_clock),
    .reset(regs_84_reset),
    .io_in(regs_84_io_in),
    .io_reset(regs_84_io_reset),
    .io_out(regs_84_io_out),
    .io_enable(regs_84_io_enable)
  );
  FringeFF regs_85 ( // @[RegFile.scala 66:20:@50920.4]
    .clock(regs_85_clock),
    .reset(regs_85_reset),
    .io_in(regs_85_io_in),
    .io_reset(regs_85_io_reset),
    .io_out(regs_85_io_out),
    .io_enable(regs_85_io_enable)
  );
  FringeFF regs_86 ( // @[RegFile.scala 66:20:@50934.4]
    .clock(regs_86_clock),
    .reset(regs_86_reset),
    .io_in(regs_86_io_in),
    .io_reset(regs_86_io_reset),
    .io_out(regs_86_io_out),
    .io_enable(regs_86_io_enable)
  );
  FringeFF regs_87 ( // @[RegFile.scala 66:20:@50948.4]
    .clock(regs_87_clock),
    .reset(regs_87_reset),
    .io_in(regs_87_io_in),
    .io_reset(regs_87_io_reset),
    .io_out(regs_87_io_out),
    .io_enable(regs_87_io_enable)
  );
  FringeFF regs_88 ( // @[RegFile.scala 66:20:@50962.4]
    .clock(regs_88_clock),
    .reset(regs_88_reset),
    .io_in(regs_88_io_in),
    .io_reset(regs_88_io_reset),
    .io_out(regs_88_io_out),
    .io_enable(regs_88_io_enable)
  );
  FringeFF regs_89 ( // @[RegFile.scala 66:20:@50976.4]
    .clock(regs_89_clock),
    .reset(regs_89_reset),
    .io_in(regs_89_io_in),
    .io_reset(regs_89_io_reset),
    .io_out(regs_89_io_out),
    .io_enable(regs_89_io_enable)
  );
  FringeFF regs_90 ( // @[RegFile.scala 66:20:@50990.4]
    .clock(regs_90_clock),
    .reset(regs_90_reset),
    .io_in(regs_90_io_in),
    .io_reset(regs_90_io_reset),
    .io_out(regs_90_io_out),
    .io_enable(regs_90_io_enable)
  );
  FringeFF regs_91 ( // @[RegFile.scala 66:20:@51004.4]
    .clock(regs_91_clock),
    .reset(regs_91_reset),
    .io_in(regs_91_io_in),
    .io_reset(regs_91_io_reset),
    .io_out(regs_91_io_out),
    .io_enable(regs_91_io_enable)
  );
  FringeFF regs_92 ( // @[RegFile.scala 66:20:@51018.4]
    .clock(regs_92_clock),
    .reset(regs_92_reset),
    .io_in(regs_92_io_in),
    .io_reset(regs_92_io_reset),
    .io_out(regs_92_io_out),
    .io_enable(regs_92_io_enable)
  );
  FringeFF regs_93 ( // @[RegFile.scala 66:20:@51032.4]
    .clock(regs_93_clock),
    .reset(regs_93_reset),
    .io_in(regs_93_io_in),
    .io_reset(regs_93_io_reset),
    .io_out(regs_93_io_out),
    .io_enable(regs_93_io_enable)
  );
  FringeFF regs_94 ( // @[RegFile.scala 66:20:@51046.4]
    .clock(regs_94_clock),
    .reset(regs_94_reset),
    .io_in(regs_94_io_in),
    .io_reset(regs_94_io_reset),
    .io_out(regs_94_io_out),
    .io_enable(regs_94_io_enable)
  );
  FringeFF regs_95 ( // @[RegFile.scala 66:20:@51060.4]
    .clock(regs_95_clock),
    .reset(regs_95_reset),
    .io_in(regs_95_io_in),
    .io_reset(regs_95_io_reset),
    .io_out(regs_95_io_out),
    .io_enable(regs_95_io_enable)
  );
  FringeFF regs_96 ( // @[RegFile.scala 66:20:@51074.4]
    .clock(regs_96_clock),
    .reset(regs_96_reset),
    .io_in(regs_96_io_in),
    .io_reset(regs_96_io_reset),
    .io_out(regs_96_io_out),
    .io_enable(regs_96_io_enable)
  );
  FringeFF regs_97 ( // @[RegFile.scala 66:20:@51088.4]
    .clock(regs_97_clock),
    .reset(regs_97_reset),
    .io_in(regs_97_io_in),
    .io_reset(regs_97_io_reset),
    .io_out(regs_97_io_out),
    .io_enable(regs_97_io_enable)
  );
  FringeFF regs_98 ( // @[RegFile.scala 66:20:@51102.4]
    .clock(regs_98_clock),
    .reset(regs_98_reset),
    .io_in(regs_98_io_in),
    .io_reset(regs_98_io_reset),
    .io_out(regs_98_io_out),
    .io_enable(regs_98_io_enable)
  );
  FringeFF regs_99 ( // @[RegFile.scala 66:20:@51116.4]
    .clock(regs_99_clock),
    .reset(regs_99_reset),
    .io_in(regs_99_io_in),
    .io_reset(regs_99_io_reset),
    .io_out(regs_99_io_out),
    .io_enable(regs_99_io_enable)
  );
  FringeFF regs_100 ( // @[RegFile.scala 66:20:@51130.4]
    .clock(regs_100_clock),
    .reset(regs_100_reset),
    .io_in(regs_100_io_in),
    .io_reset(regs_100_io_reset),
    .io_out(regs_100_io_out),
    .io_enable(regs_100_io_enable)
  );
  FringeFF regs_101 ( // @[RegFile.scala 66:20:@51144.4]
    .clock(regs_101_clock),
    .reset(regs_101_reset),
    .io_in(regs_101_io_in),
    .io_reset(regs_101_io_reset),
    .io_out(regs_101_io_out),
    .io_enable(regs_101_io_enable)
  );
  FringeFF regs_102 ( // @[RegFile.scala 66:20:@51158.4]
    .clock(regs_102_clock),
    .reset(regs_102_reset),
    .io_in(regs_102_io_in),
    .io_reset(regs_102_io_reset),
    .io_out(regs_102_io_out),
    .io_enable(regs_102_io_enable)
  );
  FringeFF regs_103 ( // @[RegFile.scala 66:20:@51172.4]
    .clock(regs_103_clock),
    .reset(regs_103_reset),
    .io_in(regs_103_io_in),
    .io_reset(regs_103_io_reset),
    .io_out(regs_103_io_out),
    .io_enable(regs_103_io_enable)
  );
  FringeFF regs_104 ( // @[RegFile.scala 66:20:@51186.4]
    .clock(regs_104_clock),
    .reset(regs_104_reset),
    .io_in(regs_104_io_in),
    .io_reset(regs_104_io_reset),
    .io_out(regs_104_io_out),
    .io_enable(regs_104_io_enable)
  );
  FringeFF regs_105 ( // @[RegFile.scala 66:20:@51200.4]
    .clock(regs_105_clock),
    .reset(regs_105_reset),
    .io_in(regs_105_io_in),
    .io_reset(regs_105_io_reset),
    .io_out(regs_105_io_out),
    .io_enable(regs_105_io_enable)
  );
  FringeFF regs_106 ( // @[RegFile.scala 66:20:@51214.4]
    .clock(regs_106_clock),
    .reset(regs_106_reset),
    .io_in(regs_106_io_in),
    .io_reset(regs_106_io_reset),
    .io_out(regs_106_io_out),
    .io_enable(regs_106_io_enable)
  );
  FringeFF regs_107 ( // @[RegFile.scala 66:20:@51228.4]
    .clock(regs_107_clock),
    .reset(regs_107_reset),
    .io_in(regs_107_io_in),
    .io_reset(regs_107_io_reset),
    .io_out(regs_107_io_out),
    .io_enable(regs_107_io_enable)
  );
  FringeFF regs_108 ( // @[RegFile.scala 66:20:@51242.4]
    .clock(regs_108_clock),
    .reset(regs_108_reset),
    .io_in(regs_108_io_in),
    .io_reset(regs_108_io_reset),
    .io_out(regs_108_io_out),
    .io_enable(regs_108_io_enable)
  );
  FringeFF regs_109 ( // @[RegFile.scala 66:20:@51256.4]
    .clock(regs_109_clock),
    .reset(regs_109_reset),
    .io_in(regs_109_io_in),
    .io_reset(regs_109_io_reset),
    .io_out(regs_109_io_out),
    .io_enable(regs_109_io_enable)
  );
  FringeFF regs_110 ( // @[RegFile.scala 66:20:@51270.4]
    .clock(regs_110_clock),
    .reset(regs_110_reset),
    .io_in(regs_110_io_in),
    .io_reset(regs_110_io_reset),
    .io_out(regs_110_io_out),
    .io_enable(regs_110_io_enable)
  );
  FringeFF regs_111 ( // @[RegFile.scala 66:20:@51284.4]
    .clock(regs_111_clock),
    .reset(regs_111_reset),
    .io_in(regs_111_io_in),
    .io_reset(regs_111_io_reset),
    .io_out(regs_111_io_out),
    .io_enable(regs_111_io_enable)
  );
  FringeFF regs_112 ( // @[RegFile.scala 66:20:@51298.4]
    .clock(regs_112_clock),
    .reset(regs_112_reset),
    .io_in(regs_112_io_in),
    .io_reset(regs_112_io_reset),
    .io_out(regs_112_io_out),
    .io_enable(regs_112_io_enable)
  );
  FringeFF regs_113 ( // @[RegFile.scala 66:20:@51312.4]
    .clock(regs_113_clock),
    .reset(regs_113_reset),
    .io_in(regs_113_io_in),
    .io_reset(regs_113_io_reset),
    .io_out(regs_113_io_out),
    .io_enable(regs_113_io_enable)
  );
  FringeFF regs_114 ( // @[RegFile.scala 66:20:@51326.4]
    .clock(regs_114_clock),
    .reset(regs_114_reset),
    .io_in(regs_114_io_in),
    .io_reset(regs_114_io_reset),
    .io_out(regs_114_io_out),
    .io_enable(regs_114_io_enable)
  );
  FringeFF regs_115 ( // @[RegFile.scala 66:20:@51340.4]
    .clock(regs_115_clock),
    .reset(regs_115_reset),
    .io_in(regs_115_io_in),
    .io_reset(regs_115_io_reset),
    .io_out(regs_115_io_out),
    .io_enable(regs_115_io_enable)
  );
  FringeFF regs_116 ( // @[RegFile.scala 66:20:@51354.4]
    .clock(regs_116_clock),
    .reset(regs_116_reset),
    .io_in(regs_116_io_in),
    .io_reset(regs_116_io_reset),
    .io_out(regs_116_io_out),
    .io_enable(regs_116_io_enable)
  );
  FringeFF regs_117 ( // @[RegFile.scala 66:20:@51368.4]
    .clock(regs_117_clock),
    .reset(regs_117_reset),
    .io_in(regs_117_io_in),
    .io_reset(regs_117_io_reset),
    .io_out(regs_117_io_out),
    .io_enable(regs_117_io_enable)
  );
  FringeFF regs_118 ( // @[RegFile.scala 66:20:@51382.4]
    .clock(regs_118_clock),
    .reset(regs_118_reset),
    .io_in(regs_118_io_in),
    .io_reset(regs_118_io_reset),
    .io_out(regs_118_io_out),
    .io_enable(regs_118_io_enable)
  );
  FringeFF regs_119 ( // @[RegFile.scala 66:20:@51396.4]
    .clock(regs_119_clock),
    .reset(regs_119_reset),
    .io_in(regs_119_io_in),
    .io_reset(regs_119_io_reset),
    .io_out(regs_119_io_out),
    .io_enable(regs_119_io_enable)
  );
  FringeFF regs_120 ( // @[RegFile.scala 66:20:@51410.4]
    .clock(regs_120_clock),
    .reset(regs_120_reset),
    .io_in(regs_120_io_in),
    .io_reset(regs_120_io_reset),
    .io_out(regs_120_io_out),
    .io_enable(regs_120_io_enable)
  );
  FringeFF regs_121 ( // @[RegFile.scala 66:20:@51424.4]
    .clock(regs_121_clock),
    .reset(regs_121_reset),
    .io_in(regs_121_io_in),
    .io_reset(regs_121_io_reset),
    .io_out(regs_121_io_out),
    .io_enable(regs_121_io_enable)
  );
  FringeFF regs_122 ( // @[RegFile.scala 66:20:@51438.4]
    .clock(regs_122_clock),
    .reset(regs_122_reset),
    .io_in(regs_122_io_in),
    .io_reset(regs_122_io_reset),
    .io_out(regs_122_io_out),
    .io_enable(regs_122_io_enable)
  );
  FringeFF regs_123 ( // @[RegFile.scala 66:20:@51452.4]
    .clock(regs_123_clock),
    .reset(regs_123_reset),
    .io_in(regs_123_io_in),
    .io_reset(regs_123_io_reset),
    .io_out(regs_123_io_out),
    .io_enable(regs_123_io_enable)
  );
  FringeFF regs_124 ( // @[RegFile.scala 66:20:@51466.4]
    .clock(regs_124_clock),
    .reset(regs_124_reset),
    .io_in(regs_124_io_in),
    .io_reset(regs_124_io_reset),
    .io_out(regs_124_io_out),
    .io_enable(regs_124_io_enable)
  );
  FringeFF regs_125 ( // @[RegFile.scala 66:20:@51480.4]
    .clock(regs_125_clock),
    .reset(regs_125_reset),
    .io_in(regs_125_io_in),
    .io_reset(regs_125_io_reset),
    .io_out(regs_125_io_out),
    .io_enable(regs_125_io_enable)
  );
  FringeFF regs_126 ( // @[RegFile.scala 66:20:@51494.4]
    .clock(regs_126_clock),
    .reset(regs_126_reset),
    .io_in(regs_126_io_in),
    .io_reset(regs_126_io_reset),
    .io_out(regs_126_io_out),
    .io_enable(regs_126_io_enable)
  );
  FringeFF regs_127 ( // @[RegFile.scala 66:20:@51508.4]
    .clock(regs_127_clock),
    .reset(regs_127_reset),
    .io_in(regs_127_io_in),
    .io_reset(regs_127_io_reset),
    .io_out(regs_127_io_out),
    .io_enable(regs_127_io_enable)
  );
  FringeFF regs_128 ( // @[RegFile.scala 66:20:@51522.4]
    .clock(regs_128_clock),
    .reset(regs_128_reset),
    .io_in(regs_128_io_in),
    .io_reset(regs_128_io_reset),
    .io_out(regs_128_io_out),
    .io_enable(regs_128_io_enable)
  );
  FringeFF regs_129 ( // @[RegFile.scala 66:20:@51536.4]
    .clock(regs_129_clock),
    .reset(regs_129_reset),
    .io_in(regs_129_io_in),
    .io_reset(regs_129_io_reset),
    .io_out(regs_129_io_out),
    .io_enable(regs_129_io_enable)
  );
  FringeFF regs_130 ( // @[RegFile.scala 66:20:@51550.4]
    .clock(regs_130_clock),
    .reset(regs_130_reset),
    .io_in(regs_130_io_in),
    .io_reset(regs_130_io_reset),
    .io_out(regs_130_io_out),
    .io_enable(regs_130_io_enable)
  );
  FringeFF regs_131 ( // @[RegFile.scala 66:20:@51564.4]
    .clock(regs_131_clock),
    .reset(regs_131_reset),
    .io_in(regs_131_io_in),
    .io_reset(regs_131_io_reset),
    .io_out(regs_131_io_out),
    .io_enable(regs_131_io_enable)
  );
  FringeFF regs_132 ( // @[RegFile.scala 66:20:@51578.4]
    .clock(regs_132_clock),
    .reset(regs_132_reset),
    .io_in(regs_132_io_in),
    .io_reset(regs_132_io_reset),
    .io_out(regs_132_io_out),
    .io_enable(regs_132_io_enable)
  );
  FringeFF regs_133 ( // @[RegFile.scala 66:20:@51592.4]
    .clock(regs_133_clock),
    .reset(regs_133_reset),
    .io_in(regs_133_io_in),
    .io_reset(regs_133_io_reset),
    .io_out(regs_133_io_out),
    .io_enable(regs_133_io_enable)
  );
  FringeFF regs_134 ( // @[RegFile.scala 66:20:@51606.4]
    .clock(regs_134_clock),
    .reset(regs_134_reset),
    .io_in(regs_134_io_in),
    .io_reset(regs_134_io_reset),
    .io_out(regs_134_io_out),
    .io_enable(regs_134_io_enable)
  );
  FringeFF regs_135 ( // @[RegFile.scala 66:20:@51620.4]
    .clock(regs_135_clock),
    .reset(regs_135_reset),
    .io_in(regs_135_io_in),
    .io_reset(regs_135_io_reset),
    .io_out(regs_135_io_out),
    .io_enable(regs_135_io_enable)
  );
  FringeFF regs_136 ( // @[RegFile.scala 66:20:@51634.4]
    .clock(regs_136_clock),
    .reset(regs_136_reset),
    .io_in(regs_136_io_in),
    .io_reset(regs_136_io_reset),
    .io_out(regs_136_io_out),
    .io_enable(regs_136_io_enable)
  );
  FringeFF regs_137 ( // @[RegFile.scala 66:20:@51648.4]
    .clock(regs_137_clock),
    .reset(regs_137_reset),
    .io_in(regs_137_io_in),
    .io_reset(regs_137_io_reset),
    .io_out(regs_137_io_out),
    .io_enable(regs_137_io_enable)
  );
  FringeFF regs_138 ( // @[RegFile.scala 66:20:@51662.4]
    .clock(regs_138_clock),
    .reset(regs_138_reset),
    .io_in(regs_138_io_in),
    .io_reset(regs_138_io_reset),
    .io_out(regs_138_io_out),
    .io_enable(regs_138_io_enable)
  );
  FringeFF regs_139 ( // @[RegFile.scala 66:20:@51676.4]
    .clock(regs_139_clock),
    .reset(regs_139_reset),
    .io_in(regs_139_io_in),
    .io_reset(regs_139_io_reset),
    .io_out(regs_139_io_out),
    .io_enable(regs_139_io_enable)
  );
  FringeFF regs_140 ( // @[RegFile.scala 66:20:@51690.4]
    .clock(regs_140_clock),
    .reset(regs_140_reset),
    .io_in(regs_140_io_in),
    .io_reset(regs_140_io_reset),
    .io_out(regs_140_io_out),
    .io_enable(regs_140_io_enable)
  );
  FringeFF regs_141 ( // @[RegFile.scala 66:20:@51704.4]
    .clock(regs_141_clock),
    .reset(regs_141_reset),
    .io_in(regs_141_io_in),
    .io_reset(regs_141_io_reset),
    .io_out(regs_141_io_out),
    .io_enable(regs_141_io_enable)
  );
  FringeFF regs_142 ( // @[RegFile.scala 66:20:@51718.4]
    .clock(regs_142_clock),
    .reset(regs_142_reset),
    .io_in(regs_142_io_in),
    .io_reset(regs_142_io_reset),
    .io_out(regs_142_io_out),
    .io_enable(regs_142_io_enable)
  );
  FringeFF regs_143 ( // @[RegFile.scala 66:20:@51732.4]
    .clock(regs_143_clock),
    .reset(regs_143_reset),
    .io_in(regs_143_io_in),
    .io_reset(regs_143_io_reset),
    .io_out(regs_143_io_out),
    .io_enable(regs_143_io_enable)
  );
  FringeFF regs_144 ( // @[RegFile.scala 66:20:@51746.4]
    .clock(regs_144_clock),
    .reset(regs_144_reset),
    .io_in(regs_144_io_in),
    .io_reset(regs_144_io_reset),
    .io_out(regs_144_io_out),
    .io_enable(regs_144_io_enable)
  );
  FringeFF regs_145 ( // @[RegFile.scala 66:20:@51760.4]
    .clock(regs_145_clock),
    .reset(regs_145_reset),
    .io_in(regs_145_io_in),
    .io_reset(regs_145_io_reset),
    .io_out(regs_145_io_out),
    .io_enable(regs_145_io_enable)
  );
  FringeFF regs_146 ( // @[RegFile.scala 66:20:@51774.4]
    .clock(regs_146_clock),
    .reset(regs_146_reset),
    .io_in(regs_146_io_in),
    .io_reset(regs_146_io_reset),
    .io_out(regs_146_io_out),
    .io_enable(regs_146_io_enable)
  );
  FringeFF regs_147 ( // @[RegFile.scala 66:20:@51788.4]
    .clock(regs_147_clock),
    .reset(regs_147_reset),
    .io_in(regs_147_io_in),
    .io_reset(regs_147_io_reset),
    .io_out(regs_147_io_out),
    .io_enable(regs_147_io_enable)
  );
  FringeFF regs_148 ( // @[RegFile.scala 66:20:@51802.4]
    .clock(regs_148_clock),
    .reset(regs_148_reset),
    .io_in(regs_148_io_in),
    .io_reset(regs_148_io_reset),
    .io_out(regs_148_io_out),
    .io_enable(regs_148_io_enable)
  );
  FringeFF regs_149 ( // @[RegFile.scala 66:20:@51816.4]
    .clock(regs_149_clock),
    .reset(regs_149_reset),
    .io_in(regs_149_io_in),
    .io_reset(regs_149_io_reset),
    .io_out(regs_149_io_out),
    .io_enable(regs_149_io_enable)
  );
  FringeFF regs_150 ( // @[RegFile.scala 66:20:@51830.4]
    .clock(regs_150_clock),
    .reset(regs_150_reset),
    .io_in(regs_150_io_in),
    .io_reset(regs_150_io_reset),
    .io_out(regs_150_io_out),
    .io_enable(regs_150_io_enable)
  );
  FringeFF regs_151 ( // @[RegFile.scala 66:20:@51844.4]
    .clock(regs_151_clock),
    .reset(regs_151_reset),
    .io_in(regs_151_io_in),
    .io_reset(regs_151_io_reset),
    .io_out(regs_151_io_out),
    .io_enable(regs_151_io_enable)
  );
  FringeFF regs_152 ( // @[RegFile.scala 66:20:@51858.4]
    .clock(regs_152_clock),
    .reset(regs_152_reset),
    .io_in(regs_152_io_in),
    .io_reset(regs_152_io_reset),
    .io_out(regs_152_io_out),
    .io_enable(regs_152_io_enable)
  );
  FringeFF regs_153 ( // @[RegFile.scala 66:20:@51872.4]
    .clock(regs_153_clock),
    .reset(regs_153_reset),
    .io_in(regs_153_io_in),
    .io_reset(regs_153_io_reset),
    .io_out(regs_153_io_out),
    .io_enable(regs_153_io_enable)
  );
  FringeFF regs_154 ( // @[RegFile.scala 66:20:@51886.4]
    .clock(regs_154_clock),
    .reset(regs_154_reset),
    .io_in(regs_154_io_in),
    .io_reset(regs_154_io_reset),
    .io_out(regs_154_io_out),
    .io_enable(regs_154_io_enable)
  );
  FringeFF regs_155 ( // @[RegFile.scala 66:20:@51900.4]
    .clock(regs_155_clock),
    .reset(regs_155_reset),
    .io_in(regs_155_io_in),
    .io_reset(regs_155_io_reset),
    .io_out(regs_155_io_out),
    .io_enable(regs_155_io_enable)
  );
  FringeFF regs_156 ( // @[RegFile.scala 66:20:@51914.4]
    .clock(regs_156_clock),
    .reset(regs_156_reset),
    .io_in(regs_156_io_in),
    .io_reset(regs_156_io_reset),
    .io_out(regs_156_io_out),
    .io_enable(regs_156_io_enable)
  );
  FringeFF regs_157 ( // @[RegFile.scala 66:20:@51928.4]
    .clock(regs_157_clock),
    .reset(regs_157_reset),
    .io_in(regs_157_io_in),
    .io_reset(regs_157_io_reset),
    .io_out(regs_157_io_out),
    .io_enable(regs_157_io_enable)
  );
  FringeFF regs_158 ( // @[RegFile.scala 66:20:@51942.4]
    .clock(regs_158_clock),
    .reset(regs_158_reset),
    .io_in(regs_158_io_in),
    .io_reset(regs_158_io_reset),
    .io_out(regs_158_io_out),
    .io_enable(regs_158_io_enable)
  );
  FringeFF regs_159 ( // @[RegFile.scala 66:20:@51956.4]
    .clock(regs_159_clock),
    .reset(regs_159_reset),
    .io_in(regs_159_io_in),
    .io_reset(regs_159_io_reset),
    .io_out(regs_159_io_out),
    .io_enable(regs_159_io_enable)
  );
  FringeFF regs_160 ( // @[RegFile.scala 66:20:@51970.4]
    .clock(regs_160_clock),
    .reset(regs_160_reset),
    .io_in(regs_160_io_in),
    .io_reset(regs_160_io_reset),
    .io_out(regs_160_io_out),
    .io_enable(regs_160_io_enable)
  );
  FringeFF regs_161 ( // @[RegFile.scala 66:20:@51984.4]
    .clock(regs_161_clock),
    .reset(regs_161_reset),
    .io_in(regs_161_io_in),
    .io_reset(regs_161_io_reset),
    .io_out(regs_161_io_out),
    .io_enable(regs_161_io_enable)
  );
  FringeFF regs_162 ( // @[RegFile.scala 66:20:@51998.4]
    .clock(regs_162_clock),
    .reset(regs_162_reset),
    .io_in(regs_162_io_in),
    .io_reset(regs_162_io_reset),
    .io_out(regs_162_io_out),
    .io_enable(regs_162_io_enable)
  );
  FringeFF regs_163 ( // @[RegFile.scala 66:20:@52012.4]
    .clock(regs_163_clock),
    .reset(regs_163_reset),
    .io_in(regs_163_io_in),
    .io_reset(regs_163_io_reset),
    .io_out(regs_163_io_out),
    .io_enable(regs_163_io_enable)
  );
  FringeFF regs_164 ( // @[RegFile.scala 66:20:@52026.4]
    .clock(regs_164_clock),
    .reset(regs_164_reset),
    .io_in(regs_164_io_in),
    .io_reset(regs_164_io_reset),
    .io_out(regs_164_io_out),
    .io_enable(regs_164_io_enable)
  );
  FringeFF regs_165 ( // @[RegFile.scala 66:20:@52040.4]
    .clock(regs_165_clock),
    .reset(regs_165_reset),
    .io_in(regs_165_io_in),
    .io_reset(regs_165_io_reset),
    .io_out(regs_165_io_out),
    .io_enable(regs_165_io_enable)
  );
  FringeFF regs_166 ( // @[RegFile.scala 66:20:@52054.4]
    .clock(regs_166_clock),
    .reset(regs_166_reset),
    .io_in(regs_166_io_in),
    .io_reset(regs_166_io_reset),
    .io_out(regs_166_io_out),
    .io_enable(regs_166_io_enable)
  );
  FringeFF regs_167 ( // @[RegFile.scala 66:20:@52068.4]
    .clock(regs_167_clock),
    .reset(regs_167_reset),
    .io_in(regs_167_io_in),
    .io_reset(regs_167_io_reset),
    .io_out(regs_167_io_out),
    .io_enable(regs_167_io_enable)
  );
  FringeFF regs_168 ( // @[RegFile.scala 66:20:@52082.4]
    .clock(regs_168_clock),
    .reset(regs_168_reset),
    .io_in(regs_168_io_in),
    .io_reset(regs_168_io_reset),
    .io_out(regs_168_io_out),
    .io_enable(regs_168_io_enable)
  );
  FringeFF regs_169 ( // @[RegFile.scala 66:20:@52096.4]
    .clock(regs_169_clock),
    .reset(regs_169_reset),
    .io_in(regs_169_io_in),
    .io_reset(regs_169_io_reset),
    .io_out(regs_169_io_out),
    .io_enable(regs_169_io_enable)
  );
  FringeFF regs_170 ( // @[RegFile.scala 66:20:@52110.4]
    .clock(regs_170_clock),
    .reset(regs_170_reset),
    .io_in(regs_170_io_in),
    .io_reset(regs_170_io_reset),
    .io_out(regs_170_io_out),
    .io_enable(regs_170_io_enable)
  );
  FringeFF regs_171 ( // @[RegFile.scala 66:20:@52124.4]
    .clock(regs_171_clock),
    .reset(regs_171_reset),
    .io_in(regs_171_io_in),
    .io_reset(regs_171_io_reset),
    .io_out(regs_171_io_out),
    .io_enable(regs_171_io_enable)
  );
  FringeFF regs_172 ( // @[RegFile.scala 66:20:@52138.4]
    .clock(regs_172_clock),
    .reset(regs_172_reset),
    .io_in(regs_172_io_in),
    .io_reset(regs_172_io_reset),
    .io_out(regs_172_io_out),
    .io_enable(regs_172_io_enable)
  );
  FringeFF regs_173 ( // @[RegFile.scala 66:20:@52152.4]
    .clock(regs_173_clock),
    .reset(regs_173_reset),
    .io_in(regs_173_io_in),
    .io_reset(regs_173_io_reset),
    .io_out(regs_173_io_out),
    .io_enable(regs_173_io_enable)
  );
  FringeFF regs_174 ( // @[RegFile.scala 66:20:@52166.4]
    .clock(regs_174_clock),
    .reset(regs_174_reset),
    .io_in(regs_174_io_in),
    .io_reset(regs_174_io_reset),
    .io_out(regs_174_io_out),
    .io_enable(regs_174_io_enable)
  );
  FringeFF regs_175 ( // @[RegFile.scala 66:20:@52180.4]
    .clock(regs_175_clock),
    .reset(regs_175_reset),
    .io_in(regs_175_io_in),
    .io_reset(regs_175_io_reset),
    .io_out(regs_175_io_out),
    .io_enable(regs_175_io_enable)
  );
  FringeFF regs_176 ( // @[RegFile.scala 66:20:@52194.4]
    .clock(regs_176_clock),
    .reset(regs_176_reset),
    .io_in(regs_176_io_in),
    .io_reset(regs_176_io_reset),
    .io_out(regs_176_io_out),
    .io_enable(regs_176_io_enable)
  );
  FringeFF regs_177 ( // @[RegFile.scala 66:20:@52208.4]
    .clock(regs_177_clock),
    .reset(regs_177_reset),
    .io_in(regs_177_io_in),
    .io_reset(regs_177_io_reset),
    .io_out(regs_177_io_out),
    .io_enable(regs_177_io_enable)
  );
  FringeFF regs_178 ( // @[RegFile.scala 66:20:@52222.4]
    .clock(regs_178_clock),
    .reset(regs_178_reset),
    .io_in(regs_178_io_in),
    .io_reset(regs_178_io_reset),
    .io_out(regs_178_io_out),
    .io_enable(regs_178_io_enable)
  );
  FringeFF regs_179 ( // @[RegFile.scala 66:20:@52236.4]
    .clock(regs_179_clock),
    .reset(regs_179_reset),
    .io_in(regs_179_io_in),
    .io_reset(regs_179_io_reset),
    .io_out(regs_179_io_out),
    .io_enable(regs_179_io_enable)
  );
  FringeFF regs_180 ( // @[RegFile.scala 66:20:@52250.4]
    .clock(regs_180_clock),
    .reset(regs_180_reset),
    .io_in(regs_180_io_in),
    .io_reset(regs_180_io_reset),
    .io_out(regs_180_io_out),
    .io_enable(regs_180_io_enable)
  );
  FringeFF regs_181 ( // @[RegFile.scala 66:20:@52264.4]
    .clock(regs_181_clock),
    .reset(regs_181_reset),
    .io_in(regs_181_io_in),
    .io_reset(regs_181_io_reset),
    .io_out(regs_181_io_out),
    .io_enable(regs_181_io_enable)
  );
  FringeFF regs_182 ( // @[RegFile.scala 66:20:@52278.4]
    .clock(regs_182_clock),
    .reset(regs_182_reset),
    .io_in(regs_182_io_in),
    .io_reset(regs_182_io_reset),
    .io_out(regs_182_io_out),
    .io_enable(regs_182_io_enable)
  );
  FringeFF regs_183 ( // @[RegFile.scala 66:20:@52292.4]
    .clock(regs_183_clock),
    .reset(regs_183_reset),
    .io_in(regs_183_io_in),
    .io_reset(regs_183_io_reset),
    .io_out(regs_183_io_out),
    .io_enable(regs_183_io_enable)
  );
  FringeFF regs_184 ( // @[RegFile.scala 66:20:@52306.4]
    .clock(regs_184_clock),
    .reset(regs_184_reset),
    .io_in(regs_184_io_in),
    .io_reset(regs_184_io_reset),
    .io_out(regs_184_io_out),
    .io_enable(regs_184_io_enable)
  );
  FringeFF regs_185 ( // @[RegFile.scala 66:20:@52320.4]
    .clock(regs_185_clock),
    .reset(regs_185_reset),
    .io_in(regs_185_io_in),
    .io_reset(regs_185_io_reset),
    .io_out(regs_185_io_out),
    .io_enable(regs_185_io_enable)
  );
  FringeFF regs_186 ( // @[RegFile.scala 66:20:@52334.4]
    .clock(regs_186_clock),
    .reset(regs_186_reset),
    .io_in(regs_186_io_in),
    .io_reset(regs_186_io_reset),
    .io_out(regs_186_io_out),
    .io_enable(regs_186_io_enable)
  );
  FringeFF regs_187 ( // @[RegFile.scala 66:20:@52348.4]
    .clock(regs_187_clock),
    .reset(regs_187_reset),
    .io_in(regs_187_io_in),
    .io_reset(regs_187_io_reset),
    .io_out(regs_187_io_out),
    .io_enable(regs_187_io_enable)
  );
  FringeFF regs_188 ( // @[RegFile.scala 66:20:@52362.4]
    .clock(regs_188_clock),
    .reset(regs_188_reset),
    .io_in(regs_188_io_in),
    .io_reset(regs_188_io_reset),
    .io_out(regs_188_io_out),
    .io_enable(regs_188_io_enable)
  );
  FringeFF regs_189 ( // @[RegFile.scala 66:20:@52376.4]
    .clock(regs_189_clock),
    .reset(regs_189_reset),
    .io_in(regs_189_io_in),
    .io_reset(regs_189_io_reset),
    .io_out(regs_189_io_out),
    .io_enable(regs_189_io_enable)
  );
  FringeFF regs_190 ( // @[RegFile.scala 66:20:@52390.4]
    .clock(regs_190_clock),
    .reset(regs_190_reset),
    .io_in(regs_190_io_in),
    .io_reset(regs_190_io_reset),
    .io_out(regs_190_io_out),
    .io_enable(regs_190_io_enable)
  );
  FringeFF regs_191 ( // @[RegFile.scala 66:20:@52404.4]
    .clock(regs_191_clock),
    .reset(regs_191_reset),
    .io_in(regs_191_io_in),
    .io_reset(regs_191_io_reset),
    .io_out(regs_191_io_out),
    .io_enable(regs_191_io_enable)
  );
  FringeFF regs_192 ( // @[RegFile.scala 66:20:@52418.4]
    .clock(regs_192_clock),
    .reset(regs_192_reset),
    .io_in(regs_192_io_in),
    .io_reset(regs_192_io_reset),
    .io_out(regs_192_io_out),
    .io_enable(regs_192_io_enable)
  );
  FringeFF regs_193 ( // @[RegFile.scala 66:20:@52432.4]
    .clock(regs_193_clock),
    .reset(regs_193_reset),
    .io_in(regs_193_io_in),
    .io_reset(regs_193_io_reset),
    .io_out(regs_193_io_out),
    .io_enable(regs_193_io_enable)
  );
  FringeFF regs_194 ( // @[RegFile.scala 66:20:@52446.4]
    .clock(regs_194_clock),
    .reset(regs_194_reset),
    .io_in(regs_194_io_in),
    .io_reset(regs_194_io_reset),
    .io_out(regs_194_io_out),
    .io_enable(regs_194_io_enable)
  );
  FringeFF regs_195 ( // @[RegFile.scala 66:20:@52460.4]
    .clock(regs_195_clock),
    .reset(regs_195_reset),
    .io_in(regs_195_io_in),
    .io_reset(regs_195_io_reset),
    .io_out(regs_195_io_out),
    .io_enable(regs_195_io_enable)
  );
  FringeFF regs_196 ( // @[RegFile.scala 66:20:@52474.4]
    .clock(regs_196_clock),
    .reset(regs_196_reset),
    .io_in(regs_196_io_in),
    .io_reset(regs_196_io_reset),
    .io_out(regs_196_io_out),
    .io_enable(regs_196_io_enable)
  );
  FringeFF regs_197 ( // @[RegFile.scala 66:20:@52488.4]
    .clock(regs_197_clock),
    .reset(regs_197_reset),
    .io_in(regs_197_io_in),
    .io_reset(regs_197_io_reset),
    .io_out(regs_197_io_out),
    .io_enable(regs_197_io_enable)
  );
  FringeFF regs_198 ( // @[RegFile.scala 66:20:@52502.4]
    .clock(regs_198_clock),
    .reset(regs_198_reset),
    .io_in(regs_198_io_in),
    .io_reset(regs_198_io_reset),
    .io_out(regs_198_io_out),
    .io_enable(regs_198_io_enable)
  );
  FringeFF regs_199 ( // @[RegFile.scala 66:20:@52516.4]
    .clock(regs_199_clock),
    .reset(regs_199_reset),
    .io_in(regs_199_io_in),
    .io_reset(regs_199_io_reset),
    .io_out(regs_199_io_out),
    .io_enable(regs_199_io_enable)
  );
  FringeFF regs_200 ( // @[RegFile.scala 66:20:@52530.4]
    .clock(regs_200_clock),
    .reset(regs_200_reset),
    .io_in(regs_200_io_in),
    .io_reset(regs_200_io_reset),
    .io_out(regs_200_io_out),
    .io_enable(regs_200_io_enable)
  );
  FringeFF regs_201 ( // @[RegFile.scala 66:20:@52544.4]
    .clock(regs_201_clock),
    .reset(regs_201_reset),
    .io_in(regs_201_io_in),
    .io_reset(regs_201_io_reset),
    .io_out(regs_201_io_out),
    .io_enable(regs_201_io_enable)
  );
  FringeFF regs_202 ( // @[RegFile.scala 66:20:@52558.4]
    .clock(regs_202_clock),
    .reset(regs_202_reset),
    .io_in(regs_202_io_in),
    .io_reset(regs_202_io_reset),
    .io_out(regs_202_io_out),
    .io_enable(regs_202_io_enable)
  );
  FringeFF regs_203 ( // @[RegFile.scala 66:20:@52572.4]
    .clock(regs_203_clock),
    .reset(regs_203_reset),
    .io_in(regs_203_io_in),
    .io_reset(regs_203_io_reset),
    .io_out(regs_203_io_out),
    .io_enable(regs_203_io_enable)
  );
  FringeFF regs_204 ( // @[RegFile.scala 66:20:@52586.4]
    .clock(regs_204_clock),
    .reset(regs_204_reset),
    .io_in(regs_204_io_in),
    .io_reset(regs_204_io_reset),
    .io_out(regs_204_io_out),
    .io_enable(regs_204_io_enable)
  );
  FringeFF regs_205 ( // @[RegFile.scala 66:20:@52600.4]
    .clock(regs_205_clock),
    .reset(regs_205_reset),
    .io_in(regs_205_io_in),
    .io_reset(regs_205_io_reset),
    .io_out(regs_205_io_out),
    .io_enable(regs_205_io_enable)
  );
  FringeFF regs_206 ( // @[RegFile.scala 66:20:@52614.4]
    .clock(regs_206_clock),
    .reset(regs_206_reset),
    .io_in(regs_206_io_in),
    .io_reset(regs_206_io_reset),
    .io_out(regs_206_io_out),
    .io_enable(regs_206_io_enable)
  );
  FringeFF regs_207 ( // @[RegFile.scala 66:20:@52628.4]
    .clock(regs_207_clock),
    .reset(regs_207_reset),
    .io_in(regs_207_io_in),
    .io_reset(regs_207_io_reset),
    .io_out(regs_207_io_out),
    .io_enable(regs_207_io_enable)
  );
  FringeFF regs_208 ( // @[RegFile.scala 66:20:@52642.4]
    .clock(regs_208_clock),
    .reset(regs_208_reset),
    .io_in(regs_208_io_in),
    .io_reset(regs_208_io_reset),
    .io_out(regs_208_io_out),
    .io_enable(regs_208_io_enable)
  );
  FringeFF regs_209 ( // @[RegFile.scala 66:20:@52656.4]
    .clock(regs_209_clock),
    .reset(regs_209_reset),
    .io_in(regs_209_io_in),
    .io_reset(regs_209_io_reset),
    .io_out(regs_209_io_out),
    .io_enable(regs_209_io_enable)
  );
  FringeFF regs_210 ( // @[RegFile.scala 66:20:@52670.4]
    .clock(regs_210_clock),
    .reset(regs_210_reset),
    .io_in(regs_210_io_in),
    .io_reset(regs_210_io_reset),
    .io_out(regs_210_io_out),
    .io_enable(regs_210_io_enable)
  );
  FringeFF regs_211 ( // @[RegFile.scala 66:20:@52684.4]
    .clock(regs_211_clock),
    .reset(regs_211_reset),
    .io_in(regs_211_io_in),
    .io_reset(regs_211_io_reset),
    .io_out(regs_211_io_out),
    .io_enable(regs_211_io_enable)
  );
  FringeFF regs_212 ( // @[RegFile.scala 66:20:@52698.4]
    .clock(regs_212_clock),
    .reset(regs_212_reset),
    .io_in(regs_212_io_in),
    .io_reset(regs_212_io_reset),
    .io_out(regs_212_io_out),
    .io_enable(regs_212_io_enable)
  );
  FringeFF regs_213 ( // @[RegFile.scala 66:20:@52712.4]
    .clock(regs_213_clock),
    .reset(regs_213_reset),
    .io_in(regs_213_io_in),
    .io_reset(regs_213_io_reset),
    .io_out(regs_213_io_out),
    .io_enable(regs_213_io_enable)
  );
  FringeFF regs_214 ( // @[RegFile.scala 66:20:@52726.4]
    .clock(regs_214_clock),
    .reset(regs_214_reset),
    .io_in(regs_214_io_in),
    .io_reset(regs_214_io_reset),
    .io_out(regs_214_io_out),
    .io_enable(regs_214_io_enable)
  );
  FringeFF regs_215 ( // @[RegFile.scala 66:20:@52740.4]
    .clock(regs_215_clock),
    .reset(regs_215_reset),
    .io_in(regs_215_io_in),
    .io_reset(regs_215_io_reset),
    .io_out(regs_215_io_out),
    .io_enable(regs_215_io_enable)
  );
  FringeFF regs_216 ( // @[RegFile.scala 66:20:@52754.4]
    .clock(regs_216_clock),
    .reset(regs_216_reset),
    .io_in(regs_216_io_in),
    .io_reset(regs_216_io_reset),
    .io_out(regs_216_io_out),
    .io_enable(regs_216_io_enable)
  );
  FringeFF regs_217 ( // @[RegFile.scala 66:20:@52768.4]
    .clock(regs_217_clock),
    .reset(regs_217_reset),
    .io_in(regs_217_io_in),
    .io_reset(regs_217_io_reset),
    .io_out(regs_217_io_out),
    .io_enable(regs_217_io_enable)
  );
  FringeFF regs_218 ( // @[RegFile.scala 66:20:@52782.4]
    .clock(regs_218_clock),
    .reset(regs_218_reset),
    .io_in(regs_218_io_in),
    .io_reset(regs_218_io_reset),
    .io_out(regs_218_io_out),
    .io_enable(regs_218_io_enable)
  );
  FringeFF regs_219 ( // @[RegFile.scala 66:20:@52796.4]
    .clock(regs_219_clock),
    .reset(regs_219_reset),
    .io_in(regs_219_io_in),
    .io_reset(regs_219_io_reset),
    .io_out(regs_219_io_out),
    .io_enable(regs_219_io_enable)
  );
  FringeFF regs_220 ( // @[RegFile.scala 66:20:@52810.4]
    .clock(regs_220_clock),
    .reset(regs_220_reset),
    .io_in(regs_220_io_in),
    .io_reset(regs_220_io_reset),
    .io_out(regs_220_io_out),
    .io_enable(regs_220_io_enable)
  );
  FringeFF regs_221 ( // @[RegFile.scala 66:20:@52824.4]
    .clock(regs_221_clock),
    .reset(regs_221_reset),
    .io_in(regs_221_io_in),
    .io_reset(regs_221_io_reset),
    .io_out(regs_221_io_out),
    .io_enable(regs_221_io_enable)
  );
  FringeFF regs_222 ( // @[RegFile.scala 66:20:@52838.4]
    .clock(regs_222_clock),
    .reset(regs_222_reset),
    .io_in(regs_222_io_in),
    .io_reset(regs_222_io_reset),
    .io_out(regs_222_io_out),
    .io_enable(regs_222_io_enable)
  );
  FringeFF regs_223 ( // @[RegFile.scala 66:20:@52852.4]
    .clock(regs_223_clock),
    .reset(regs_223_reset),
    .io_in(regs_223_io_in),
    .io_reset(regs_223_io_reset),
    .io_out(regs_223_io_out),
    .io_enable(regs_223_io_enable)
  );
  FringeFF regs_224 ( // @[RegFile.scala 66:20:@52866.4]
    .clock(regs_224_clock),
    .reset(regs_224_reset),
    .io_in(regs_224_io_in),
    .io_reset(regs_224_io_reset),
    .io_out(regs_224_io_out),
    .io_enable(regs_224_io_enable)
  );
  FringeFF regs_225 ( // @[RegFile.scala 66:20:@52880.4]
    .clock(regs_225_clock),
    .reset(regs_225_reset),
    .io_in(regs_225_io_in),
    .io_reset(regs_225_io_reset),
    .io_out(regs_225_io_out),
    .io_enable(regs_225_io_enable)
  );
  FringeFF regs_226 ( // @[RegFile.scala 66:20:@52894.4]
    .clock(regs_226_clock),
    .reset(regs_226_reset),
    .io_in(regs_226_io_in),
    .io_reset(regs_226_io_reset),
    .io_out(regs_226_io_out),
    .io_enable(regs_226_io_enable)
  );
  FringeFF regs_227 ( // @[RegFile.scala 66:20:@52908.4]
    .clock(regs_227_clock),
    .reset(regs_227_reset),
    .io_in(regs_227_io_in),
    .io_reset(regs_227_io_reset),
    .io_out(regs_227_io_out),
    .io_enable(regs_227_io_enable)
  );
  FringeFF regs_228 ( // @[RegFile.scala 66:20:@52922.4]
    .clock(regs_228_clock),
    .reset(regs_228_reset),
    .io_in(regs_228_io_in),
    .io_reset(regs_228_io_reset),
    .io_out(regs_228_io_out),
    .io_enable(regs_228_io_enable)
  );
  FringeFF regs_229 ( // @[RegFile.scala 66:20:@52936.4]
    .clock(regs_229_clock),
    .reset(regs_229_reset),
    .io_in(regs_229_io_in),
    .io_reset(regs_229_io_reset),
    .io_out(regs_229_io_out),
    .io_enable(regs_229_io_enable)
  );
  FringeFF regs_230 ( // @[RegFile.scala 66:20:@52950.4]
    .clock(regs_230_clock),
    .reset(regs_230_reset),
    .io_in(regs_230_io_in),
    .io_reset(regs_230_io_reset),
    .io_out(regs_230_io_out),
    .io_enable(regs_230_io_enable)
  );
  FringeFF regs_231 ( // @[RegFile.scala 66:20:@52964.4]
    .clock(regs_231_clock),
    .reset(regs_231_reset),
    .io_in(regs_231_io_in),
    .io_reset(regs_231_io_reset),
    .io_out(regs_231_io_out),
    .io_enable(regs_231_io_enable)
  );
  FringeFF regs_232 ( // @[RegFile.scala 66:20:@52978.4]
    .clock(regs_232_clock),
    .reset(regs_232_reset),
    .io_in(regs_232_io_in),
    .io_reset(regs_232_io_reset),
    .io_out(regs_232_io_out),
    .io_enable(regs_232_io_enable)
  );
  FringeFF regs_233 ( // @[RegFile.scala 66:20:@52992.4]
    .clock(regs_233_clock),
    .reset(regs_233_reset),
    .io_in(regs_233_io_in),
    .io_reset(regs_233_io_reset),
    .io_out(regs_233_io_out),
    .io_enable(regs_233_io_enable)
  );
  FringeFF regs_234 ( // @[RegFile.scala 66:20:@53006.4]
    .clock(regs_234_clock),
    .reset(regs_234_reset),
    .io_in(regs_234_io_in),
    .io_reset(regs_234_io_reset),
    .io_out(regs_234_io_out),
    .io_enable(regs_234_io_enable)
  );
  FringeFF regs_235 ( // @[RegFile.scala 66:20:@53020.4]
    .clock(regs_235_clock),
    .reset(regs_235_reset),
    .io_in(regs_235_io_in),
    .io_reset(regs_235_io_reset),
    .io_out(regs_235_io_out),
    .io_enable(regs_235_io_enable)
  );
  FringeFF regs_236 ( // @[RegFile.scala 66:20:@53034.4]
    .clock(regs_236_clock),
    .reset(regs_236_reset),
    .io_in(regs_236_io_in),
    .io_reset(regs_236_io_reset),
    .io_out(regs_236_io_out),
    .io_enable(regs_236_io_enable)
  );
  FringeFF regs_237 ( // @[RegFile.scala 66:20:@53048.4]
    .clock(regs_237_clock),
    .reset(regs_237_reset),
    .io_in(regs_237_io_in),
    .io_reset(regs_237_io_reset),
    .io_out(regs_237_io_out),
    .io_enable(regs_237_io_enable)
  );
  FringeFF regs_238 ( // @[RegFile.scala 66:20:@53062.4]
    .clock(regs_238_clock),
    .reset(regs_238_reset),
    .io_in(regs_238_io_in),
    .io_reset(regs_238_io_reset),
    .io_out(regs_238_io_out),
    .io_enable(regs_238_io_enable)
  );
  FringeFF regs_239 ( // @[RegFile.scala 66:20:@53076.4]
    .clock(regs_239_clock),
    .reset(regs_239_reset),
    .io_in(regs_239_io_in),
    .io_reset(regs_239_io_reset),
    .io_out(regs_239_io_out),
    .io_enable(regs_239_io_enable)
  );
  FringeFF regs_240 ( // @[RegFile.scala 66:20:@53090.4]
    .clock(regs_240_clock),
    .reset(regs_240_reset),
    .io_in(regs_240_io_in),
    .io_reset(regs_240_io_reset),
    .io_out(regs_240_io_out),
    .io_enable(regs_240_io_enable)
  );
  FringeFF regs_241 ( // @[RegFile.scala 66:20:@53104.4]
    .clock(regs_241_clock),
    .reset(regs_241_reset),
    .io_in(regs_241_io_in),
    .io_reset(regs_241_io_reset),
    .io_out(regs_241_io_out),
    .io_enable(regs_241_io_enable)
  );
  FringeFF regs_242 ( // @[RegFile.scala 66:20:@53118.4]
    .clock(regs_242_clock),
    .reset(regs_242_reset),
    .io_in(regs_242_io_in),
    .io_reset(regs_242_io_reset),
    .io_out(regs_242_io_out),
    .io_enable(regs_242_io_enable)
  );
  FringeFF regs_243 ( // @[RegFile.scala 66:20:@53132.4]
    .clock(regs_243_clock),
    .reset(regs_243_reset),
    .io_in(regs_243_io_in),
    .io_reset(regs_243_io_reset),
    .io_out(regs_243_io_out),
    .io_enable(regs_243_io_enable)
  );
  FringeFF regs_244 ( // @[RegFile.scala 66:20:@53146.4]
    .clock(regs_244_clock),
    .reset(regs_244_reset),
    .io_in(regs_244_io_in),
    .io_reset(regs_244_io_reset),
    .io_out(regs_244_io_out),
    .io_enable(regs_244_io_enable)
  );
  FringeFF regs_245 ( // @[RegFile.scala 66:20:@53160.4]
    .clock(regs_245_clock),
    .reset(regs_245_reset),
    .io_in(regs_245_io_in),
    .io_reset(regs_245_io_reset),
    .io_out(regs_245_io_out),
    .io_enable(regs_245_io_enable)
  );
  FringeFF regs_246 ( // @[RegFile.scala 66:20:@53174.4]
    .clock(regs_246_clock),
    .reset(regs_246_reset),
    .io_in(regs_246_io_in),
    .io_reset(regs_246_io_reset),
    .io_out(regs_246_io_out),
    .io_enable(regs_246_io_enable)
  );
  FringeFF regs_247 ( // @[RegFile.scala 66:20:@53188.4]
    .clock(regs_247_clock),
    .reset(regs_247_reset),
    .io_in(regs_247_io_in),
    .io_reset(regs_247_io_reset),
    .io_out(regs_247_io_out),
    .io_enable(regs_247_io_enable)
  );
  FringeFF regs_248 ( // @[RegFile.scala 66:20:@53202.4]
    .clock(regs_248_clock),
    .reset(regs_248_reset),
    .io_in(regs_248_io_in),
    .io_reset(regs_248_io_reset),
    .io_out(regs_248_io_out),
    .io_enable(regs_248_io_enable)
  );
  FringeFF regs_249 ( // @[RegFile.scala 66:20:@53216.4]
    .clock(regs_249_clock),
    .reset(regs_249_reset),
    .io_in(regs_249_io_in),
    .io_reset(regs_249_io_reset),
    .io_out(regs_249_io_out),
    .io_enable(regs_249_io_enable)
  );
  FringeFF regs_250 ( // @[RegFile.scala 66:20:@53230.4]
    .clock(regs_250_clock),
    .reset(regs_250_reset),
    .io_in(regs_250_io_in),
    .io_reset(regs_250_io_reset),
    .io_out(regs_250_io_out),
    .io_enable(regs_250_io_enable)
  );
  FringeFF regs_251 ( // @[RegFile.scala 66:20:@53244.4]
    .clock(regs_251_clock),
    .reset(regs_251_reset),
    .io_in(regs_251_io_in),
    .io_reset(regs_251_io_reset),
    .io_out(regs_251_io_out),
    .io_enable(regs_251_io_enable)
  );
  FringeFF regs_252 ( // @[RegFile.scala 66:20:@53258.4]
    .clock(regs_252_clock),
    .reset(regs_252_reset),
    .io_in(regs_252_io_in),
    .io_reset(regs_252_io_reset),
    .io_out(regs_252_io_out),
    .io_enable(regs_252_io_enable)
  );
  FringeFF regs_253 ( // @[RegFile.scala 66:20:@53272.4]
    .clock(regs_253_clock),
    .reset(regs_253_reset),
    .io_in(regs_253_io_in),
    .io_reset(regs_253_io_reset),
    .io_out(regs_253_io_out),
    .io_enable(regs_253_io_enable)
  );
  FringeFF regs_254 ( // @[RegFile.scala 66:20:@53286.4]
    .clock(regs_254_clock),
    .reset(regs_254_reset),
    .io_in(regs_254_io_in),
    .io_reset(regs_254_io_reset),
    .io_out(regs_254_io_out),
    .io_enable(regs_254_io_enable)
  );
  FringeFF regs_255 ( // @[RegFile.scala 66:20:@53300.4]
    .clock(regs_255_clock),
    .reset(regs_255_reset),
    .io_in(regs_255_io_in),
    .io_reset(regs_255_io_reset),
    .io_out(regs_255_io_out),
    .io_enable(regs_255_io_enable)
  );
  FringeFF regs_256 ( // @[RegFile.scala 66:20:@53314.4]
    .clock(regs_256_clock),
    .reset(regs_256_reset),
    .io_in(regs_256_io_in),
    .io_reset(regs_256_io_reset),
    .io_out(regs_256_io_out),
    .io_enable(regs_256_io_enable)
  );
  FringeFF regs_257 ( // @[RegFile.scala 66:20:@53328.4]
    .clock(regs_257_clock),
    .reset(regs_257_reset),
    .io_in(regs_257_io_in),
    .io_reset(regs_257_io_reset),
    .io_out(regs_257_io_out),
    .io_enable(regs_257_io_enable)
  );
  FringeFF regs_258 ( // @[RegFile.scala 66:20:@53342.4]
    .clock(regs_258_clock),
    .reset(regs_258_reset),
    .io_in(regs_258_io_in),
    .io_reset(regs_258_io_reset),
    .io_out(regs_258_io_out),
    .io_enable(regs_258_io_enable)
  );
  FringeFF regs_259 ( // @[RegFile.scala 66:20:@53356.4]
    .clock(regs_259_clock),
    .reset(regs_259_reset),
    .io_in(regs_259_io_in),
    .io_reset(regs_259_io_reset),
    .io_out(regs_259_io_out),
    .io_enable(regs_259_io_enable)
  );
  FringeFF regs_260 ( // @[RegFile.scala 66:20:@53370.4]
    .clock(regs_260_clock),
    .reset(regs_260_reset),
    .io_in(regs_260_io_in),
    .io_reset(regs_260_io_reset),
    .io_out(regs_260_io_out),
    .io_enable(regs_260_io_enable)
  );
  FringeFF regs_261 ( // @[RegFile.scala 66:20:@53384.4]
    .clock(regs_261_clock),
    .reset(regs_261_reset),
    .io_in(regs_261_io_in),
    .io_reset(regs_261_io_reset),
    .io_out(regs_261_io_out),
    .io_enable(regs_261_io_enable)
  );
  FringeFF regs_262 ( // @[RegFile.scala 66:20:@53398.4]
    .clock(regs_262_clock),
    .reset(regs_262_reset),
    .io_in(regs_262_io_in),
    .io_reset(regs_262_io_reset),
    .io_out(regs_262_io_out),
    .io_enable(regs_262_io_enable)
  );
  FringeFF regs_263 ( // @[RegFile.scala 66:20:@53412.4]
    .clock(regs_263_clock),
    .reset(regs_263_reset),
    .io_in(regs_263_io_in),
    .io_reset(regs_263_io_reset),
    .io_out(regs_263_io_out),
    .io_enable(regs_263_io_enable)
  );
  FringeFF regs_264 ( // @[RegFile.scala 66:20:@53426.4]
    .clock(regs_264_clock),
    .reset(regs_264_reset),
    .io_in(regs_264_io_in),
    .io_reset(regs_264_io_reset),
    .io_out(regs_264_io_out),
    .io_enable(regs_264_io_enable)
  );
  FringeFF regs_265 ( // @[RegFile.scala 66:20:@53440.4]
    .clock(regs_265_clock),
    .reset(regs_265_reset),
    .io_in(regs_265_io_in),
    .io_reset(regs_265_io_reset),
    .io_out(regs_265_io_out),
    .io_enable(regs_265_io_enable)
  );
  FringeFF regs_266 ( // @[RegFile.scala 66:20:@53454.4]
    .clock(regs_266_clock),
    .reset(regs_266_reset),
    .io_in(regs_266_io_in),
    .io_reset(regs_266_io_reset),
    .io_out(regs_266_io_out),
    .io_enable(regs_266_io_enable)
  );
  FringeFF regs_267 ( // @[RegFile.scala 66:20:@53468.4]
    .clock(regs_267_clock),
    .reset(regs_267_reset),
    .io_in(regs_267_io_in),
    .io_reset(regs_267_io_reset),
    .io_out(regs_267_io_out),
    .io_enable(regs_267_io_enable)
  );
  FringeFF regs_268 ( // @[RegFile.scala 66:20:@53482.4]
    .clock(regs_268_clock),
    .reset(regs_268_reset),
    .io_in(regs_268_io_in),
    .io_reset(regs_268_io_reset),
    .io_out(regs_268_io_out),
    .io_enable(regs_268_io_enable)
  );
  FringeFF regs_269 ( // @[RegFile.scala 66:20:@53496.4]
    .clock(regs_269_clock),
    .reset(regs_269_reset),
    .io_in(regs_269_io_in),
    .io_reset(regs_269_io_reset),
    .io_out(regs_269_io_out),
    .io_enable(regs_269_io_enable)
  );
  FringeFF regs_270 ( // @[RegFile.scala 66:20:@53510.4]
    .clock(regs_270_clock),
    .reset(regs_270_reset),
    .io_in(regs_270_io_in),
    .io_reset(regs_270_io_reset),
    .io_out(regs_270_io_out),
    .io_enable(regs_270_io_enable)
  );
  FringeFF regs_271 ( // @[RegFile.scala 66:20:@53524.4]
    .clock(regs_271_clock),
    .reset(regs_271_reset),
    .io_in(regs_271_io_in),
    .io_reset(regs_271_io_reset),
    .io_out(regs_271_io_out),
    .io_enable(regs_271_io_enable)
  );
  FringeFF regs_272 ( // @[RegFile.scala 66:20:@53538.4]
    .clock(regs_272_clock),
    .reset(regs_272_reset),
    .io_in(regs_272_io_in),
    .io_reset(regs_272_io_reset),
    .io_out(regs_272_io_out),
    .io_enable(regs_272_io_enable)
  );
  FringeFF regs_273 ( // @[RegFile.scala 66:20:@53552.4]
    .clock(regs_273_clock),
    .reset(regs_273_reset),
    .io_in(regs_273_io_in),
    .io_reset(regs_273_io_reset),
    .io_out(regs_273_io_out),
    .io_enable(regs_273_io_enable)
  );
  FringeFF regs_274 ( // @[RegFile.scala 66:20:@53566.4]
    .clock(regs_274_clock),
    .reset(regs_274_reset),
    .io_in(regs_274_io_in),
    .io_reset(regs_274_io_reset),
    .io_out(regs_274_io_out),
    .io_enable(regs_274_io_enable)
  );
  FringeFF regs_275 ( // @[RegFile.scala 66:20:@53580.4]
    .clock(regs_275_clock),
    .reset(regs_275_reset),
    .io_in(regs_275_io_in),
    .io_reset(regs_275_io_reset),
    .io_out(regs_275_io_out),
    .io_enable(regs_275_io_enable)
  );
  FringeFF regs_276 ( // @[RegFile.scala 66:20:@53594.4]
    .clock(regs_276_clock),
    .reset(regs_276_reset),
    .io_in(regs_276_io_in),
    .io_reset(regs_276_io_reset),
    .io_out(regs_276_io_out),
    .io_enable(regs_276_io_enable)
  );
  FringeFF regs_277 ( // @[RegFile.scala 66:20:@53608.4]
    .clock(regs_277_clock),
    .reset(regs_277_reset),
    .io_in(regs_277_io_in),
    .io_reset(regs_277_io_reset),
    .io_out(regs_277_io_out),
    .io_enable(regs_277_io_enable)
  );
  FringeFF regs_278 ( // @[RegFile.scala 66:20:@53622.4]
    .clock(regs_278_clock),
    .reset(regs_278_reset),
    .io_in(regs_278_io_in),
    .io_reset(regs_278_io_reset),
    .io_out(regs_278_io_out),
    .io_enable(regs_278_io_enable)
  );
  FringeFF regs_279 ( // @[RegFile.scala 66:20:@53636.4]
    .clock(regs_279_clock),
    .reset(regs_279_reset),
    .io_in(regs_279_io_in),
    .io_reset(regs_279_io_reset),
    .io_out(regs_279_io_out),
    .io_enable(regs_279_io_enable)
  );
  FringeFF regs_280 ( // @[RegFile.scala 66:20:@53650.4]
    .clock(regs_280_clock),
    .reset(regs_280_reset),
    .io_in(regs_280_io_in),
    .io_reset(regs_280_io_reset),
    .io_out(regs_280_io_out),
    .io_enable(regs_280_io_enable)
  );
  FringeFF regs_281 ( // @[RegFile.scala 66:20:@53664.4]
    .clock(regs_281_clock),
    .reset(regs_281_reset),
    .io_in(regs_281_io_in),
    .io_reset(regs_281_io_reset),
    .io_out(regs_281_io_out),
    .io_enable(regs_281_io_enable)
  );
  FringeFF regs_282 ( // @[RegFile.scala 66:20:@53678.4]
    .clock(regs_282_clock),
    .reset(regs_282_reset),
    .io_in(regs_282_io_in),
    .io_reset(regs_282_io_reset),
    .io_out(regs_282_io_out),
    .io_enable(regs_282_io_enable)
  );
  FringeFF regs_283 ( // @[RegFile.scala 66:20:@53692.4]
    .clock(regs_283_clock),
    .reset(regs_283_reset),
    .io_in(regs_283_io_in),
    .io_reset(regs_283_io_reset),
    .io_out(regs_283_io_out),
    .io_enable(regs_283_io_enable)
  );
  FringeFF regs_284 ( // @[RegFile.scala 66:20:@53706.4]
    .clock(regs_284_clock),
    .reset(regs_284_reset),
    .io_in(regs_284_io_in),
    .io_reset(regs_284_io_reset),
    .io_out(regs_284_io_out),
    .io_enable(regs_284_io_enable)
  );
  FringeFF regs_285 ( // @[RegFile.scala 66:20:@53720.4]
    .clock(regs_285_clock),
    .reset(regs_285_reset),
    .io_in(regs_285_io_in),
    .io_reset(regs_285_io_reset),
    .io_out(regs_285_io_out),
    .io_enable(regs_285_io_enable)
  );
  FringeFF regs_286 ( // @[RegFile.scala 66:20:@53734.4]
    .clock(regs_286_clock),
    .reset(regs_286_reset),
    .io_in(regs_286_io_in),
    .io_reset(regs_286_io_reset),
    .io_out(regs_286_io_out),
    .io_enable(regs_286_io_enable)
  );
  FringeFF regs_287 ( // @[RegFile.scala 66:20:@53748.4]
    .clock(regs_287_clock),
    .reset(regs_287_reset),
    .io_in(regs_287_io_in),
    .io_reset(regs_287_io_reset),
    .io_out(regs_287_io_out),
    .io_enable(regs_287_io_enable)
  );
  FringeFF regs_288 ( // @[RegFile.scala 66:20:@53762.4]
    .clock(regs_288_clock),
    .reset(regs_288_reset),
    .io_in(regs_288_io_in),
    .io_reset(regs_288_io_reset),
    .io_out(regs_288_io_out),
    .io_enable(regs_288_io_enable)
  );
  FringeFF regs_289 ( // @[RegFile.scala 66:20:@53776.4]
    .clock(regs_289_clock),
    .reset(regs_289_reset),
    .io_in(regs_289_io_in),
    .io_reset(regs_289_io_reset),
    .io_out(regs_289_io_out),
    .io_enable(regs_289_io_enable)
  );
  FringeFF regs_290 ( // @[RegFile.scala 66:20:@53790.4]
    .clock(regs_290_clock),
    .reset(regs_290_reset),
    .io_in(regs_290_io_in),
    .io_reset(regs_290_io_reset),
    .io_out(regs_290_io_out),
    .io_enable(regs_290_io_enable)
  );
  FringeFF regs_291 ( // @[RegFile.scala 66:20:@53804.4]
    .clock(regs_291_clock),
    .reset(regs_291_reset),
    .io_in(regs_291_io_in),
    .io_reset(regs_291_io_reset),
    .io_out(regs_291_io_out),
    .io_enable(regs_291_io_enable)
  );
  FringeFF regs_292 ( // @[RegFile.scala 66:20:@53818.4]
    .clock(regs_292_clock),
    .reset(regs_292_reset),
    .io_in(regs_292_io_in),
    .io_reset(regs_292_io_reset),
    .io_out(regs_292_io_out),
    .io_enable(regs_292_io_enable)
  );
  FringeFF regs_293 ( // @[RegFile.scala 66:20:@53832.4]
    .clock(regs_293_clock),
    .reset(regs_293_reset),
    .io_in(regs_293_io_in),
    .io_reset(regs_293_io_reset),
    .io_out(regs_293_io_out),
    .io_enable(regs_293_io_enable)
  );
  FringeFF regs_294 ( // @[RegFile.scala 66:20:@53846.4]
    .clock(regs_294_clock),
    .reset(regs_294_reset),
    .io_in(regs_294_io_in),
    .io_reset(regs_294_io_reset),
    .io_out(regs_294_io_out),
    .io_enable(regs_294_io_enable)
  );
  FringeFF regs_295 ( // @[RegFile.scala 66:20:@53860.4]
    .clock(regs_295_clock),
    .reset(regs_295_reset),
    .io_in(regs_295_io_in),
    .io_reset(regs_295_io_reset),
    .io_out(regs_295_io_out),
    .io_enable(regs_295_io_enable)
  );
  FringeFF regs_296 ( // @[RegFile.scala 66:20:@53874.4]
    .clock(regs_296_clock),
    .reset(regs_296_reset),
    .io_in(regs_296_io_in),
    .io_reset(regs_296_io_reset),
    .io_out(regs_296_io_out),
    .io_enable(regs_296_io_enable)
  );
  FringeFF regs_297 ( // @[RegFile.scala 66:20:@53888.4]
    .clock(regs_297_clock),
    .reset(regs_297_reset),
    .io_in(regs_297_io_in),
    .io_reset(regs_297_io_reset),
    .io_out(regs_297_io_out),
    .io_enable(regs_297_io_enable)
  );
  FringeFF regs_298 ( // @[RegFile.scala 66:20:@53902.4]
    .clock(regs_298_clock),
    .reset(regs_298_reset),
    .io_in(regs_298_io_in),
    .io_reset(regs_298_io_reset),
    .io_out(regs_298_io_out),
    .io_enable(regs_298_io_enable)
  );
  FringeFF regs_299 ( // @[RegFile.scala 66:20:@53916.4]
    .clock(regs_299_clock),
    .reset(regs_299_reset),
    .io_in(regs_299_io_in),
    .io_reset(regs_299_io_reset),
    .io_out(regs_299_io_out),
    .io_enable(regs_299_io_enable)
  );
  FringeFF regs_300 ( // @[RegFile.scala 66:20:@53930.4]
    .clock(regs_300_clock),
    .reset(regs_300_reset),
    .io_in(regs_300_io_in),
    .io_reset(regs_300_io_reset),
    .io_out(regs_300_io_out),
    .io_enable(regs_300_io_enable)
  );
  FringeFF regs_301 ( // @[RegFile.scala 66:20:@53944.4]
    .clock(regs_301_clock),
    .reset(regs_301_reset),
    .io_in(regs_301_io_in),
    .io_reset(regs_301_io_reset),
    .io_out(regs_301_io_out),
    .io_enable(regs_301_io_enable)
  );
  FringeFF regs_302 ( // @[RegFile.scala 66:20:@53958.4]
    .clock(regs_302_clock),
    .reset(regs_302_reset),
    .io_in(regs_302_io_in),
    .io_reset(regs_302_io_reset),
    .io_out(regs_302_io_out),
    .io_enable(regs_302_io_enable)
  );
  FringeFF regs_303 ( // @[RegFile.scala 66:20:@53972.4]
    .clock(regs_303_clock),
    .reset(regs_303_reset),
    .io_in(regs_303_io_in),
    .io_reset(regs_303_io_reset),
    .io_out(regs_303_io_out),
    .io_enable(regs_303_io_enable)
  );
  FringeFF regs_304 ( // @[RegFile.scala 66:20:@53986.4]
    .clock(regs_304_clock),
    .reset(regs_304_reset),
    .io_in(regs_304_io_in),
    .io_reset(regs_304_io_reset),
    .io_out(regs_304_io_out),
    .io_enable(regs_304_io_enable)
  );
  FringeFF regs_305 ( // @[RegFile.scala 66:20:@54000.4]
    .clock(regs_305_clock),
    .reset(regs_305_reset),
    .io_in(regs_305_io_in),
    .io_reset(regs_305_io_reset),
    .io_out(regs_305_io_out),
    .io_enable(regs_305_io_enable)
  );
  FringeFF regs_306 ( // @[RegFile.scala 66:20:@54014.4]
    .clock(regs_306_clock),
    .reset(regs_306_reset),
    .io_in(regs_306_io_in),
    .io_reset(regs_306_io_reset),
    .io_out(regs_306_io_out),
    .io_enable(regs_306_io_enable)
  );
  FringeFF regs_307 ( // @[RegFile.scala 66:20:@54028.4]
    .clock(regs_307_clock),
    .reset(regs_307_reset),
    .io_in(regs_307_io_in),
    .io_reset(regs_307_io_reset),
    .io_out(regs_307_io_out),
    .io_enable(regs_307_io_enable)
  );
  FringeFF regs_308 ( // @[RegFile.scala 66:20:@54042.4]
    .clock(regs_308_clock),
    .reset(regs_308_reset),
    .io_in(regs_308_io_in),
    .io_reset(regs_308_io_reset),
    .io_out(regs_308_io_out),
    .io_enable(regs_308_io_enable)
  );
  FringeFF regs_309 ( // @[RegFile.scala 66:20:@54056.4]
    .clock(regs_309_clock),
    .reset(regs_309_reset),
    .io_in(regs_309_io_in),
    .io_reset(regs_309_io_reset),
    .io_out(regs_309_io_out),
    .io_enable(regs_309_io_enable)
  );
  FringeFF regs_310 ( // @[RegFile.scala 66:20:@54070.4]
    .clock(regs_310_clock),
    .reset(regs_310_reset),
    .io_in(regs_310_io_in),
    .io_reset(regs_310_io_reset),
    .io_out(regs_310_io_out),
    .io_enable(regs_310_io_enable)
  );
  FringeFF regs_311 ( // @[RegFile.scala 66:20:@54084.4]
    .clock(regs_311_clock),
    .reset(regs_311_reset),
    .io_in(regs_311_io_in),
    .io_reset(regs_311_io_reset),
    .io_out(regs_311_io_out),
    .io_enable(regs_311_io_enable)
  );
  FringeFF regs_312 ( // @[RegFile.scala 66:20:@54098.4]
    .clock(regs_312_clock),
    .reset(regs_312_reset),
    .io_in(regs_312_io_in),
    .io_reset(regs_312_io_reset),
    .io_out(regs_312_io_out),
    .io_enable(regs_312_io_enable)
  );
  FringeFF regs_313 ( // @[RegFile.scala 66:20:@54112.4]
    .clock(regs_313_clock),
    .reset(regs_313_reset),
    .io_in(regs_313_io_in),
    .io_reset(regs_313_io_reset),
    .io_out(regs_313_io_out),
    .io_enable(regs_313_io_enable)
  );
  FringeFF regs_314 ( // @[RegFile.scala 66:20:@54126.4]
    .clock(regs_314_clock),
    .reset(regs_314_reset),
    .io_in(regs_314_io_in),
    .io_reset(regs_314_io_reset),
    .io_out(regs_314_io_out),
    .io_enable(regs_314_io_enable)
  );
  FringeFF regs_315 ( // @[RegFile.scala 66:20:@54140.4]
    .clock(regs_315_clock),
    .reset(regs_315_reset),
    .io_in(regs_315_io_in),
    .io_reset(regs_315_io_reset),
    .io_out(regs_315_io_out),
    .io_enable(regs_315_io_enable)
  );
  FringeFF regs_316 ( // @[RegFile.scala 66:20:@54154.4]
    .clock(regs_316_clock),
    .reset(regs_316_reset),
    .io_in(regs_316_io_in),
    .io_reset(regs_316_io_reset),
    .io_out(regs_316_io_out),
    .io_enable(regs_316_io_enable)
  );
  FringeFF regs_317 ( // @[RegFile.scala 66:20:@54168.4]
    .clock(regs_317_clock),
    .reset(regs_317_reset),
    .io_in(regs_317_io_in),
    .io_reset(regs_317_io_reset),
    .io_out(regs_317_io_out),
    .io_enable(regs_317_io_enable)
  );
  FringeFF regs_318 ( // @[RegFile.scala 66:20:@54182.4]
    .clock(regs_318_clock),
    .reset(regs_318_reset),
    .io_in(regs_318_io_in),
    .io_reset(regs_318_io_reset),
    .io_out(regs_318_io_out),
    .io_enable(regs_318_io_enable)
  );
  FringeFF regs_319 ( // @[RegFile.scala 66:20:@54196.4]
    .clock(regs_319_clock),
    .reset(regs_319_reset),
    .io_in(regs_319_io_in),
    .io_reset(regs_319_io_reset),
    .io_out(regs_319_io_out),
    .io_enable(regs_319_io_enable)
  );
  FringeFF regs_320 ( // @[RegFile.scala 66:20:@54210.4]
    .clock(regs_320_clock),
    .reset(regs_320_reset),
    .io_in(regs_320_io_in),
    .io_reset(regs_320_io_reset),
    .io_out(regs_320_io_out),
    .io_enable(regs_320_io_enable)
  );
  FringeFF regs_321 ( // @[RegFile.scala 66:20:@54224.4]
    .clock(regs_321_clock),
    .reset(regs_321_reset),
    .io_in(regs_321_io_in),
    .io_reset(regs_321_io_reset),
    .io_out(regs_321_io_out),
    .io_enable(regs_321_io_enable)
  );
  FringeFF regs_322 ( // @[RegFile.scala 66:20:@54238.4]
    .clock(regs_322_clock),
    .reset(regs_322_reset),
    .io_in(regs_322_io_in),
    .io_reset(regs_322_io_reset),
    .io_out(regs_322_io_out),
    .io_enable(regs_322_io_enable)
  );
  FringeFF regs_323 ( // @[RegFile.scala 66:20:@54252.4]
    .clock(regs_323_clock),
    .reset(regs_323_reset),
    .io_in(regs_323_io_in),
    .io_reset(regs_323_io_reset),
    .io_out(regs_323_io_out),
    .io_enable(regs_323_io_enable)
  );
  FringeFF regs_324 ( // @[RegFile.scala 66:20:@54266.4]
    .clock(regs_324_clock),
    .reset(regs_324_reset),
    .io_in(regs_324_io_in),
    .io_reset(regs_324_io_reset),
    .io_out(regs_324_io_out),
    .io_enable(regs_324_io_enable)
  );
  FringeFF regs_325 ( // @[RegFile.scala 66:20:@54280.4]
    .clock(regs_325_clock),
    .reset(regs_325_reset),
    .io_in(regs_325_io_in),
    .io_reset(regs_325_io_reset),
    .io_out(regs_325_io_out),
    .io_enable(regs_325_io_enable)
  );
  FringeFF regs_326 ( // @[RegFile.scala 66:20:@54294.4]
    .clock(regs_326_clock),
    .reset(regs_326_reset),
    .io_in(regs_326_io_in),
    .io_reset(regs_326_io_reset),
    .io_out(regs_326_io_out),
    .io_enable(regs_326_io_enable)
  );
  FringeFF regs_327 ( // @[RegFile.scala 66:20:@54308.4]
    .clock(regs_327_clock),
    .reset(regs_327_reset),
    .io_in(regs_327_io_in),
    .io_reset(regs_327_io_reset),
    .io_out(regs_327_io_out),
    .io_enable(regs_327_io_enable)
  );
  FringeFF regs_328 ( // @[RegFile.scala 66:20:@54322.4]
    .clock(regs_328_clock),
    .reset(regs_328_reset),
    .io_in(regs_328_io_in),
    .io_reset(regs_328_io_reset),
    .io_out(regs_328_io_out),
    .io_enable(regs_328_io_enable)
  );
  FringeFF regs_329 ( // @[RegFile.scala 66:20:@54336.4]
    .clock(regs_329_clock),
    .reset(regs_329_reset),
    .io_in(regs_329_io_in),
    .io_reset(regs_329_io_reset),
    .io_out(regs_329_io_out),
    .io_enable(regs_329_io_enable)
  );
  FringeFF regs_330 ( // @[RegFile.scala 66:20:@54350.4]
    .clock(regs_330_clock),
    .reset(regs_330_reset),
    .io_in(regs_330_io_in),
    .io_reset(regs_330_io_reset),
    .io_out(regs_330_io_out),
    .io_enable(regs_330_io_enable)
  );
  FringeFF regs_331 ( // @[RegFile.scala 66:20:@54364.4]
    .clock(regs_331_clock),
    .reset(regs_331_reset),
    .io_in(regs_331_io_in),
    .io_reset(regs_331_io_reset),
    .io_out(regs_331_io_out),
    .io_enable(regs_331_io_enable)
  );
  FringeFF regs_332 ( // @[RegFile.scala 66:20:@54378.4]
    .clock(regs_332_clock),
    .reset(regs_332_reset),
    .io_in(regs_332_io_in),
    .io_reset(regs_332_io_reset),
    .io_out(regs_332_io_out),
    .io_enable(regs_332_io_enable)
  );
  FringeFF regs_333 ( // @[RegFile.scala 66:20:@54392.4]
    .clock(regs_333_clock),
    .reset(regs_333_reset),
    .io_in(regs_333_io_in),
    .io_reset(regs_333_io_reset),
    .io_out(regs_333_io_out),
    .io_enable(regs_333_io_enable)
  );
  FringeFF regs_334 ( // @[RegFile.scala 66:20:@54406.4]
    .clock(regs_334_clock),
    .reset(regs_334_reset),
    .io_in(regs_334_io_in),
    .io_reset(regs_334_io_reset),
    .io_out(regs_334_io_out),
    .io_enable(regs_334_io_enable)
  );
  FringeFF regs_335 ( // @[RegFile.scala 66:20:@54420.4]
    .clock(regs_335_clock),
    .reset(regs_335_reset),
    .io_in(regs_335_io_in),
    .io_reset(regs_335_io_reset),
    .io_out(regs_335_io_out),
    .io_enable(regs_335_io_enable)
  );
  FringeFF regs_336 ( // @[RegFile.scala 66:20:@54434.4]
    .clock(regs_336_clock),
    .reset(regs_336_reset),
    .io_in(regs_336_io_in),
    .io_reset(regs_336_io_reset),
    .io_out(regs_336_io_out),
    .io_enable(regs_336_io_enable)
  );
  FringeFF regs_337 ( // @[RegFile.scala 66:20:@54448.4]
    .clock(regs_337_clock),
    .reset(regs_337_reset),
    .io_in(regs_337_io_in),
    .io_reset(regs_337_io_reset),
    .io_out(regs_337_io_out),
    .io_enable(regs_337_io_enable)
  );
  FringeFF regs_338 ( // @[RegFile.scala 66:20:@54462.4]
    .clock(regs_338_clock),
    .reset(regs_338_reset),
    .io_in(regs_338_io_in),
    .io_reset(regs_338_io_reset),
    .io_out(regs_338_io_out),
    .io_enable(regs_338_io_enable)
  );
  FringeFF regs_339 ( // @[RegFile.scala 66:20:@54476.4]
    .clock(regs_339_clock),
    .reset(regs_339_reset),
    .io_in(regs_339_io_in),
    .io_reset(regs_339_io_reset),
    .io_out(regs_339_io_out),
    .io_enable(regs_339_io_enable)
  );
  FringeFF regs_340 ( // @[RegFile.scala 66:20:@54490.4]
    .clock(regs_340_clock),
    .reset(regs_340_reset),
    .io_in(regs_340_io_in),
    .io_reset(regs_340_io_reset),
    .io_out(regs_340_io_out),
    .io_enable(regs_340_io_enable)
  );
  FringeFF regs_341 ( // @[RegFile.scala 66:20:@54504.4]
    .clock(regs_341_clock),
    .reset(regs_341_reset),
    .io_in(regs_341_io_in),
    .io_reset(regs_341_io_reset),
    .io_out(regs_341_io_out),
    .io_enable(regs_341_io_enable)
  );
  FringeFF regs_342 ( // @[RegFile.scala 66:20:@54518.4]
    .clock(regs_342_clock),
    .reset(regs_342_reset),
    .io_in(regs_342_io_in),
    .io_reset(regs_342_io_reset),
    .io_out(regs_342_io_out),
    .io_enable(regs_342_io_enable)
  );
  FringeFF regs_343 ( // @[RegFile.scala 66:20:@54532.4]
    .clock(regs_343_clock),
    .reset(regs_343_reset),
    .io_in(regs_343_io_in),
    .io_reset(regs_343_io_reset),
    .io_out(regs_343_io_out),
    .io_enable(regs_343_io_enable)
  );
  FringeFF regs_344 ( // @[RegFile.scala 66:20:@54546.4]
    .clock(regs_344_clock),
    .reset(regs_344_reset),
    .io_in(regs_344_io_in),
    .io_reset(regs_344_io_reset),
    .io_out(regs_344_io_out),
    .io_enable(regs_344_io_enable)
  );
  FringeFF regs_345 ( // @[RegFile.scala 66:20:@54560.4]
    .clock(regs_345_clock),
    .reset(regs_345_reset),
    .io_in(regs_345_io_in),
    .io_reset(regs_345_io_reset),
    .io_out(regs_345_io_out),
    .io_enable(regs_345_io_enable)
  );
  FringeFF regs_346 ( // @[RegFile.scala 66:20:@54574.4]
    .clock(regs_346_clock),
    .reset(regs_346_reset),
    .io_in(regs_346_io_in),
    .io_reset(regs_346_io_reset),
    .io_out(regs_346_io_out),
    .io_enable(regs_346_io_enable)
  );
  FringeFF regs_347 ( // @[RegFile.scala 66:20:@54588.4]
    .clock(regs_347_clock),
    .reset(regs_347_reset),
    .io_in(regs_347_io_in),
    .io_reset(regs_347_io_reset),
    .io_out(regs_347_io_out),
    .io_enable(regs_347_io_enable)
  );
  FringeFF regs_348 ( // @[RegFile.scala 66:20:@54602.4]
    .clock(regs_348_clock),
    .reset(regs_348_reset),
    .io_in(regs_348_io_in),
    .io_reset(regs_348_io_reset),
    .io_out(regs_348_io_out),
    .io_enable(regs_348_io_enable)
  );
  FringeFF regs_349 ( // @[RegFile.scala 66:20:@54616.4]
    .clock(regs_349_clock),
    .reset(regs_349_reset),
    .io_in(regs_349_io_in),
    .io_reset(regs_349_io_reset),
    .io_out(regs_349_io_out),
    .io_enable(regs_349_io_enable)
  );
  FringeFF regs_350 ( // @[RegFile.scala 66:20:@54630.4]
    .clock(regs_350_clock),
    .reset(regs_350_reset),
    .io_in(regs_350_io_in),
    .io_reset(regs_350_io_reset),
    .io_out(regs_350_io_out),
    .io_enable(regs_350_io_enable)
  );
  FringeFF regs_351 ( // @[RegFile.scala 66:20:@54644.4]
    .clock(regs_351_clock),
    .reset(regs_351_reset),
    .io_in(regs_351_io_in),
    .io_reset(regs_351_io_reset),
    .io_out(regs_351_io_out),
    .io_enable(regs_351_io_enable)
  );
  FringeFF regs_352 ( // @[RegFile.scala 66:20:@54658.4]
    .clock(regs_352_clock),
    .reset(regs_352_reset),
    .io_in(regs_352_io_in),
    .io_reset(regs_352_io_reset),
    .io_out(regs_352_io_out),
    .io_enable(regs_352_io_enable)
  );
  FringeFF regs_353 ( // @[RegFile.scala 66:20:@54672.4]
    .clock(regs_353_clock),
    .reset(regs_353_reset),
    .io_in(regs_353_io_in),
    .io_reset(regs_353_io_reset),
    .io_out(regs_353_io_out),
    .io_enable(regs_353_io_enable)
  );
  FringeFF regs_354 ( // @[RegFile.scala 66:20:@54686.4]
    .clock(regs_354_clock),
    .reset(regs_354_reset),
    .io_in(regs_354_io_in),
    .io_reset(regs_354_io_reset),
    .io_out(regs_354_io_out),
    .io_enable(regs_354_io_enable)
  );
  FringeFF regs_355 ( // @[RegFile.scala 66:20:@54700.4]
    .clock(regs_355_clock),
    .reset(regs_355_reset),
    .io_in(regs_355_io_in),
    .io_reset(regs_355_io_reset),
    .io_out(regs_355_io_out),
    .io_enable(regs_355_io_enable)
  );
  FringeFF regs_356 ( // @[RegFile.scala 66:20:@54714.4]
    .clock(regs_356_clock),
    .reset(regs_356_reset),
    .io_in(regs_356_io_in),
    .io_reset(regs_356_io_reset),
    .io_out(regs_356_io_out),
    .io_enable(regs_356_io_enable)
  );
  FringeFF regs_357 ( // @[RegFile.scala 66:20:@54728.4]
    .clock(regs_357_clock),
    .reset(regs_357_reset),
    .io_in(regs_357_io_in),
    .io_reset(regs_357_io_reset),
    .io_out(regs_357_io_out),
    .io_enable(regs_357_io_enable)
  );
  FringeFF regs_358 ( // @[RegFile.scala 66:20:@54742.4]
    .clock(regs_358_clock),
    .reset(regs_358_reset),
    .io_in(regs_358_io_in),
    .io_reset(regs_358_io_reset),
    .io_out(regs_358_io_out),
    .io_enable(regs_358_io_enable)
  );
  FringeFF regs_359 ( // @[RegFile.scala 66:20:@54756.4]
    .clock(regs_359_clock),
    .reset(regs_359_reset),
    .io_in(regs_359_io_in),
    .io_reset(regs_359_io_reset),
    .io_out(regs_359_io_out),
    .io_enable(regs_359_io_enable)
  );
  FringeFF regs_360 ( // @[RegFile.scala 66:20:@54770.4]
    .clock(regs_360_clock),
    .reset(regs_360_reset),
    .io_in(regs_360_io_in),
    .io_reset(regs_360_io_reset),
    .io_out(regs_360_io_out),
    .io_enable(regs_360_io_enable)
  );
  FringeFF regs_361 ( // @[RegFile.scala 66:20:@54784.4]
    .clock(regs_361_clock),
    .reset(regs_361_reset),
    .io_in(regs_361_io_in),
    .io_reset(regs_361_io_reset),
    .io_out(regs_361_io_out),
    .io_enable(regs_361_io_enable)
  );
  FringeFF regs_362 ( // @[RegFile.scala 66:20:@54798.4]
    .clock(regs_362_clock),
    .reset(regs_362_reset),
    .io_in(regs_362_io_in),
    .io_reset(regs_362_io_reset),
    .io_out(regs_362_io_out),
    .io_enable(regs_362_io_enable)
  );
  FringeFF regs_363 ( // @[RegFile.scala 66:20:@54812.4]
    .clock(regs_363_clock),
    .reset(regs_363_reset),
    .io_in(regs_363_io_in),
    .io_reset(regs_363_io_reset),
    .io_out(regs_363_io_out),
    .io_enable(regs_363_io_enable)
  );
  FringeFF regs_364 ( // @[RegFile.scala 66:20:@54826.4]
    .clock(regs_364_clock),
    .reset(regs_364_reset),
    .io_in(regs_364_io_in),
    .io_reset(regs_364_io_reset),
    .io_out(regs_364_io_out),
    .io_enable(regs_364_io_enable)
  );
  FringeFF regs_365 ( // @[RegFile.scala 66:20:@54840.4]
    .clock(regs_365_clock),
    .reset(regs_365_reset),
    .io_in(regs_365_io_in),
    .io_reset(regs_365_io_reset),
    .io_out(regs_365_io_out),
    .io_enable(regs_365_io_enable)
  );
  FringeFF regs_366 ( // @[RegFile.scala 66:20:@54854.4]
    .clock(regs_366_clock),
    .reset(regs_366_reset),
    .io_in(regs_366_io_in),
    .io_reset(regs_366_io_reset),
    .io_out(regs_366_io_out),
    .io_enable(regs_366_io_enable)
  );
  FringeFF regs_367 ( // @[RegFile.scala 66:20:@54868.4]
    .clock(regs_367_clock),
    .reset(regs_367_reset),
    .io_in(regs_367_io_in),
    .io_reset(regs_367_io_reset),
    .io_out(regs_367_io_out),
    .io_enable(regs_367_io_enable)
  );
  FringeFF regs_368 ( // @[RegFile.scala 66:20:@54882.4]
    .clock(regs_368_clock),
    .reset(regs_368_reset),
    .io_in(regs_368_io_in),
    .io_reset(regs_368_io_reset),
    .io_out(regs_368_io_out),
    .io_enable(regs_368_io_enable)
  );
  FringeFF regs_369 ( // @[RegFile.scala 66:20:@54896.4]
    .clock(regs_369_clock),
    .reset(regs_369_reset),
    .io_in(regs_369_io_in),
    .io_reset(regs_369_io_reset),
    .io_out(regs_369_io_out),
    .io_enable(regs_369_io_enable)
  );
  FringeFF regs_370 ( // @[RegFile.scala 66:20:@54910.4]
    .clock(regs_370_clock),
    .reset(regs_370_reset),
    .io_in(regs_370_io_in),
    .io_reset(regs_370_io_reset),
    .io_out(regs_370_io_out),
    .io_enable(regs_370_io_enable)
  );
  FringeFF regs_371 ( // @[RegFile.scala 66:20:@54924.4]
    .clock(regs_371_clock),
    .reset(regs_371_reset),
    .io_in(regs_371_io_in),
    .io_reset(regs_371_io_reset),
    .io_out(regs_371_io_out),
    .io_enable(regs_371_io_enable)
  );
  FringeFF regs_372 ( // @[RegFile.scala 66:20:@54938.4]
    .clock(regs_372_clock),
    .reset(regs_372_reset),
    .io_in(regs_372_io_in),
    .io_reset(regs_372_io_reset),
    .io_out(regs_372_io_out),
    .io_enable(regs_372_io_enable)
  );
  FringeFF regs_373 ( // @[RegFile.scala 66:20:@54952.4]
    .clock(regs_373_clock),
    .reset(regs_373_reset),
    .io_in(regs_373_io_in),
    .io_reset(regs_373_io_reset),
    .io_out(regs_373_io_out),
    .io_enable(regs_373_io_enable)
  );
  FringeFF regs_374 ( // @[RegFile.scala 66:20:@54966.4]
    .clock(regs_374_clock),
    .reset(regs_374_reset),
    .io_in(regs_374_io_in),
    .io_reset(regs_374_io_reset),
    .io_out(regs_374_io_out),
    .io_enable(regs_374_io_enable)
  );
  FringeFF regs_375 ( // @[RegFile.scala 66:20:@54980.4]
    .clock(regs_375_clock),
    .reset(regs_375_reset),
    .io_in(regs_375_io_in),
    .io_reset(regs_375_io_reset),
    .io_out(regs_375_io_out),
    .io_enable(regs_375_io_enable)
  );
  FringeFF regs_376 ( // @[RegFile.scala 66:20:@54994.4]
    .clock(regs_376_clock),
    .reset(regs_376_reset),
    .io_in(regs_376_io_in),
    .io_reset(regs_376_io_reset),
    .io_out(regs_376_io_out),
    .io_enable(regs_376_io_enable)
  );
  FringeFF regs_377 ( // @[RegFile.scala 66:20:@55008.4]
    .clock(regs_377_clock),
    .reset(regs_377_reset),
    .io_in(regs_377_io_in),
    .io_reset(regs_377_io_reset),
    .io_out(regs_377_io_out),
    .io_enable(regs_377_io_enable)
  );
  FringeFF regs_378 ( // @[RegFile.scala 66:20:@55022.4]
    .clock(regs_378_clock),
    .reset(regs_378_reset),
    .io_in(regs_378_io_in),
    .io_reset(regs_378_io_reset),
    .io_out(regs_378_io_out),
    .io_enable(regs_378_io_enable)
  );
  FringeFF regs_379 ( // @[RegFile.scala 66:20:@55036.4]
    .clock(regs_379_clock),
    .reset(regs_379_reset),
    .io_in(regs_379_io_in),
    .io_reset(regs_379_io_reset),
    .io_out(regs_379_io_out),
    .io_enable(regs_379_io_enable)
  );
  FringeFF regs_380 ( // @[RegFile.scala 66:20:@55050.4]
    .clock(regs_380_clock),
    .reset(regs_380_reset),
    .io_in(regs_380_io_in),
    .io_reset(regs_380_io_reset),
    .io_out(regs_380_io_out),
    .io_enable(regs_380_io_enable)
  );
  FringeFF regs_381 ( // @[RegFile.scala 66:20:@55064.4]
    .clock(regs_381_clock),
    .reset(regs_381_reset),
    .io_in(regs_381_io_in),
    .io_reset(regs_381_io_reset),
    .io_out(regs_381_io_out),
    .io_enable(regs_381_io_enable)
  );
  FringeFF regs_382 ( // @[RegFile.scala 66:20:@55078.4]
    .clock(regs_382_clock),
    .reset(regs_382_reset),
    .io_in(regs_382_io_in),
    .io_reset(regs_382_io_reset),
    .io_out(regs_382_io_out),
    .io_enable(regs_382_io_enable)
  );
  FringeFF regs_383 ( // @[RegFile.scala 66:20:@55092.4]
    .clock(regs_383_clock),
    .reset(regs_383_reset),
    .io_in(regs_383_io_in),
    .io_reset(regs_383_io_reset),
    .io_out(regs_383_io_out),
    .io_enable(regs_383_io_enable)
  );
  FringeFF regs_384 ( // @[RegFile.scala 66:20:@55106.4]
    .clock(regs_384_clock),
    .reset(regs_384_reset),
    .io_in(regs_384_io_in),
    .io_reset(regs_384_io_reset),
    .io_out(regs_384_io_out),
    .io_enable(regs_384_io_enable)
  );
  FringeFF regs_385 ( // @[RegFile.scala 66:20:@55120.4]
    .clock(regs_385_clock),
    .reset(regs_385_reset),
    .io_in(regs_385_io_in),
    .io_reset(regs_385_io_reset),
    .io_out(regs_385_io_out),
    .io_enable(regs_385_io_enable)
  );
  FringeFF regs_386 ( // @[RegFile.scala 66:20:@55134.4]
    .clock(regs_386_clock),
    .reset(regs_386_reset),
    .io_in(regs_386_io_in),
    .io_reset(regs_386_io_reset),
    .io_out(regs_386_io_out),
    .io_enable(regs_386_io_enable)
  );
  FringeFF regs_387 ( // @[RegFile.scala 66:20:@55148.4]
    .clock(regs_387_clock),
    .reset(regs_387_reset),
    .io_in(regs_387_io_in),
    .io_reset(regs_387_io_reset),
    .io_out(regs_387_io_out),
    .io_enable(regs_387_io_enable)
  );
  FringeFF regs_388 ( // @[RegFile.scala 66:20:@55162.4]
    .clock(regs_388_clock),
    .reset(regs_388_reset),
    .io_in(regs_388_io_in),
    .io_reset(regs_388_io_reset),
    .io_out(regs_388_io_out),
    .io_enable(regs_388_io_enable)
  );
  FringeFF regs_389 ( // @[RegFile.scala 66:20:@55176.4]
    .clock(regs_389_clock),
    .reset(regs_389_reset),
    .io_in(regs_389_io_in),
    .io_reset(regs_389_io_reset),
    .io_out(regs_389_io_out),
    .io_enable(regs_389_io_enable)
  );
  FringeFF regs_390 ( // @[RegFile.scala 66:20:@55190.4]
    .clock(regs_390_clock),
    .reset(regs_390_reset),
    .io_in(regs_390_io_in),
    .io_reset(regs_390_io_reset),
    .io_out(regs_390_io_out),
    .io_enable(regs_390_io_enable)
  );
  FringeFF regs_391 ( // @[RegFile.scala 66:20:@55204.4]
    .clock(regs_391_clock),
    .reset(regs_391_reset),
    .io_in(regs_391_io_in),
    .io_reset(regs_391_io_reset),
    .io_out(regs_391_io_out),
    .io_enable(regs_391_io_enable)
  );
  FringeFF regs_392 ( // @[RegFile.scala 66:20:@55218.4]
    .clock(regs_392_clock),
    .reset(regs_392_reset),
    .io_in(regs_392_io_in),
    .io_reset(regs_392_io_reset),
    .io_out(regs_392_io_out),
    .io_enable(regs_392_io_enable)
  );
  FringeFF regs_393 ( // @[RegFile.scala 66:20:@55232.4]
    .clock(regs_393_clock),
    .reset(regs_393_reset),
    .io_in(regs_393_io_in),
    .io_reset(regs_393_io_reset),
    .io_out(regs_393_io_out),
    .io_enable(regs_393_io_enable)
  );
  FringeFF regs_394 ( // @[RegFile.scala 66:20:@55246.4]
    .clock(regs_394_clock),
    .reset(regs_394_reset),
    .io_in(regs_394_io_in),
    .io_reset(regs_394_io_reset),
    .io_out(regs_394_io_out),
    .io_enable(regs_394_io_enable)
  );
  FringeFF regs_395 ( // @[RegFile.scala 66:20:@55260.4]
    .clock(regs_395_clock),
    .reset(regs_395_reset),
    .io_in(regs_395_io_in),
    .io_reset(regs_395_io_reset),
    .io_out(regs_395_io_out),
    .io_enable(regs_395_io_enable)
  );
  FringeFF regs_396 ( // @[RegFile.scala 66:20:@55274.4]
    .clock(regs_396_clock),
    .reset(regs_396_reset),
    .io_in(regs_396_io_in),
    .io_reset(regs_396_io_reset),
    .io_out(regs_396_io_out),
    .io_enable(regs_396_io_enable)
  );
  FringeFF regs_397 ( // @[RegFile.scala 66:20:@55288.4]
    .clock(regs_397_clock),
    .reset(regs_397_reset),
    .io_in(regs_397_io_in),
    .io_reset(regs_397_io_reset),
    .io_out(regs_397_io_out),
    .io_enable(regs_397_io_enable)
  );
  FringeFF regs_398 ( // @[RegFile.scala 66:20:@55302.4]
    .clock(regs_398_clock),
    .reset(regs_398_reset),
    .io_in(regs_398_io_in),
    .io_reset(regs_398_io_reset),
    .io_out(regs_398_io_out),
    .io_enable(regs_398_io_enable)
  );
  FringeFF regs_399 ( // @[RegFile.scala 66:20:@55316.4]
    .clock(regs_399_clock),
    .reset(regs_399_reset),
    .io_in(regs_399_io_in),
    .io_reset(regs_399_io_reset),
    .io_out(regs_399_io_out),
    .io_enable(regs_399_io_enable)
  );
  FringeFF regs_400 ( // @[RegFile.scala 66:20:@55330.4]
    .clock(regs_400_clock),
    .reset(regs_400_reset),
    .io_in(regs_400_io_in),
    .io_reset(regs_400_io_reset),
    .io_out(regs_400_io_out),
    .io_enable(regs_400_io_enable)
  );
  FringeFF regs_401 ( // @[RegFile.scala 66:20:@55344.4]
    .clock(regs_401_clock),
    .reset(regs_401_reset),
    .io_in(regs_401_io_in),
    .io_reset(regs_401_io_reset),
    .io_out(regs_401_io_out),
    .io_enable(regs_401_io_enable)
  );
  FringeFF regs_402 ( // @[RegFile.scala 66:20:@55358.4]
    .clock(regs_402_clock),
    .reset(regs_402_reset),
    .io_in(regs_402_io_in),
    .io_reset(regs_402_io_reset),
    .io_out(regs_402_io_out),
    .io_enable(regs_402_io_enable)
  );
  FringeFF regs_403 ( // @[RegFile.scala 66:20:@55372.4]
    .clock(regs_403_clock),
    .reset(regs_403_reset),
    .io_in(regs_403_io_in),
    .io_reset(regs_403_io_reset),
    .io_out(regs_403_io_out),
    .io_enable(regs_403_io_enable)
  );
  FringeFF regs_404 ( // @[RegFile.scala 66:20:@55386.4]
    .clock(regs_404_clock),
    .reset(regs_404_reset),
    .io_in(regs_404_io_in),
    .io_reset(regs_404_io_reset),
    .io_out(regs_404_io_out),
    .io_enable(regs_404_io_enable)
  );
  FringeFF regs_405 ( // @[RegFile.scala 66:20:@55400.4]
    .clock(regs_405_clock),
    .reset(regs_405_reset),
    .io_in(regs_405_io_in),
    .io_reset(regs_405_io_reset),
    .io_out(regs_405_io_out),
    .io_enable(regs_405_io_enable)
  );
  FringeFF regs_406 ( // @[RegFile.scala 66:20:@55414.4]
    .clock(regs_406_clock),
    .reset(regs_406_reset),
    .io_in(regs_406_io_in),
    .io_reset(regs_406_io_reset),
    .io_out(regs_406_io_out),
    .io_enable(regs_406_io_enable)
  );
  FringeFF regs_407 ( // @[RegFile.scala 66:20:@55428.4]
    .clock(regs_407_clock),
    .reset(regs_407_reset),
    .io_in(regs_407_io_in),
    .io_reset(regs_407_io_reset),
    .io_out(regs_407_io_out),
    .io_enable(regs_407_io_enable)
  );
  FringeFF regs_408 ( // @[RegFile.scala 66:20:@55442.4]
    .clock(regs_408_clock),
    .reset(regs_408_reset),
    .io_in(regs_408_io_in),
    .io_reset(regs_408_io_reset),
    .io_out(regs_408_io_out),
    .io_enable(regs_408_io_enable)
  );
  FringeFF regs_409 ( // @[RegFile.scala 66:20:@55456.4]
    .clock(regs_409_clock),
    .reset(regs_409_reset),
    .io_in(regs_409_io_in),
    .io_reset(regs_409_io_reset),
    .io_out(regs_409_io_out),
    .io_enable(regs_409_io_enable)
  );
  FringeFF regs_410 ( // @[RegFile.scala 66:20:@55470.4]
    .clock(regs_410_clock),
    .reset(regs_410_reset),
    .io_in(regs_410_io_in),
    .io_reset(regs_410_io_reset),
    .io_out(regs_410_io_out),
    .io_enable(regs_410_io_enable)
  );
  FringeFF regs_411 ( // @[RegFile.scala 66:20:@55484.4]
    .clock(regs_411_clock),
    .reset(regs_411_reset),
    .io_in(regs_411_io_in),
    .io_reset(regs_411_io_reset),
    .io_out(regs_411_io_out),
    .io_enable(regs_411_io_enable)
  );
  FringeFF regs_412 ( // @[RegFile.scala 66:20:@55498.4]
    .clock(regs_412_clock),
    .reset(regs_412_reset),
    .io_in(regs_412_io_in),
    .io_reset(regs_412_io_reset),
    .io_out(regs_412_io_out),
    .io_enable(regs_412_io_enable)
  );
  FringeFF regs_413 ( // @[RegFile.scala 66:20:@55512.4]
    .clock(regs_413_clock),
    .reset(regs_413_reset),
    .io_in(regs_413_io_in),
    .io_reset(regs_413_io_reset),
    .io_out(regs_413_io_out),
    .io_enable(regs_413_io_enable)
  );
  FringeFF regs_414 ( // @[RegFile.scala 66:20:@55526.4]
    .clock(regs_414_clock),
    .reset(regs_414_reset),
    .io_in(regs_414_io_in),
    .io_reset(regs_414_io_reset),
    .io_out(regs_414_io_out),
    .io_enable(regs_414_io_enable)
  );
  FringeFF regs_415 ( // @[RegFile.scala 66:20:@55540.4]
    .clock(regs_415_clock),
    .reset(regs_415_reset),
    .io_in(regs_415_io_in),
    .io_reset(regs_415_io_reset),
    .io_out(regs_415_io_out),
    .io_enable(regs_415_io_enable)
  );
  FringeFF regs_416 ( // @[RegFile.scala 66:20:@55554.4]
    .clock(regs_416_clock),
    .reset(regs_416_reset),
    .io_in(regs_416_io_in),
    .io_reset(regs_416_io_reset),
    .io_out(regs_416_io_out),
    .io_enable(regs_416_io_enable)
  );
  FringeFF regs_417 ( // @[RegFile.scala 66:20:@55568.4]
    .clock(regs_417_clock),
    .reset(regs_417_reset),
    .io_in(regs_417_io_in),
    .io_reset(regs_417_io_reset),
    .io_out(regs_417_io_out),
    .io_enable(regs_417_io_enable)
  );
  FringeFF regs_418 ( // @[RegFile.scala 66:20:@55582.4]
    .clock(regs_418_clock),
    .reset(regs_418_reset),
    .io_in(regs_418_io_in),
    .io_reset(regs_418_io_reset),
    .io_out(regs_418_io_out),
    .io_enable(regs_418_io_enable)
  );
  FringeFF regs_419 ( // @[RegFile.scala 66:20:@55596.4]
    .clock(regs_419_clock),
    .reset(regs_419_reset),
    .io_in(regs_419_io_in),
    .io_reset(regs_419_io_reset),
    .io_out(regs_419_io_out),
    .io_enable(regs_419_io_enable)
  );
  FringeFF regs_420 ( // @[RegFile.scala 66:20:@55610.4]
    .clock(regs_420_clock),
    .reset(regs_420_reset),
    .io_in(regs_420_io_in),
    .io_reset(regs_420_io_reset),
    .io_out(regs_420_io_out),
    .io_enable(regs_420_io_enable)
  );
  FringeFF regs_421 ( // @[RegFile.scala 66:20:@55624.4]
    .clock(regs_421_clock),
    .reset(regs_421_reset),
    .io_in(regs_421_io_in),
    .io_reset(regs_421_io_reset),
    .io_out(regs_421_io_out),
    .io_enable(regs_421_io_enable)
  );
  FringeFF regs_422 ( // @[RegFile.scala 66:20:@55638.4]
    .clock(regs_422_clock),
    .reset(regs_422_reset),
    .io_in(regs_422_io_in),
    .io_reset(regs_422_io_reset),
    .io_out(regs_422_io_out),
    .io_enable(regs_422_io_enable)
  );
  FringeFF regs_423 ( // @[RegFile.scala 66:20:@55652.4]
    .clock(regs_423_clock),
    .reset(regs_423_reset),
    .io_in(regs_423_io_in),
    .io_reset(regs_423_io_reset),
    .io_out(regs_423_io_out),
    .io_enable(regs_423_io_enable)
  );
  FringeFF regs_424 ( // @[RegFile.scala 66:20:@55666.4]
    .clock(regs_424_clock),
    .reset(regs_424_reset),
    .io_in(regs_424_io_in),
    .io_reset(regs_424_io_reset),
    .io_out(regs_424_io_out),
    .io_enable(regs_424_io_enable)
  );
  FringeFF regs_425 ( // @[RegFile.scala 66:20:@55680.4]
    .clock(regs_425_clock),
    .reset(regs_425_reset),
    .io_in(regs_425_io_in),
    .io_reset(regs_425_io_reset),
    .io_out(regs_425_io_out),
    .io_enable(regs_425_io_enable)
  );
  FringeFF regs_426 ( // @[RegFile.scala 66:20:@55694.4]
    .clock(regs_426_clock),
    .reset(regs_426_reset),
    .io_in(regs_426_io_in),
    .io_reset(regs_426_io_reset),
    .io_out(regs_426_io_out),
    .io_enable(regs_426_io_enable)
  );
  FringeFF regs_427 ( // @[RegFile.scala 66:20:@55708.4]
    .clock(regs_427_clock),
    .reset(regs_427_reset),
    .io_in(regs_427_io_in),
    .io_reset(regs_427_io_reset),
    .io_out(regs_427_io_out),
    .io_enable(regs_427_io_enable)
  );
  FringeFF regs_428 ( // @[RegFile.scala 66:20:@55722.4]
    .clock(regs_428_clock),
    .reset(regs_428_reset),
    .io_in(regs_428_io_in),
    .io_reset(regs_428_io_reset),
    .io_out(regs_428_io_out),
    .io_enable(regs_428_io_enable)
  );
  FringeFF regs_429 ( // @[RegFile.scala 66:20:@55736.4]
    .clock(regs_429_clock),
    .reset(regs_429_reset),
    .io_in(regs_429_io_in),
    .io_reset(regs_429_io_reset),
    .io_out(regs_429_io_out),
    .io_enable(regs_429_io_enable)
  );
  FringeFF regs_430 ( // @[RegFile.scala 66:20:@55750.4]
    .clock(regs_430_clock),
    .reset(regs_430_reset),
    .io_in(regs_430_io_in),
    .io_reset(regs_430_io_reset),
    .io_out(regs_430_io_out),
    .io_enable(regs_430_io_enable)
  );
  FringeFF regs_431 ( // @[RegFile.scala 66:20:@55764.4]
    .clock(regs_431_clock),
    .reset(regs_431_reset),
    .io_in(regs_431_io_in),
    .io_reset(regs_431_io_reset),
    .io_out(regs_431_io_out),
    .io_enable(regs_431_io_enable)
  );
  FringeFF regs_432 ( // @[RegFile.scala 66:20:@55778.4]
    .clock(regs_432_clock),
    .reset(regs_432_reset),
    .io_in(regs_432_io_in),
    .io_reset(regs_432_io_reset),
    .io_out(regs_432_io_out),
    .io_enable(regs_432_io_enable)
  );
  FringeFF regs_433 ( // @[RegFile.scala 66:20:@55792.4]
    .clock(regs_433_clock),
    .reset(regs_433_reset),
    .io_in(regs_433_io_in),
    .io_reset(regs_433_io_reset),
    .io_out(regs_433_io_out),
    .io_enable(regs_433_io_enable)
  );
  FringeFF regs_434 ( // @[RegFile.scala 66:20:@55806.4]
    .clock(regs_434_clock),
    .reset(regs_434_reset),
    .io_in(regs_434_io_in),
    .io_reset(regs_434_io_reset),
    .io_out(regs_434_io_out),
    .io_enable(regs_434_io_enable)
  );
  FringeFF regs_435 ( // @[RegFile.scala 66:20:@55820.4]
    .clock(regs_435_clock),
    .reset(regs_435_reset),
    .io_in(regs_435_io_in),
    .io_reset(regs_435_io_reset),
    .io_out(regs_435_io_out),
    .io_enable(regs_435_io_enable)
  );
  FringeFF regs_436 ( // @[RegFile.scala 66:20:@55834.4]
    .clock(regs_436_clock),
    .reset(regs_436_reset),
    .io_in(regs_436_io_in),
    .io_reset(regs_436_io_reset),
    .io_out(regs_436_io_out),
    .io_enable(regs_436_io_enable)
  );
  FringeFF regs_437 ( // @[RegFile.scala 66:20:@55848.4]
    .clock(regs_437_clock),
    .reset(regs_437_reset),
    .io_in(regs_437_io_in),
    .io_reset(regs_437_io_reset),
    .io_out(regs_437_io_out),
    .io_enable(regs_437_io_enable)
  );
  FringeFF regs_438 ( // @[RegFile.scala 66:20:@55862.4]
    .clock(regs_438_clock),
    .reset(regs_438_reset),
    .io_in(regs_438_io_in),
    .io_reset(regs_438_io_reset),
    .io_out(regs_438_io_out),
    .io_enable(regs_438_io_enable)
  );
  FringeFF regs_439 ( // @[RegFile.scala 66:20:@55876.4]
    .clock(regs_439_clock),
    .reset(regs_439_reset),
    .io_in(regs_439_io_in),
    .io_reset(regs_439_io_reset),
    .io_out(regs_439_io_out),
    .io_enable(regs_439_io_enable)
  );
  FringeFF regs_440 ( // @[RegFile.scala 66:20:@55890.4]
    .clock(regs_440_clock),
    .reset(regs_440_reset),
    .io_in(regs_440_io_in),
    .io_reset(regs_440_io_reset),
    .io_out(regs_440_io_out),
    .io_enable(regs_440_io_enable)
  );
  FringeFF regs_441 ( // @[RegFile.scala 66:20:@55904.4]
    .clock(regs_441_clock),
    .reset(regs_441_reset),
    .io_in(regs_441_io_in),
    .io_reset(regs_441_io_reset),
    .io_out(regs_441_io_out),
    .io_enable(regs_441_io_enable)
  );
  FringeFF regs_442 ( // @[RegFile.scala 66:20:@55918.4]
    .clock(regs_442_clock),
    .reset(regs_442_reset),
    .io_in(regs_442_io_in),
    .io_reset(regs_442_io_reset),
    .io_out(regs_442_io_out),
    .io_enable(regs_442_io_enable)
  );
  FringeFF regs_443 ( // @[RegFile.scala 66:20:@55932.4]
    .clock(regs_443_clock),
    .reset(regs_443_reset),
    .io_in(regs_443_io_in),
    .io_reset(regs_443_io_reset),
    .io_out(regs_443_io_out),
    .io_enable(regs_443_io_enable)
  );
  FringeFF regs_444 ( // @[RegFile.scala 66:20:@55946.4]
    .clock(regs_444_clock),
    .reset(regs_444_reset),
    .io_in(regs_444_io_in),
    .io_reset(regs_444_io_reset),
    .io_out(regs_444_io_out),
    .io_enable(regs_444_io_enable)
  );
  FringeFF regs_445 ( // @[RegFile.scala 66:20:@55960.4]
    .clock(regs_445_clock),
    .reset(regs_445_reset),
    .io_in(regs_445_io_in),
    .io_reset(regs_445_io_reset),
    .io_out(regs_445_io_out),
    .io_enable(regs_445_io_enable)
  );
  FringeFF regs_446 ( // @[RegFile.scala 66:20:@55974.4]
    .clock(regs_446_clock),
    .reset(regs_446_reset),
    .io_in(regs_446_io_in),
    .io_reset(regs_446_io_reset),
    .io_out(regs_446_io_out),
    .io_enable(regs_446_io_enable)
  );
  FringeFF regs_447 ( // @[RegFile.scala 66:20:@55988.4]
    .clock(regs_447_clock),
    .reset(regs_447_reset),
    .io_in(regs_447_io_in),
    .io_reset(regs_447_io_reset),
    .io_out(regs_447_io_out),
    .io_enable(regs_447_io_enable)
  );
  FringeFF regs_448 ( // @[RegFile.scala 66:20:@56002.4]
    .clock(regs_448_clock),
    .reset(regs_448_reset),
    .io_in(regs_448_io_in),
    .io_reset(regs_448_io_reset),
    .io_out(regs_448_io_out),
    .io_enable(regs_448_io_enable)
  );
  FringeFF regs_449 ( // @[RegFile.scala 66:20:@56016.4]
    .clock(regs_449_clock),
    .reset(regs_449_reset),
    .io_in(regs_449_io_in),
    .io_reset(regs_449_io_reset),
    .io_out(regs_449_io_out),
    .io_enable(regs_449_io_enable)
  );
  FringeFF regs_450 ( // @[RegFile.scala 66:20:@56030.4]
    .clock(regs_450_clock),
    .reset(regs_450_reset),
    .io_in(regs_450_io_in),
    .io_reset(regs_450_io_reset),
    .io_out(regs_450_io_out),
    .io_enable(regs_450_io_enable)
  );
  FringeFF regs_451 ( // @[RegFile.scala 66:20:@56044.4]
    .clock(regs_451_clock),
    .reset(regs_451_reset),
    .io_in(regs_451_io_in),
    .io_reset(regs_451_io_reset),
    .io_out(regs_451_io_out),
    .io_enable(regs_451_io_enable)
  );
  FringeFF regs_452 ( // @[RegFile.scala 66:20:@56058.4]
    .clock(regs_452_clock),
    .reset(regs_452_reset),
    .io_in(regs_452_io_in),
    .io_reset(regs_452_io_reset),
    .io_out(regs_452_io_out),
    .io_enable(regs_452_io_enable)
  );
  FringeFF regs_453 ( // @[RegFile.scala 66:20:@56072.4]
    .clock(regs_453_clock),
    .reset(regs_453_reset),
    .io_in(regs_453_io_in),
    .io_reset(regs_453_io_reset),
    .io_out(regs_453_io_out),
    .io_enable(regs_453_io_enable)
  );
  FringeFF regs_454 ( // @[RegFile.scala 66:20:@56086.4]
    .clock(regs_454_clock),
    .reset(regs_454_reset),
    .io_in(regs_454_io_in),
    .io_reset(regs_454_io_reset),
    .io_out(regs_454_io_out),
    .io_enable(regs_454_io_enable)
  );
  FringeFF regs_455 ( // @[RegFile.scala 66:20:@56100.4]
    .clock(regs_455_clock),
    .reset(regs_455_reset),
    .io_in(regs_455_io_in),
    .io_reset(regs_455_io_reset),
    .io_out(regs_455_io_out),
    .io_enable(regs_455_io_enable)
  );
  FringeFF regs_456 ( // @[RegFile.scala 66:20:@56114.4]
    .clock(regs_456_clock),
    .reset(regs_456_reset),
    .io_in(regs_456_io_in),
    .io_reset(regs_456_io_reset),
    .io_out(regs_456_io_out),
    .io_enable(regs_456_io_enable)
  );
  FringeFF regs_457 ( // @[RegFile.scala 66:20:@56128.4]
    .clock(regs_457_clock),
    .reset(regs_457_reset),
    .io_in(regs_457_io_in),
    .io_reset(regs_457_io_reset),
    .io_out(regs_457_io_out),
    .io_enable(regs_457_io_enable)
  );
  FringeFF regs_458 ( // @[RegFile.scala 66:20:@56142.4]
    .clock(regs_458_clock),
    .reset(regs_458_reset),
    .io_in(regs_458_io_in),
    .io_reset(regs_458_io_reset),
    .io_out(regs_458_io_out),
    .io_enable(regs_458_io_enable)
  );
  FringeFF regs_459 ( // @[RegFile.scala 66:20:@56156.4]
    .clock(regs_459_clock),
    .reset(regs_459_reset),
    .io_in(regs_459_io_in),
    .io_reset(regs_459_io_reset),
    .io_out(regs_459_io_out),
    .io_enable(regs_459_io_enable)
  );
  FringeFF regs_460 ( // @[RegFile.scala 66:20:@56170.4]
    .clock(regs_460_clock),
    .reset(regs_460_reset),
    .io_in(regs_460_io_in),
    .io_reset(regs_460_io_reset),
    .io_out(regs_460_io_out),
    .io_enable(regs_460_io_enable)
  );
  FringeFF regs_461 ( // @[RegFile.scala 66:20:@56184.4]
    .clock(regs_461_clock),
    .reset(regs_461_reset),
    .io_in(regs_461_io_in),
    .io_reset(regs_461_io_reset),
    .io_out(regs_461_io_out),
    .io_enable(regs_461_io_enable)
  );
  FringeFF regs_462 ( // @[RegFile.scala 66:20:@56198.4]
    .clock(regs_462_clock),
    .reset(regs_462_reset),
    .io_in(regs_462_io_in),
    .io_reset(regs_462_io_reset),
    .io_out(regs_462_io_out),
    .io_enable(regs_462_io_enable)
  );
  FringeFF regs_463 ( // @[RegFile.scala 66:20:@56212.4]
    .clock(regs_463_clock),
    .reset(regs_463_reset),
    .io_in(regs_463_io_in),
    .io_reset(regs_463_io_reset),
    .io_out(regs_463_io_out),
    .io_enable(regs_463_io_enable)
  );
  FringeFF regs_464 ( // @[RegFile.scala 66:20:@56226.4]
    .clock(regs_464_clock),
    .reset(regs_464_reset),
    .io_in(regs_464_io_in),
    .io_reset(regs_464_io_reset),
    .io_out(regs_464_io_out),
    .io_enable(regs_464_io_enable)
  );
  FringeFF regs_465 ( // @[RegFile.scala 66:20:@56240.4]
    .clock(regs_465_clock),
    .reset(regs_465_reset),
    .io_in(regs_465_io_in),
    .io_reset(regs_465_io_reset),
    .io_out(regs_465_io_out),
    .io_enable(regs_465_io_enable)
  );
  FringeFF regs_466 ( // @[RegFile.scala 66:20:@56254.4]
    .clock(regs_466_clock),
    .reset(regs_466_reset),
    .io_in(regs_466_io_in),
    .io_reset(regs_466_io_reset),
    .io_out(regs_466_io_out),
    .io_enable(regs_466_io_enable)
  );
  FringeFF regs_467 ( // @[RegFile.scala 66:20:@56268.4]
    .clock(regs_467_clock),
    .reset(regs_467_reset),
    .io_in(regs_467_io_in),
    .io_reset(regs_467_io_reset),
    .io_out(regs_467_io_out),
    .io_enable(regs_467_io_enable)
  );
  FringeFF regs_468 ( // @[RegFile.scala 66:20:@56282.4]
    .clock(regs_468_clock),
    .reset(regs_468_reset),
    .io_in(regs_468_io_in),
    .io_reset(regs_468_io_reset),
    .io_out(regs_468_io_out),
    .io_enable(regs_468_io_enable)
  );
  FringeFF regs_469 ( // @[RegFile.scala 66:20:@56296.4]
    .clock(regs_469_clock),
    .reset(regs_469_reset),
    .io_in(regs_469_io_in),
    .io_reset(regs_469_io_reset),
    .io_out(regs_469_io_out),
    .io_enable(regs_469_io_enable)
  );
  FringeFF regs_470 ( // @[RegFile.scala 66:20:@56310.4]
    .clock(regs_470_clock),
    .reset(regs_470_reset),
    .io_in(regs_470_io_in),
    .io_reset(regs_470_io_reset),
    .io_out(regs_470_io_out),
    .io_enable(regs_470_io_enable)
  );
  FringeFF regs_471 ( // @[RegFile.scala 66:20:@56324.4]
    .clock(regs_471_clock),
    .reset(regs_471_reset),
    .io_in(regs_471_io_in),
    .io_reset(regs_471_io_reset),
    .io_out(regs_471_io_out),
    .io_enable(regs_471_io_enable)
  );
  FringeFF regs_472 ( // @[RegFile.scala 66:20:@56338.4]
    .clock(regs_472_clock),
    .reset(regs_472_reset),
    .io_in(regs_472_io_in),
    .io_reset(regs_472_io_reset),
    .io_out(regs_472_io_out),
    .io_enable(regs_472_io_enable)
  );
  FringeFF regs_473 ( // @[RegFile.scala 66:20:@56352.4]
    .clock(regs_473_clock),
    .reset(regs_473_reset),
    .io_in(regs_473_io_in),
    .io_reset(regs_473_io_reset),
    .io_out(regs_473_io_out),
    .io_enable(regs_473_io_enable)
  );
  FringeFF regs_474 ( // @[RegFile.scala 66:20:@56366.4]
    .clock(regs_474_clock),
    .reset(regs_474_reset),
    .io_in(regs_474_io_in),
    .io_reset(regs_474_io_reset),
    .io_out(regs_474_io_out),
    .io_enable(regs_474_io_enable)
  );
  FringeFF regs_475 ( // @[RegFile.scala 66:20:@56380.4]
    .clock(regs_475_clock),
    .reset(regs_475_reset),
    .io_in(regs_475_io_in),
    .io_reset(regs_475_io_reset),
    .io_out(regs_475_io_out),
    .io_enable(regs_475_io_enable)
  );
  FringeFF regs_476 ( // @[RegFile.scala 66:20:@56394.4]
    .clock(regs_476_clock),
    .reset(regs_476_reset),
    .io_in(regs_476_io_in),
    .io_reset(regs_476_io_reset),
    .io_out(regs_476_io_out),
    .io_enable(regs_476_io_enable)
  );
  FringeFF regs_477 ( // @[RegFile.scala 66:20:@56408.4]
    .clock(regs_477_clock),
    .reset(regs_477_reset),
    .io_in(regs_477_io_in),
    .io_reset(regs_477_io_reset),
    .io_out(regs_477_io_out),
    .io_enable(regs_477_io_enable)
  );
  FringeFF regs_478 ( // @[RegFile.scala 66:20:@56422.4]
    .clock(regs_478_clock),
    .reset(regs_478_reset),
    .io_in(regs_478_io_in),
    .io_reset(regs_478_io_reset),
    .io_out(regs_478_io_out),
    .io_enable(regs_478_io_enable)
  );
  FringeFF regs_479 ( // @[RegFile.scala 66:20:@56436.4]
    .clock(regs_479_clock),
    .reset(regs_479_reset),
    .io_in(regs_479_io_in),
    .io_reset(regs_479_io_reset),
    .io_out(regs_479_io_out),
    .io_enable(regs_479_io_enable)
  );
  FringeFF regs_480 ( // @[RegFile.scala 66:20:@56450.4]
    .clock(regs_480_clock),
    .reset(regs_480_reset),
    .io_in(regs_480_io_in),
    .io_reset(regs_480_io_reset),
    .io_out(regs_480_io_out),
    .io_enable(regs_480_io_enable)
  );
  FringeFF regs_481 ( // @[RegFile.scala 66:20:@56464.4]
    .clock(regs_481_clock),
    .reset(regs_481_reset),
    .io_in(regs_481_io_in),
    .io_reset(regs_481_io_reset),
    .io_out(regs_481_io_out),
    .io_enable(regs_481_io_enable)
  );
  FringeFF regs_482 ( // @[RegFile.scala 66:20:@56478.4]
    .clock(regs_482_clock),
    .reset(regs_482_reset),
    .io_in(regs_482_io_in),
    .io_reset(regs_482_io_reset),
    .io_out(regs_482_io_out),
    .io_enable(regs_482_io_enable)
  );
  FringeFF regs_483 ( // @[RegFile.scala 66:20:@56492.4]
    .clock(regs_483_clock),
    .reset(regs_483_reset),
    .io_in(regs_483_io_in),
    .io_reset(regs_483_io_reset),
    .io_out(regs_483_io_out),
    .io_enable(regs_483_io_enable)
  );
  FringeFF regs_484 ( // @[RegFile.scala 66:20:@56506.4]
    .clock(regs_484_clock),
    .reset(regs_484_reset),
    .io_in(regs_484_io_in),
    .io_reset(regs_484_io_reset),
    .io_out(regs_484_io_out),
    .io_enable(regs_484_io_enable)
  );
  FringeFF regs_485 ( // @[RegFile.scala 66:20:@56520.4]
    .clock(regs_485_clock),
    .reset(regs_485_reset),
    .io_in(regs_485_io_in),
    .io_reset(regs_485_io_reset),
    .io_out(regs_485_io_out),
    .io_enable(regs_485_io_enable)
  );
  FringeFF regs_486 ( // @[RegFile.scala 66:20:@56534.4]
    .clock(regs_486_clock),
    .reset(regs_486_reset),
    .io_in(regs_486_io_in),
    .io_reset(regs_486_io_reset),
    .io_out(regs_486_io_out),
    .io_enable(regs_486_io_enable)
  );
  FringeFF regs_487 ( // @[RegFile.scala 66:20:@56548.4]
    .clock(regs_487_clock),
    .reset(regs_487_reset),
    .io_in(regs_487_io_in),
    .io_reset(regs_487_io_reset),
    .io_out(regs_487_io_out),
    .io_enable(regs_487_io_enable)
  );
  FringeFF regs_488 ( // @[RegFile.scala 66:20:@56562.4]
    .clock(regs_488_clock),
    .reset(regs_488_reset),
    .io_in(regs_488_io_in),
    .io_reset(regs_488_io_reset),
    .io_out(regs_488_io_out),
    .io_enable(regs_488_io_enable)
  );
  FringeFF regs_489 ( // @[RegFile.scala 66:20:@56576.4]
    .clock(regs_489_clock),
    .reset(regs_489_reset),
    .io_in(regs_489_io_in),
    .io_reset(regs_489_io_reset),
    .io_out(regs_489_io_out),
    .io_enable(regs_489_io_enable)
  );
  FringeFF regs_490 ( // @[RegFile.scala 66:20:@56590.4]
    .clock(regs_490_clock),
    .reset(regs_490_reset),
    .io_in(regs_490_io_in),
    .io_reset(regs_490_io_reset),
    .io_out(regs_490_io_out),
    .io_enable(regs_490_io_enable)
  );
  FringeFF regs_491 ( // @[RegFile.scala 66:20:@56604.4]
    .clock(regs_491_clock),
    .reset(regs_491_reset),
    .io_in(regs_491_io_in),
    .io_reset(regs_491_io_reset),
    .io_out(regs_491_io_out),
    .io_enable(regs_491_io_enable)
  );
  FringeFF regs_492 ( // @[RegFile.scala 66:20:@56618.4]
    .clock(regs_492_clock),
    .reset(regs_492_reset),
    .io_in(regs_492_io_in),
    .io_reset(regs_492_io_reset),
    .io_out(regs_492_io_out),
    .io_enable(regs_492_io_enable)
  );
  FringeFF regs_493 ( // @[RegFile.scala 66:20:@56632.4]
    .clock(regs_493_clock),
    .reset(regs_493_reset),
    .io_in(regs_493_io_in),
    .io_reset(regs_493_io_reset),
    .io_out(regs_493_io_out),
    .io_enable(regs_493_io_enable)
  );
  FringeFF regs_494 ( // @[RegFile.scala 66:20:@56646.4]
    .clock(regs_494_clock),
    .reset(regs_494_reset),
    .io_in(regs_494_io_in),
    .io_reset(regs_494_io_reset),
    .io_out(regs_494_io_out),
    .io_enable(regs_494_io_enable)
  );
  FringeFF regs_495 ( // @[RegFile.scala 66:20:@56660.4]
    .clock(regs_495_clock),
    .reset(regs_495_reset),
    .io_in(regs_495_io_in),
    .io_reset(regs_495_io_reset),
    .io_out(regs_495_io_out),
    .io_enable(regs_495_io_enable)
  );
  FringeFF regs_496 ( // @[RegFile.scala 66:20:@56674.4]
    .clock(regs_496_clock),
    .reset(regs_496_reset),
    .io_in(regs_496_io_in),
    .io_reset(regs_496_io_reset),
    .io_out(regs_496_io_out),
    .io_enable(regs_496_io_enable)
  );
  FringeFF regs_497 ( // @[RegFile.scala 66:20:@56688.4]
    .clock(regs_497_clock),
    .reset(regs_497_reset),
    .io_in(regs_497_io_in),
    .io_reset(regs_497_io_reset),
    .io_out(regs_497_io_out),
    .io_enable(regs_497_io_enable)
  );
  FringeFF regs_498 ( // @[RegFile.scala 66:20:@56702.4]
    .clock(regs_498_clock),
    .reset(regs_498_reset),
    .io_in(regs_498_io_in),
    .io_reset(regs_498_io_reset),
    .io_out(regs_498_io_out),
    .io_enable(regs_498_io_enable)
  );
  FringeFF regs_499 ( // @[RegFile.scala 66:20:@56716.4]
    .clock(regs_499_clock),
    .reset(regs_499_reset),
    .io_in(regs_499_io_in),
    .io_reset(regs_499_io_reset),
    .io_out(regs_499_io_out),
    .io_enable(regs_499_io_enable)
  );
  FringeFF regs_500 ( // @[RegFile.scala 66:20:@56730.4]
    .clock(regs_500_clock),
    .reset(regs_500_reset),
    .io_in(regs_500_io_in),
    .io_reset(regs_500_io_reset),
    .io_out(regs_500_io_out),
    .io_enable(regs_500_io_enable)
  );
  FringeFF regs_501 ( // @[RegFile.scala 66:20:@56744.4]
    .clock(regs_501_clock),
    .reset(regs_501_reset),
    .io_in(regs_501_io_in),
    .io_reset(regs_501_io_reset),
    .io_out(regs_501_io_out),
    .io_enable(regs_501_io_enable)
  );
  FringeFF regs_502 ( // @[RegFile.scala 66:20:@56758.4]
    .clock(regs_502_clock),
    .reset(regs_502_reset),
    .io_in(regs_502_io_in),
    .io_reset(regs_502_io_reset),
    .io_out(regs_502_io_out),
    .io_enable(regs_502_io_enable)
  );
  FringeFF regs_503 ( // @[RegFile.scala 66:20:@56772.4]
    .clock(regs_503_clock),
    .reset(regs_503_reset),
    .io_in(regs_503_io_in),
    .io_reset(regs_503_io_reset),
    .io_out(regs_503_io_out),
    .io_enable(regs_503_io_enable)
  );
  FringeFF regs_504 ( // @[RegFile.scala 66:20:@56786.4]
    .clock(regs_504_clock),
    .reset(regs_504_reset),
    .io_in(regs_504_io_in),
    .io_reset(regs_504_io_reset),
    .io_out(regs_504_io_out),
    .io_enable(regs_504_io_enable)
  );
  FringeFF regs_505 ( // @[RegFile.scala 66:20:@56800.4]
    .clock(regs_505_clock),
    .reset(regs_505_reset),
    .io_in(regs_505_io_in),
    .io_reset(regs_505_io_reset),
    .io_out(regs_505_io_out),
    .io_enable(regs_505_io_enable)
  );
  FringeFF regs_506 ( // @[RegFile.scala 66:20:@56814.4]
    .clock(regs_506_clock),
    .reset(regs_506_reset),
    .io_in(regs_506_io_in),
    .io_reset(regs_506_io_reset),
    .io_out(regs_506_io_out),
    .io_enable(regs_506_io_enable)
  );
  FringeFF regs_507 ( // @[RegFile.scala 66:20:@56828.4]
    .clock(regs_507_clock),
    .reset(regs_507_reset),
    .io_in(regs_507_io_in),
    .io_reset(regs_507_io_reset),
    .io_out(regs_507_io_out),
    .io_enable(regs_507_io_enable)
  );
  FringeFF regs_508 ( // @[RegFile.scala 66:20:@56842.4]
    .clock(regs_508_clock),
    .reset(regs_508_reset),
    .io_in(regs_508_io_in),
    .io_reset(regs_508_io_reset),
    .io_out(regs_508_io_out),
    .io_enable(regs_508_io_enable)
  );
  FringeFF regs_509 ( // @[RegFile.scala 66:20:@56856.4]
    .clock(regs_509_clock),
    .reset(regs_509_reset),
    .io_in(regs_509_io_in),
    .io_reset(regs_509_io_reset),
    .io_out(regs_509_io_out),
    .io_enable(regs_509_io_enable)
  );
  FringeFF regs_510 ( // @[RegFile.scala 66:20:@56870.4]
    .clock(regs_510_clock),
    .reset(regs_510_reset),
    .io_in(regs_510_io_in),
    .io_reset(regs_510_io_reset),
    .io_out(regs_510_io_out),
    .io_enable(regs_510_io_enable)
  );
  FringeFF regs_511 ( // @[RegFile.scala 66:20:@56884.4]
    .clock(regs_511_clock),
    .reset(regs_511_reset),
    .io_in(regs_511_io_in),
    .io_reset(regs_511_io_reset),
    .io_out(regs_511_io_out),
    .io_enable(regs_511_io_enable)
  );
  FringeFF regs_512 ( // @[RegFile.scala 66:20:@56898.4]
    .clock(regs_512_clock),
    .reset(regs_512_reset),
    .io_in(regs_512_io_in),
    .io_reset(regs_512_io_reset),
    .io_out(regs_512_io_out),
    .io_enable(regs_512_io_enable)
  );
  FringeFF regs_513 ( // @[RegFile.scala 66:20:@56912.4]
    .clock(regs_513_clock),
    .reset(regs_513_reset),
    .io_in(regs_513_io_in),
    .io_reset(regs_513_io_reset),
    .io_out(regs_513_io_out),
    .io_enable(regs_513_io_enable)
  );
  FringeFF regs_514 ( // @[RegFile.scala 66:20:@56926.4]
    .clock(regs_514_clock),
    .reset(regs_514_reset),
    .io_in(regs_514_io_in),
    .io_reset(regs_514_io_reset),
    .io_out(regs_514_io_out),
    .io_enable(regs_514_io_enable)
  );
  FringeFF regs_515 ( // @[RegFile.scala 66:20:@56940.4]
    .clock(regs_515_clock),
    .reset(regs_515_reset),
    .io_in(regs_515_io_in),
    .io_reset(regs_515_io_reset),
    .io_out(regs_515_io_out),
    .io_enable(regs_515_io_enable)
  );
  FringeFF regs_516 ( // @[RegFile.scala 66:20:@56954.4]
    .clock(regs_516_clock),
    .reset(regs_516_reset),
    .io_in(regs_516_io_in),
    .io_reset(regs_516_io_reset),
    .io_out(regs_516_io_out),
    .io_enable(regs_516_io_enable)
  );
  FringeFF regs_517 ( // @[RegFile.scala 66:20:@56968.4]
    .clock(regs_517_clock),
    .reset(regs_517_reset),
    .io_in(regs_517_io_in),
    .io_reset(regs_517_io_reset),
    .io_out(regs_517_io_out),
    .io_enable(regs_517_io_enable)
  );
  MuxN rport ( // @[RegFile.scala 95:21:@56982.4]
    .io_ins_0(rport_io_ins_0),
    .io_ins_1(rport_io_ins_1),
    .io_ins_2(rport_io_ins_2),
    .io_ins_3(rport_io_ins_3),
    .io_ins_4(rport_io_ins_4),
    .io_ins_5(rport_io_ins_5),
    .io_ins_6(rport_io_ins_6),
    .io_ins_7(rport_io_ins_7),
    .io_ins_8(rport_io_ins_8),
    .io_ins_9(rport_io_ins_9),
    .io_ins_10(rport_io_ins_10),
    .io_ins_11(rport_io_ins_11),
    .io_ins_12(rport_io_ins_12),
    .io_ins_13(rport_io_ins_13),
    .io_ins_14(rport_io_ins_14),
    .io_ins_15(rport_io_ins_15),
    .io_ins_16(rport_io_ins_16),
    .io_ins_17(rport_io_ins_17),
    .io_ins_18(rport_io_ins_18),
    .io_ins_19(rport_io_ins_19),
    .io_ins_20(rport_io_ins_20),
    .io_ins_21(rport_io_ins_21),
    .io_ins_22(rport_io_ins_22),
    .io_ins_23(rport_io_ins_23),
    .io_ins_24(rport_io_ins_24),
    .io_ins_25(rport_io_ins_25),
    .io_ins_26(rport_io_ins_26),
    .io_ins_27(rport_io_ins_27),
    .io_ins_28(rport_io_ins_28),
    .io_ins_29(rport_io_ins_29),
    .io_ins_30(rport_io_ins_30),
    .io_ins_31(rport_io_ins_31),
    .io_ins_32(rport_io_ins_32),
    .io_ins_33(rport_io_ins_33),
    .io_ins_34(rport_io_ins_34),
    .io_ins_35(rport_io_ins_35),
    .io_ins_36(rport_io_ins_36),
    .io_ins_37(rport_io_ins_37),
    .io_ins_38(rport_io_ins_38),
    .io_ins_39(rport_io_ins_39),
    .io_ins_40(rport_io_ins_40),
    .io_ins_41(rport_io_ins_41),
    .io_ins_42(rport_io_ins_42),
    .io_ins_43(rport_io_ins_43),
    .io_ins_44(rport_io_ins_44),
    .io_ins_45(rport_io_ins_45),
    .io_ins_46(rport_io_ins_46),
    .io_ins_47(rport_io_ins_47),
    .io_ins_48(rport_io_ins_48),
    .io_ins_49(rport_io_ins_49),
    .io_ins_50(rport_io_ins_50),
    .io_ins_51(rport_io_ins_51),
    .io_ins_52(rport_io_ins_52),
    .io_ins_53(rport_io_ins_53),
    .io_ins_54(rport_io_ins_54),
    .io_ins_55(rport_io_ins_55),
    .io_ins_56(rport_io_ins_56),
    .io_ins_57(rport_io_ins_57),
    .io_ins_58(rport_io_ins_58),
    .io_ins_59(rport_io_ins_59),
    .io_ins_60(rport_io_ins_60),
    .io_ins_61(rport_io_ins_61),
    .io_ins_62(rport_io_ins_62),
    .io_ins_63(rport_io_ins_63),
    .io_ins_64(rport_io_ins_64),
    .io_ins_65(rport_io_ins_65),
    .io_ins_66(rport_io_ins_66),
    .io_ins_67(rport_io_ins_67),
    .io_ins_68(rport_io_ins_68),
    .io_ins_69(rport_io_ins_69),
    .io_ins_70(rport_io_ins_70),
    .io_ins_71(rport_io_ins_71),
    .io_ins_72(rport_io_ins_72),
    .io_ins_73(rport_io_ins_73),
    .io_ins_74(rport_io_ins_74),
    .io_ins_75(rport_io_ins_75),
    .io_ins_76(rport_io_ins_76),
    .io_ins_77(rport_io_ins_77),
    .io_ins_78(rport_io_ins_78),
    .io_ins_79(rport_io_ins_79),
    .io_ins_80(rport_io_ins_80),
    .io_ins_81(rport_io_ins_81),
    .io_ins_82(rport_io_ins_82),
    .io_ins_83(rport_io_ins_83),
    .io_ins_84(rport_io_ins_84),
    .io_ins_85(rport_io_ins_85),
    .io_ins_86(rport_io_ins_86),
    .io_ins_87(rport_io_ins_87),
    .io_ins_88(rport_io_ins_88),
    .io_ins_89(rport_io_ins_89),
    .io_ins_90(rport_io_ins_90),
    .io_ins_91(rport_io_ins_91),
    .io_ins_92(rport_io_ins_92),
    .io_ins_93(rport_io_ins_93),
    .io_ins_94(rport_io_ins_94),
    .io_ins_95(rport_io_ins_95),
    .io_ins_96(rport_io_ins_96),
    .io_ins_97(rport_io_ins_97),
    .io_ins_98(rport_io_ins_98),
    .io_ins_99(rport_io_ins_99),
    .io_ins_100(rport_io_ins_100),
    .io_ins_101(rport_io_ins_101),
    .io_ins_102(rport_io_ins_102),
    .io_ins_103(rport_io_ins_103),
    .io_ins_104(rport_io_ins_104),
    .io_ins_105(rport_io_ins_105),
    .io_ins_106(rport_io_ins_106),
    .io_ins_107(rport_io_ins_107),
    .io_ins_108(rport_io_ins_108),
    .io_ins_109(rport_io_ins_109),
    .io_ins_110(rport_io_ins_110),
    .io_ins_111(rport_io_ins_111),
    .io_ins_112(rport_io_ins_112),
    .io_ins_113(rport_io_ins_113),
    .io_ins_114(rport_io_ins_114),
    .io_ins_115(rport_io_ins_115),
    .io_ins_116(rport_io_ins_116),
    .io_ins_117(rport_io_ins_117),
    .io_ins_118(rport_io_ins_118),
    .io_ins_119(rport_io_ins_119),
    .io_ins_120(rport_io_ins_120),
    .io_ins_121(rport_io_ins_121),
    .io_ins_122(rport_io_ins_122),
    .io_ins_123(rport_io_ins_123),
    .io_ins_124(rport_io_ins_124),
    .io_ins_125(rport_io_ins_125),
    .io_ins_126(rport_io_ins_126),
    .io_ins_127(rport_io_ins_127),
    .io_ins_128(rport_io_ins_128),
    .io_ins_129(rport_io_ins_129),
    .io_ins_130(rport_io_ins_130),
    .io_ins_131(rport_io_ins_131),
    .io_ins_132(rport_io_ins_132),
    .io_ins_133(rport_io_ins_133),
    .io_ins_134(rport_io_ins_134),
    .io_ins_135(rport_io_ins_135),
    .io_ins_136(rport_io_ins_136),
    .io_ins_137(rport_io_ins_137),
    .io_ins_138(rport_io_ins_138),
    .io_ins_139(rport_io_ins_139),
    .io_ins_140(rport_io_ins_140),
    .io_ins_141(rport_io_ins_141),
    .io_ins_142(rport_io_ins_142),
    .io_ins_143(rport_io_ins_143),
    .io_ins_144(rport_io_ins_144),
    .io_ins_145(rport_io_ins_145),
    .io_ins_146(rport_io_ins_146),
    .io_ins_147(rport_io_ins_147),
    .io_ins_148(rport_io_ins_148),
    .io_ins_149(rport_io_ins_149),
    .io_ins_150(rport_io_ins_150),
    .io_ins_151(rport_io_ins_151),
    .io_ins_152(rport_io_ins_152),
    .io_ins_153(rport_io_ins_153),
    .io_ins_154(rport_io_ins_154),
    .io_ins_155(rport_io_ins_155),
    .io_ins_156(rport_io_ins_156),
    .io_ins_157(rport_io_ins_157),
    .io_ins_158(rport_io_ins_158),
    .io_ins_159(rport_io_ins_159),
    .io_ins_160(rport_io_ins_160),
    .io_ins_161(rport_io_ins_161),
    .io_ins_162(rport_io_ins_162),
    .io_ins_163(rport_io_ins_163),
    .io_ins_164(rport_io_ins_164),
    .io_ins_165(rport_io_ins_165),
    .io_ins_166(rport_io_ins_166),
    .io_ins_167(rport_io_ins_167),
    .io_ins_168(rport_io_ins_168),
    .io_ins_169(rport_io_ins_169),
    .io_ins_170(rport_io_ins_170),
    .io_ins_171(rport_io_ins_171),
    .io_ins_172(rport_io_ins_172),
    .io_ins_173(rport_io_ins_173),
    .io_ins_174(rport_io_ins_174),
    .io_ins_175(rport_io_ins_175),
    .io_ins_176(rport_io_ins_176),
    .io_ins_177(rport_io_ins_177),
    .io_ins_178(rport_io_ins_178),
    .io_ins_179(rport_io_ins_179),
    .io_ins_180(rport_io_ins_180),
    .io_ins_181(rport_io_ins_181),
    .io_ins_182(rport_io_ins_182),
    .io_ins_183(rport_io_ins_183),
    .io_ins_184(rport_io_ins_184),
    .io_ins_185(rport_io_ins_185),
    .io_ins_186(rport_io_ins_186),
    .io_ins_187(rport_io_ins_187),
    .io_ins_188(rport_io_ins_188),
    .io_ins_189(rport_io_ins_189),
    .io_ins_190(rport_io_ins_190),
    .io_ins_191(rport_io_ins_191),
    .io_ins_192(rport_io_ins_192),
    .io_ins_193(rport_io_ins_193),
    .io_ins_194(rport_io_ins_194),
    .io_ins_195(rport_io_ins_195),
    .io_ins_196(rport_io_ins_196),
    .io_ins_197(rport_io_ins_197),
    .io_ins_198(rport_io_ins_198),
    .io_ins_199(rport_io_ins_199),
    .io_ins_200(rport_io_ins_200),
    .io_ins_201(rport_io_ins_201),
    .io_ins_202(rport_io_ins_202),
    .io_ins_203(rport_io_ins_203),
    .io_ins_204(rport_io_ins_204),
    .io_ins_205(rport_io_ins_205),
    .io_ins_206(rport_io_ins_206),
    .io_ins_207(rport_io_ins_207),
    .io_ins_208(rport_io_ins_208),
    .io_ins_209(rport_io_ins_209),
    .io_ins_210(rport_io_ins_210),
    .io_ins_211(rport_io_ins_211),
    .io_ins_212(rport_io_ins_212),
    .io_ins_213(rport_io_ins_213),
    .io_ins_214(rport_io_ins_214),
    .io_ins_215(rport_io_ins_215),
    .io_ins_216(rport_io_ins_216),
    .io_ins_217(rport_io_ins_217),
    .io_ins_218(rport_io_ins_218),
    .io_ins_219(rport_io_ins_219),
    .io_ins_220(rport_io_ins_220),
    .io_ins_221(rport_io_ins_221),
    .io_ins_222(rport_io_ins_222),
    .io_ins_223(rport_io_ins_223),
    .io_ins_224(rport_io_ins_224),
    .io_ins_225(rport_io_ins_225),
    .io_ins_226(rport_io_ins_226),
    .io_ins_227(rport_io_ins_227),
    .io_ins_228(rport_io_ins_228),
    .io_ins_229(rport_io_ins_229),
    .io_ins_230(rport_io_ins_230),
    .io_ins_231(rport_io_ins_231),
    .io_ins_232(rport_io_ins_232),
    .io_ins_233(rport_io_ins_233),
    .io_ins_234(rport_io_ins_234),
    .io_ins_235(rport_io_ins_235),
    .io_ins_236(rport_io_ins_236),
    .io_ins_237(rport_io_ins_237),
    .io_ins_238(rport_io_ins_238),
    .io_ins_239(rport_io_ins_239),
    .io_ins_240(rport_io_ins_240),
    .io_ins_241(rport_io_ins_241),
    .io_ins_242(rport_io_ins_242),
    .io_ins_243(rport_io_ins_243),
    .io_ins_244(rport_io_ins_244),
    .io_ins_245(rport_io_ins_245),
    .io_ins_246(rport_io_ins_246),
    .io_ins_247(rport_io_ins_247),
    .io_ins_248(rport_io_ins_248),
    .io_ins_249(rport_io_ins_249),
    .io_ins_250(rport_io_ins_250),
    .io_ins_251(rport_io_ins_251),
    .io_ins_252(rport_io_ins_252),
    .io_ins_253(rport_io_ins_253),
    .io_ins_254(rport_io_ins_254),
    .io_ins_255(rport_io_ins_255),
    .io_ins_256(rport_io_ins_256),
    .io_ins_257(rport_io_ins_257),
    .io_ins_258(rport_io_ins_258),
    .io_ins_259(rport_io_ins_259),
    .io_ins_260(rport_io_ins_260),
    .io_ins_261(rport_io_ins_261),
    .io_ins_262(rport_io_ins_262),
    .io_ins_263(rport_io_ins_263),
    .io_ins_264(rport_io_ins_264),
    .io_ins_265(rport_io_ins_265),
    .io_ins_266(rport_io_ins_266),
    .io_ins_267(rport_io_ins_267),
    .io_ins_268(rport_io_ins_268),
    .io_ins_269(rport_io_ins_269),
    .io_ins_270(rport_io_ins_270),
    .io_ins_271(rport_io_ins_271),
    .io_ins_272(rport_io_ins_272),
    .io_ins_273(rport_io_ins_273),
    .io_ins_274(rport_io_ins_274),
    .io_ins_275(rport_io_ins_275),
    .io_ins_276(rport_io_ins_276),
    .io_ins_277(rport_io_ins_277),
    .io_ins_278(rport_io_ins_278),
    .io_ins_279(rport_io_ins_279),
    .io_ins_280(rport_io_ins_280),
    .io_ins_281(rport_io_ins_281),
    .io_ins_282(rport_io_ins_282),
    .io_ins_283(rport_io_ins_283),
    .io_ins_284(rport_io_ins_284),
    .io_ins_285(rport_io_ins_285),
    .io_ins_286(rport_io_ins_286),
    .io_ins_287(rport_io_ins_287),
    .io_ins_288(rport_io_ins_288),
    .io_ins_289(rport_io_ins_289),
    .io_ins_290(rport_io_ins_290),
    .io_ins_291(rport_io_ins_291),
    .io_ins_292(rport_io_ins_292),
    .io_ins_293(rport_io_ins_293),
    .io_ins_294(rport_io_ins_294),
    .io_ins_295(rport_io_ins_295),
    .io_ins_296(rport_io_ins_296),
    .io_ins_297(rport_io_ins_297),
    .io_ins_298(rport_io_ins_298),
    .io_ins_299(rport_io_ins_299),
    .io_ins_300(rport_io_ins_300),
    .io_ins_301(rport_io_ins_301),
    .io_ins_302(rport_io_ins_302),
    .io_ins_303(rport_io_ins_303),
    .io_ins_304(rport_io_ins_304),
    .io_ins_305(rport_io_ins_305),
    .io_ins_306(rport_io_ins_306),
    .io_ins_307(rport_io_ins_307),
    .io_ins_308(rport_io_ins_308),
    .io_ins_309(rport_io_ins_309),
    .io_ins_310(rport_io_ins_310),
    .io_ins_311(rport_io_ins_311),
    .io_ins_312(rport_io_ins_312),
    .io_ins_313(rport_io_ins_313),
    .io_ins_314(rport_io_ins_314),
    .io_ins_315(rport_io_ins_315),
    .io_ins_316(rport_io_ins_316),
    .io_ins_317(rport_io_ins_317),
    .io_ins_318(rport_io_ins_318),
    .io_ins_319(rport_io_ins_319),
    .io_ins_320(rport_io_ins_320),
    .io_ins_321(rport_io_ins_321),
    .io_ins_322(rport_io_ins_322),
    .io_ins_323(rport_io_ins_323),
    .io_ins_324(rport_io_ins_324),
    .io_ins_325(rport_io_ins_325),
    .io_ins_326(rport_io_ins_326),
    .io_ins_327(rport_io_ins_327),
    .io_ins_328(rport_io_ins_328),
    .io_ins_329(rport_io_ins_329),
    .io_ins_330(rport_io_ins_330),
    .io_ins_331(rport_io_ins_331),
    .io_ins_332(rport_io_ins_332),
    .io_ins_333(rport_io_ins_333),
    .io_ins_334(rport_io_ins_334),
    .io_ins_335(rport_io_ins_335),
    .io_ins_336(rport_io_ins_336),
    .io_ins_337(rport_io_ins_337),
    .io_ins_338(rport_io_ins_338),
    .io_ins_339(rport_io_ins_339),
    .io_ins_340(rport_io_ins_340),
    .io_ins_341(rport_io_ins_341),
    .io_ins_342(rport_io_ins_342),
    .io_ins_343(rport_io_ins_343),
    .io_ins_344(rport_io_ins_344),
    .io_ins_345(rport_io_ins_345),
    .io_ins_346(rport_io_ins_346),
    .io_ins_347(rport_io_ins_347),
    .io_ins_348(rport_io_ins_348),
    .io_ins_349(rport_io_ins_349),
    .io_ins_350(rport_io_ins_350),
    .io_ins_351(rport_io_ins_351),
    .io_ins_352(rport_io_ins_352),
    .io_ins_353(rport_io_ins_353),
    .io_ins_354(rport_io_ins_354),
    .io_ins_355(rport_io_ins_355),
    .io_ins_356(rport_io_ins_356),
    .io_ins_357(rport_io_ins_357),
    .io_ins_358(rport_io_ins_358),
    .io_ins_359(rport_io_ins_359),
    .io_ins_360(rport_io_ins_360),
    .io_ins_361(rport_io_ins_361),
    .io_ins_362(rport_io_ins_362),
    .io_ins_363(rport_io_ins_363),
    .io_ins_364(rport_io_ins_364),
    .io_ins_365(rport_io_ins_365),
    .io_ins_366(rport_io_ins_366),
    .io_ins_367(rport_io_ins_367),
    .io_ins_368(rport_io_ins_368),
    .io_ins_369(rport_io_ins_369),
    .io_ins_370(rport_io_ins_370),
    .io_ins_371(rport_io_ins_371),
    .io_ins_372(rport_io_ins_372),
    .io_ins_373(rport_io_ins_373),
    .io_ins_374(rport_io_ins_374),
    .io_ins_375(rport_io_ins_375),
    .io_ins_376(rport_io_ins_376),
    .io_ins_377(rport_io_ins_377),
    .io_ins_378(rport_io_ins_378),
    .io_ins_379(rport_io_ins_379),
    .io_ins_380(rport_io_ins_380),
    .io_ins_381(rport_io_ins_381),
    .io_ins_382(rport_io_ins_382),
    .io_ins_383(rport_io_ins_383),
    .io_ins_384(rport_io_ins_384),
    .io_ins_385(rport_io_ins_385),
    .io_ins_386(rport_io_ins_386),
    .io_ins_387(rport_io_ins_387),
    .io_ins_388(rport_io_ins_388),
    .io_ins_389(rport_io_ins_389),
    .io_ins_390(rport_io_ins_390),
    .io_ins_391(rport_io_ins_391),
    .io_ins_392(rport_io_ins_392),
    .io_ins_393(rport_io_ins_393),
    .io_ins_394(rport_io_ins_394),
    .io_ins_395(rport_io_ins_395),
    .io_ins_396(rport_io_ins_396),
    .io_ins_397(rport_io_ins_397),
    .io_ins_398(rport_io_ins_398),
    .io_ins_399(rport_io_ins_399),
    .io_ins_400(rport_io_ins_400),
    .io_ins_401(rport_io_ins_401),
    .io_ins_402(rport_io_ins_402),
    .io_ins_403(rport_io_ins_403),
    .io_ins_404(rport_io_ins_404),
    .io_ins_405(rport_io_ins_405),
    .io_ins_406(rport_io_ins_406),
    .io_ins_407(rport_io_ins_407),
    .io_ins_408(rport_io_ins_408),
    .io_ins_409(rport_io_ins_409),
    .io_ins_410(rport_io_ins_410),
    .io_ins_411(rport_io_ins_411),
    .io_ins_412(rport_io_ins_412),
    .io_ins_413(rport_io_ins_413),
    .io_ins_414(rport_io_ins_414),
    .io_ins_415(rport_io_ins_415),
    .io_ins_416(rport_io_ins_416),
    .io_ins_417(rport_io_ins_417),
    .io_ins_418(rport_io_ins_418),
    .io_ins_419(rport_io_ins_419),
    .io_ins_420(rport_io_ins_420),
    .io_ins_421(rport_io_ins_421),
    .io_ins_422(rport_io_ins_422),
    .io_ins_423(rport_io_ins_423),
    .io_ins_424(rport_io_ins_424),
    .io_ins_425(rport_io_ins_425),
    .io_ins_426(rport_io_ins_426),
    .io_ins_427(rport_io_ins_427),
    .io_ins_428(rport_io_ins_428),
    .io_ins_429(rport_io_ins_429),
    .io_ins_430(rport_io_ins_430),
    .io_ins_431(rport_io_ins_431),
    .io_ins_432(rport_io_ins_432),
    .io_ins_433(rport_io_ins_433),
    .io_ins_434(rport_io_ins_434),
    .io_ins_435(rport_io_ins_435),
    .io_ins_436(rport_io_ins_436),
    .io_ins_437(rport_io_ins_437),
    .io_ins_438(rport_io_ins_438),
    .io_ins_439(rport_io_ins_439),
    .io_ins_440(rport_io_ins_440),
    .io_ins_441(rport_io_ins_441),
    .io_ins_442(rport_io_ins_442),
    .io_ins_443(rport_io_ins_443),
    .io_ins_444(rport_io_ins_444),
    .io_ins_445(rport_io_ins_445),
    .io_ins_446(rport_io_ins_446),
    .io_ins_447(rport_io_ins_447),
    .io_ins_448(rport_io_ins_448),
    .io_ins_449(rport_io_ins_449),
    .io_ins_450(rport_io_ins_450),
    .io_ins_451(rport_io_ins_451),
    .io_ins_452(rport_io_ins_452),
    .io_ins_453(rport_io_ins_453),
    .io_ins_454(rport_io_ins_454),
    .io_ins_455(rport_io_ins_455),
    .io_ins_456(rport_io_ins_456),
    .io_ins_457(rport_io_ins_457),
    .io_ins_458(rport_io_ins_458),
    .io_ins_459(rport_io_ins_459),
    .io_ins_460(rport_io_ins_460),
    .io_ins_461(rport_io_ins_461),
    .io_ins_462(rport_io_ins_462),
    .io_ins_463(rport_io_ins_463),
    .io_ins_464(rport_io_ins_464),
    .io_ins_465(rport_io_ins_465),
    .io_ins_466(rport_io_ins_466),
    .io_ins_467(rport_io_ins_467),
    .io_ins_468(rport_io_ins_468),
    .io_ins_469(rport_io_ins_469),
    .io_ins_470(rport_io_ins_470),
    .io_ins_471(rport_io_ins_471),
    .io_ins_472(rport_io_ins_472),
    .io_ins_473(rport_io_ins_473),
    .io_ins_474(rport_io_ins_474),
    .io_ins_475(rport_io_ins_475),
    .io_ins_476(rport_io_ins_476),
    .io_ins_477(rport_io_ins_477),
    .io_ins_478(rport_io_ins_478),
    .io_ins_479(rport_io_ins_479),
    .io_ins_480(rport_io_ins_480),
    .io_ins_481(rport_io_ins_481),
    .io_ins_482(rport_io_ins_482),
    .io_ins_483(rport_io_ins_483),
    .io_ins_484(rport_io_ins_484),
    .io_ins_485(rport_io_ins_485),
    .io_ins_486(rport_io_ins_486),
    .io_ins_487(rport_io_ins_487),
    .io_ins_488(rport_io_ins_488),
    .io_ins_489(rport_io_ins_489),
    .io_ins_490(rport_io_ins_490),
    .io_ins_491(rport_io_ins_491),
    .io_ins_492(rport_io_ins_492),
    .io_ins_493(rport_io_ins_493),
    .io_ins_494(rport_io_ins_494),
    .io_ins_495(rport_io_ins_495),
    .io_ins_496(rport_io_ins_496),
    .io_ins_497(rport_io_ins_497),
    .io_ins_498(rport_io_ins_498),
    .io_ins_499(rport_io_ins_499),
    .io_ins_500(rport_io_ins_500),
    .io_ins_501(rport_io_ins_501),
    .io_ins_502(rport_io_ins_502),
    .io_ins_503(rport_io_ins_503),
    .io_ins_504(rport_io_ins_504),
    .io_ins_505(rport_io_ins_505),
    .io_ins_506(rport_io_ins_506),
    .io_ins_507(rport_io_ins_507),
    .io_ins_508(rport_io_ins_508),
    .io_ins_509(rport_io_ins_509),
    .io_ins_510(rport_io_ins_510),
    .io_ins_511(rport_io_ins_511),
    .io_ins_512(rport_io_ins_512),
    .io_ins_513(rport_io_ins_513),
    .io_ins_514(rport_io_ins_514),
    .io_ins_515(rport_io_ins_515),
    .io_ins_516(rport_io_ins_516),
    .io_ins_517(rport_io_ins_517),
    .io_sel(rport_io_sel),
    .io_out(rport_io_out)
  );
  assign _T_3166 = io_waddr == 32'h0; // @[RegFile.scala 80:42:@49732.4]
  assign _T_3172 = io_waddr == 32'h1; // @[RegFile.scala 68:46:@49744.4]
  assign _T_3173 = io_wen & _T_3172; // @[RegFile.scala 68:34:@49745.4]
  assign _T_3186 = io_waddr == 32'h2; // @[RegFile.scala 80:42:@49763.4]
  assign _T_3192 = io_waddr == 32'h3; // @[RegFile.scala 74:80:@49775.4]
  assign _T_3193 = io_wen & _T_3192; // @[RegFile.scala 74:68:@49776.4]
  assign _T_3199 = io_waddr == 32'h4; // @[RegFile.scala 74:80:@49789.4]
  assign _T_3200 = io_wen & _T_3199; // @[RegFile.scala 74:68:@49790.4]
  assign _T_3206 = io_waddr == 32'h5; // @[RegFile.scala 74:80:@49803.4]
  assign _T_3207 = io_wen & _T_3206; // @[RegFile.scala 74:68:@49804.4]
  assign _T_3213 = io_waddr == 32'h6; // @[RegFile.scala 74:80:@49817.4]
  assign _T_3214 = io_wen & _T_3213; // @[RegFile.scala 74:68:@49818.4]
  assign _T_3220 = io_waddr == 32'h7; // @[RegFile.scala 74:80:@49831.4]
  assign _T_3221 = io_wen & _T_3220; // @[RegFile.scala 74:68:@49832.4]
  assign _T_3227 = io_waddr == 32'h8; // @[RegFile.scala 74:80:@49845.4]
  assign _T_3228 = io_wen & _T_3227; // @[RegFile.scala 74:68:@49846.4]
  assign _T_3234 = io_waddr == 32'h9; // @[RegFile.scala 74:80:@49859.4]
  assign _T_3235 = io_wen & _T_3234; // @[RegFile.scala 74:68:@49860.4]
  assign _T_3241 = io_waddr == 32'ha; // @[RegFile.scala 74:80:@49873.4]
  assign _T_3242 = io_wen & _T_3241; // @[RegFile.scala 74:68:@49874.4]
  assign _T_3248 = io_waddr == 32'hb; // @[RegFile.scala 74:80:@49887.4]
  assign _T_3249 = io_wen & _T_3248; // @[RegFile.scala 74:68:@49888.4]
  assign _T_3255 = io_waddr == 32'hc; // @[RegFile.scala 74:80:@49901.4]
  assign _T_3256 = io_wen & _T_3255; // @[RegFile.scala 74:68:@49902.4]
  assign _T_3262 = io_waddr == 32'hd; // @[RegFile.scala 74:80:@49915.4]
  assign _T_3263 = io_wen & _T_3262; // @[RegFile.scala 74:68:@49916.4]
  assign _T_3269 = io_waddr == 32'he; // @[RegFile.scala 74:80:@49929.4]
  assign _T_3270 = io_wen & _T_3269; // @[RegFile.scala 74:68:@49930.4]
  assign _T_3276 = io_waddr == 32'hf; // @[RegFile.scala 74:80:@49943.4]
  assign _T_3277 = io_wen & _T_3276; // @[RegFile.scala 74:68:@49944.4]
  assign _T_3283 = io_waddr == 32'h10; // @[RegFile.scala 74:80:@49957.4]
  assign _T_3284 = io_wen & _T_3283; // @[RegFile.scala 74:68:@49958.4]
  assign _T_3290 = io_waddr == 32'h11; // @[RegFile.scala 74:80:@49971.4]
  assign _T_3291 = io_wen & _T_3290; // @[RegFile.scala 74:68:@49972.4]
  assign _T_3297 = io_waddr == 32'h12; // @[RegFile.scala 74:80:@49985.4]
  assign _T_3298 = io_wen & _T_3297; // @[RegFile.scala 74:68:@49986.4]
  assign io_rdata = rport_io_out; // @[RegFile.scala 107:14:@58023.4]
  assign io_argIns_0 = regs_0_io_out; // @[RegFile.scala 111:13:@58028.4]
  assign io_argIns_1 = regs_1_io_out; // @[RegFile.scala 111:13:@58029.4]
  assign io_argIns_2 = regs_2_io_out; // @[RegFile.scala 111:13:@58030.4]
  assign regs_0_clock = clock; // @[:@49730.4]
  assign regs_0_reset = reset; // @[:@49731.4 RegFile.scala 82:16:@49737.4]
  assign regs_0_io_in = io_wdata; // @[RegFile.scala 81:16:@49735.4]
  assign regs_0_io_reset = reset; // @[RegFile.scala 83:19:@49739.4]
  assign regs_0_io_enable = io_wen & _T_3166; // @[RegFile.scala 80:20:@49734.4]
  assign regs_1_clock = clock; // @[:@49742.4]
  assign regs_1_reset = reset; // @[:@49743.4 RegFile.scala 70:16:@49755.4]
  assign regs_1_io_in = _T_3173 ? io_wdata : io_argOuts_0_bits; // @[RegFile.scala 69:16:@49753.4]
  assign regs_1_io_reset = reset; // @[RegFile.scala 72:19:@49758.4]
  assign regs_1_io_enable = _T_3173 ? _T_3173 : io_argOuts_0_valid; // @[RegFile.scala 68:20:@49749.4]
  assign regs_2_clock = clock; // @[:@49761.4]
  assign regs_2_reset = reset; // @[:@49762.4 RegFile.scala 82:16:@49768.4]
  assign regs_2_io_in = io_wdata; // @[RegFile.scala 81:16:@49766.4]
  assign regs_2_io_reset = reset; // @[RegFile.scala 83:19:@49770.4]
  assign regs_2_io_enable = io_wen & _T_3186; // @[RegFile.scala 80:20:@49765.4]
  assign regs_3_clock = clock; // @[:@49773.4]
  assign regs_3_reset = io_reset; // @[:@49774.4 RegFile.scala 76:16:@49781.4]
  assign regs_3_io_in = io_argOuts_1_valid ? io_argOuts_1_bits : io_wdata; // @[RegFile.scala 75:16:@49780.4]
  assign regs_3_io_reset = reset; // @[RegFile.scala 78:19:@49784.4]
  assign regs_3_io_enable = io_argOuts_1_valid | _T_3193; // @[RegFile.scala 74:20:@49778.4]
  assign regs_4_clock = clock; // @[:@49787.4]
  assign regs_4_reset = io_reset; // @[:@49788.4 RegFile.scala 76:16:@49795.4]
  assign regs_4_io_in = io_argOuts_2_valid ? io_argOuts_2_bits : io_wdata; // @[RegFile.scala 75:16:@49794.4]
  assign regs_4_io_reset = reset; // @[RegFile.scala 78:19:@49798.4]
  assign regs_4_io_enable = io_argOuts_2_valid | _T_3200; // @[RegFile.scala 74:20:@49792.4]
  assign regs_5_clock = clock; // @[:@49801.4]
  assign regs_5_reset = io_reset; // @[:@49802.4 RegFile.scala 76:16:@49809.4]
  assign regs_5_io_in = io_argOuts_3_valid ? io_argOuts_3_bits : io_wdata; // @[RegFile.scala 75:16:@49808.4]
  assign regs_5_io_reset = reset; // @[RegFile.scala 78:19:@49812.4]
  assign regs_5_io_enable = io_argOuts_3_valid | _T_3207; // @[RegFile.scala 74:20:@49806.4]
  assign regs_6_clock = clock; // @[:@49815.4]
  assign regs_6_reset = io_reset; // @[:@49816.4 RegFile.scala 76:16:@49823.4]
  assign regs_6_io_in = io_argOuts_4_valid ? io_argOuts_4_bits : io_wdata; // @[RegFile.scala 75:16:@49822.4]
  assign regs_6_io_reset = reset; // @[RegFile.scala 78:19:@49826.4]
  assign regs_6_io_enable = io_argOuts_4_valid | _T_3214; // @[RegFile.scala 74:20:@49820.4]
  assign regs_7_clock = clock; // @[:@49829.4]
  assign regs_7_reset = io_reset; // @[:@49830.4 RegFile.scala 76:16:@49837.4]
  assign regs_7_io_in = io_argOuts_5_valid ? io_argOuts_5_bits : io_wdata; // @[RegFile.scala 75:16:@49836.4]
  assign regs_7_io_reset = reset; // @[RegFile.scala 78:19:@49840.4]
  assign regs_7_io_enable = io_argOuts_5_valid | _T_3221; // @[RegFile.scala 74:20:@49834.4]
  assign regs_8_clock = clock; // @[:@49843.4]
  assign regs_8_reset = io_reset; // @[:@49844.4 RegFile.scala 76:16:@49851.4]
  assign regs_8_io_in = io_argOuts_6_valid ? io_argOuts_6_bits : io_wdata; // @[RegFile.scala 75:16:@49850.4]
  assign regs_8_io_reset = reset; // @[RegFile.scala 78:19:@49854.4]
  assign regs_8_io_enable = io_argOuts_6_valid | _T_3228; // @[RegFile.scala 74:20:@49848.4]
  assign regs_9_clock = clock; // @[:@49857.4]
  assign regs_9_reset = io_reset; // @[:@49858.4 RegFile.scala 76:16:@49865.4]
  assign regs_9_io_in = io_argOuts_7_valid ? io_argOuts_7_bits : io_wdata; // @[RegFile.scala 75:16:@49864.4]
  assign regs_9_io_reset = reset; // @[RegFile.scala 78:19:@49868.4]
  assign regs_9_io_enable = io_argOuts_7_valid | _T_3235; // @[RegFile.scala 74:20:@49862.4]
  assign regs_10_clock = clock; // @[:@49871.4]
  assign regs_10_reset = io_reset; // @[:@49872.4 RegFile.scala 76:16:@49879.4]
  assign regs_10_io_in = io_argOuts_8_valid ? io_argOuts_8_bits : io_wdata; // @[RegFile.scala 75:16:@49878.4]
  assign regs_10_io_reset = reset; // @[RegFile.scala 78:19:@49882.4]
  assign regs_10_io_enable = io_argOuts_8_valid | _T_3242; // @[RegFile.scala 74:20:@49876.4]
  assign regs_11_clock = clock; // @[:@49885.4]
  assign regs_11_reset = io_reset; // @[:@49886.4 RegFile.scala 76:16:@49893.4]
  assign regs_11_io_in = io_argOuts_9_valid ? io_argOuts_9_bits : io_wdata; // @[RegFile.scala 75:16:@49892.4]
  assign regs_11_io_reset = reset; // @[RegFile.scala 78:19:@49896.4]
  assign regs_11_io_enable = io_argOuts_9_valid | _T_3249; // @[RegFile.scala 74:20:@49890.4]
  assign regs_12_clock = clock; // @[:@49899.4]
  assign regs_12_reset = io_reset; // @[:@49900.4 RegFile.scala 76:16:@49907.4]
  assign regs_12_io_in = io_argOuts_10_valid ? io_argOuts_10_bits : io_wdata; // @[RegFile.scala 75:16:@49906.4]
  assign regs_12_io_reset = reset; // @[RegFile.scala 78:19:@49910.4]
  assign regs_12_io_enable = io_argOuts_10_valid | _T_3256; // @[RegFile.scala 74:20:@49904.4]
  assign regs_13_clock = clock; // @[:@49913.4]
  assign regs_13_reset = io_reset; // @[:@49914.4 RegFile.scala 76:16:@49921.4]
  assign regs_13_io_in = io_argOuts_11_valid ? io_argOuts_11_bits : io_wdata; // @[RegFile.scala 75:16:@49920.4]
  assign regs_13_io_reset = reset; // @[RegFile.scala 78:19:@49924.4]
  assign regs_13_io_enable = io_argOuts_11_valid | _T_3263; // @[RegFile.scala 74:20:@49918.4]
  assign regs_14_clock = clock; // @[:@49927.4]
  assign regs_14_reset = io_reset; // @[:@49928.4 RegFile.scala 76:16:@49935.4]
  assign regs_14_io_in = io_argOuts_12_valid ? io_argOuts_12_bits : io_wdata; // @[RegFile.scala 75:16:@49934.4]
  assign regs_14_io_reset = reset; // @[RegFile.scala 78:19:@49938.4]
  assign regs_14_io_enable = io_argOuts_12_valid | _T_3270; // @[RegFile.scala 74:20:@49932.4]
  assign regs_15_clock = clock; // @[:@49941.4]
  assign regs_15_reset = io_reset; // @[:@49942.4 RegFile.scala 76:16:@49949.4]
  assign regs_15_io_in = io_argOuts_13_valid ? io_argOuts_13_bits : io_wdata; // @[RegFile.scala 75:16:@49948.4]
  assign regs_15_io_reset = reset; // @[RegFile.scala 78:19:@49952.4]
  assign regs_15_io_enable = io_argOuts_13_valid | _T_3277; // @[RegFile.scala 74:20:@49946.4]
  assign regs_16_clock = clock; // @[:@49955.4]
  assign regs_16_reset = io_reset; // @[:@49956.4 RegFile.scala 76:16:@49963.4]
  assign regs_16_io_in = io_argOuts_14_valid ? io_argOuts_14_bits : io_wdata; // @[RegFile.scala 75:16:@49962.4]
  assign regs_16_io_reset = reset; // @[RegFile.scala 78:19:@49966.4]
  assign regs_16_io_enable = io_argOuts_14_valid | _T_3284; // @[RegFile.scala 74:20:@49960.4]
  assign regs_17_clock = clock; // @[:@49969.4]
  assign regs_17_reset = io_reset; // @[:@49970.4 RegFile.scala 76:16:@49977.4]
  assign regs_17_io_in = io_argOuts_15_valid ? io_argOuts_15_bits : io_wdata; // @[RegFile.scala 75:16:@49976.4]
  assign regs_17_io_reset = reset; // @[RegFile.scala 78:19:@49980.4]
  assign regs_17_io_enable = io_argOuts_15_valid | _T_3291; // @[RegFile.scala 74:20:@49974.4]
  assign regs_18_clock = clock; // @[:@49983.4]
  assign regs_18_reset = io_reset; // @[:@49984.4 RegFile.scala 76:16:@49991.4]
  assign regs_18_io_in = io_argOuts_16_valid ? io_argOuts_16_bits : io_wdata; // @[RegFile.scala 75:16:@49990.4]
  assign regs_18_io_reset = reset; // @[RegFile.scala 78:19:@49994.4]
  assign regs_18_io_enable = io_argOuts_16_valid | _T_3298; // @[RegFile.scala 74:20:@49988.4]
  assign regs_19_clock = clock; // @[:@49997.4]
  assign regs_19_reset = io_reset; // @[:@49998.4 RegFile.scala 76:16:@50005.4]
  assign regs_19_io_in = io_argOuts_17_bits; // @[RegFile.scala 75:16:@50004.4]
  assign regs_19_io_reset = reset; // @[RegFile.scala 78:19:@50008.4]
  assign regs_19_io_enable = 1'h1; // @[RegFile.scala 74:20:@50002.4]
  assign regs_20_clock = clock; // @[:@50011.4]
  assign regs_20_reset = io_reset; // @[:@50012.4 RegFile.scala 76:16:@50019.4]
  assign regs_20_io_in = io_argOuts_18_bits; // @[RegFile.scala 75:16:@50018.4]
  assign regs_20_io_reset = reset; // @[RegFile.scala 78:19:@50022.4]
  assign regs_20_io_enable = 1'h1; // @[RegFile.scala 74:20:@50016.4]
  assign regs_21_clock = clock; // @[:@50025.4]
  assign regs_21_reset = io_reset; // @[:@50026.4 RegFile.scala 76:16:@50033.4]
  assign regs_21_io_in = io_argOuts_19_bits; // @[RegFile.scala 75:16:@50032.4]
  assign regs_21_io_reset = reset; // @[RegFile.scala 78:19:@50036.4]
  assign regs_21_io_enable = 1'h1; // @[RegFile.scala 74:20:@50030.4]
  assign regs_22_clock = clock; // @[:@50039.4]
  assign regs_22_reset = io_reset; // @[:@50040.4 RegFile.scala 76:16:@50047.4]
  assign regs_22_io_in = io_argOuts_20_bits; // @[RegFile.scala 75:16:@50046.4]
  assign regs_22_io_reset = reset; // @[RegFile.scala 78:19:@50050.4]
  assign regs_22_io_enable = 1'h1; // @[RegFile.scala 74:20:@50044.4]
  assign regs_23_clock = clock; // @[:@50053.4]
  assign regs_23_reset = io_reset; // @[:@50054.4 RegFile.scala 76:16:@50061.4]
  assign regs_23_io_in = io_argOuts_21_bits; // @[RegFile.scala 75:16:@50060.4]
  assign regs_23_io_reset = reset; // @[RegFile.scala 78:19:@50064.4]
  assign regs_23_io_enable = 1'h1; // @[RegFile.scala 74:20:@50058.4]
  assign regs_24_clock = clock; // @[:@50067.4]
  assign regs_24_reset = io_reset; // @[:@50068.4 RegFile.scala 76:16:@50075.4]
  assign regs_24_io_in = io_argOuts_22_bits; // @[RegFile.scala 75:16:@50074.4]
  assign regs_24_io_reset = reset; // @[RegFile.scala 78:19:@50078.4]
  assign regs_24_io_enable = 1'h1; // @[RegFile.scala 74:20:@50072.4]
  assign regs_25_clock = clock; // @[:@50081.4]
  assign regs_25_reset = io_reset; // @[:@50082.4 RegFile.scala 76:16:@50089.4]
  assign regs_25_io_in = io_argOuts_23_bits; // @[RegFile.scala 75:16:@50088.4]
  assign regs_25_io_reset = reset; // @[RegFile.scala 78:19:@50092.4]
  assign regs_25_io_enable = 1'h1; // @[RegFile.scala 74:20:@50086.4]
  assign regs_26_clock = clock; // @[:@50095.4]
  assign regs_26_reset = io_reset; // @[:@50096.4 RegFile.scala 76:16:@50103.4]
  assign regs_26_io_in = io_argOuts_24_bits; // @[RegFile.scala 75:16:@50102.4]
  assign regs_26_io_reset = reset; // @[RegFile.scala 78:19:@50106.4]
  assign regs_26_io_enable = 1'h1; // @[RegFile.scala 74:20:@50100.4]
  assign regs_27_clock = clock; // @[:@50109.4]
  assign regs_27_reset = io_reset; // @[:@50110.4 RegFile.scala 76:16:@50117.4]
  assign regs_27_io_in = io_argOuts_25_bits; // @[RegFile.scala 75:16:@50116.4]
  assign regs_27_io_reset = reset; // @[RegFile.scala 78:19:@50120.4]
  assign regs_27_io_enable = 1'h1; // @[RegFile.scala 74:20:@50114.4]
  assign regs_28_clock = clock; // @[:@50123.4]
  assign regs_28_reset = io_reset; // @[:@50124.4 RegFile.scala 76:16:@50131.4]
  assign regs_28_io_in = io_argOuts_26_bits; // @[RegFile.scala 75:16:@50130.4]
  assign regs_28_io_reset = reset; // @[RegFile.scala 78:19:@50134.4]
  assign regs_28_io_enable = 1'h1; // @[RegFile.scala 74:20:@50128.4]
  assign regs_29_clock = clock; // @[:@50137.4]
  assign regs_29_reset = io_reset; // @[:@50138.4 RegFile.scala 76:16:@50145.4]
  assign regs_29_io_in = io_argOuts_27_bits; // @[RegFile.scala 75:16:@50144.4]
  assign regs_29_io_reset = reset; // @[RegFile.scala 78:19:@50148.4]
  assign regs_29_io_enable = 1'h1; // @[RegFile.scala 74:20:@50142.4]
  assign regs_30_clock = clock; // @[:@50151.4]
  assign regs_30_reset = io_reset; // @[:@50152.4 RegFile.scala 76:16:@50159.4]
  assign regs_30_io_in = io_argOuts_28_bits; // @[RegFile.scala 75:16:@50158.4]
  assign regs_30_io_reset = reset; // @[RegFile.scala 78:19:@50162.4]
  assign regs_30_io_enable = 1'h1; // @[RegFile.scala 74:20:@50156.4]
  assign regs_31_clock = clock; // @[:@50165.4]
  assign regs_31_reset = io_reset; // @[:@50166.4 RegFile.scala 76:16:@50173.4]
  assign regs_31_io_in = io_argOuts_29_bits; // @[RegFile.scala 75:16:@50172.4]
  assign regs_31_io_reset = reset; // @[RegFile.scala 78:19:@50176.4]
  assign regs_31_io_enable = 1'h1; // @[RegFile.scala 74:20:@50170.4]
  assign regs_32_clock = clock; // @[:@50179.4]
  assign regs_32_reset = io_reset; // @[:@50180.4 RegFile.scala 76:16:@50187.4]
  assign regs_32_io_in = io_argOuts_30_bits; // @[RegFile.scala 75:16:@50186.4]
  assign regs_32_io_reset = reset; // @[RegFile.scala 78:19:@50190.4]
  assign regs_32_io_enable = 1'h1; // @[RegFile.scala 74:20:@50184.4]
  assign regs_33_clock = clock; // @[:@50193.4]
  assign regs_33_reset = io_reset; // @[:@50194.4 RegFile.scala 76:16:@50201.4]
  assign regs_33_io_in = io_argOuts_31_bits; // @[RegFile.scala 75:16:@50200.4]
  assign regs_33_io_reset = reset; // @[RegFile.scala 78:19:@50204.4]
  assign regs_33_io_enable = 1'h1; // @[RegFile.scala 74:20:@50198.4]
  assign regs_34_clock = clock; // @[:@50207.4]
  assign regs_34_reset = io_reset; // @[:@50208.4 RegFile.scala 76:16:@50215.4]
  assign regs_34_io_in = io_argOuts_32_bits; // @[RegFile.scala 75:16:@50214.4]
  assign regs_34_io_reset = reset; // @[RegFile.scala 78:19:@50218.4]
  assign regs_34_io_enable = 1'h1; // @[RegFile.scala 74:20:@50212.4]
  assign regs_35_clock = clock; // @[:@50221.4]
  assign regs_35_reset = io_reset; // @[:@50222.4 RegFile.scala 76:16:@50229.4]
  assign regs_35_io_in = io_argOuts_33_bits; // @[RegFile.scala 75:16:@50228.4]
  assign regs_35_io_reset = reset; // @[RegFile.scala 78:19:@50232.4]
  assign regs_35_io_enable = 1'h1; // @[RegFile.scala 74:20:@50226.4]
  assign regs_36_clock = clock; // @[:@50235.4]
  assign regs_36_reset = io_reset; // @[:@50236.4 RegFile.scala 76:16:@50243.4]
  assign regs_36_io_in = io_argOuts_34_bits; // @[RegFile.scala 75:16:@50242.4]
  assign regs_36_io_reset = reset; // @[RegFile.scala 78:19:@50246.4]
  assign regs_36_io_enable = 1'h1; // @[RegFile.scala 74:20:@50240.4]
  assign regs_37_clock = clock; // @[:@50249.4]
  assign regs_37_reset = io_reset; // @[:@50250.4 RegFile.scala 76:16:@50257.4]
  assign regs_37_io_in = io_argOuts_35_bits; // @[RegFile.scala 75:16:@50256.4]
  assign regs_37_io_reset = reset; // @[RegFile.scala 78:19:@50260.4]
  assign regs_37_io_enable = 1'h1; // @[RegFile.scala 74:20:@50254.4]
  assign regs_38_clock = clock; // @[:@50263.4]
  assign regs_38_reset = io_reset; // @[:@50264.4 RegFile.scala 76:16:@50271.4]
  assign regs_38_io_in = io_argOuts_36_bits; // @[RegFile.scala 75:16:@50270.4]
  assign regs_38_io_reset = reset; // @[RegFile.scala 78:19:@50274.4]
  assign regs_38_io_enable = 1'h1; // @[RegFile.scala 74:20:@50268.4]
  assign regs_39_clock = clock; // @[:@50277.4]
  assign regs_39_reset = io_reset; // @[:@50278.4 RegFile.scala 76:16:@50285.4]
  assign regs_39_io_in = io_argOuts_37_bits; // @[RegFile.scala 75:16:@50284.4]
  assign regs_39_io_reset = reset; // @[RegFile.scala 78:19:@50288.4]
  assign regs_39_io_enable = 1'h1; // @[RegFile.scala 74:20:@50282.4]
  assign regs_40_clock = clock; // @[:@50291.4]
  assign regs_40_reset = io_reset; // @[:@50292.4 RegFile.scala 76:16:@50299.4]
  assign regs_40_io_in = io_argOuts_38_bits; // @[RegFile.scala 75:16:@50298.4]
  assign regs_40_io_reset = reset; // @[RegFile.scala 78:19:@50302.4]
  assign regs_40_io_enable = 1'h1; // @[RegFile.scala 74:20:@50296.4]
  assign regs_41_clock = clock; // @[:@50305.4]
  assign regs_41_reset = io_reset; // @[:@50306.4 RegFile.scala 76:16:@50313.4]
  assign regs_41_io_in = io_argOuts_39_bits; // @[RegFile.scala 75:16:@50312.4]
  assign regs_41_io_reset = reset; // @[RegFile.scala 78:19:@50316.4]
  assign regs_41_io_enable = 1'h1; // @[RegFile.scala 74:20:@50310.4]
  assign regs_42_clock = clock; // @[:@50319.4]
  assign regs_42_reset = io_reset; // @[:@50320.4 RegFile.scala 76:16:@50327.4]
  assign regs_42_io_in = io_argOuts_40_bits; // @[RegFile.scala 75:16:@50326.4]
  assign regs_42_io_reset = reset; // @[RegFile.scala 78:19:@50330.4]
  assign regs_42_io_enable = 1'h1; // @[RegFile.scala 74:20:@50324.4]
  assign regs_43_clock = clock; // @[:@50333.4]
  assign regs_43_reset = io_reset; // @[:@50334.4 RegFile.scala 76:16:@50341.4]
  assign regs_43_io_in = io_argOuts_41_bits; // @[RegFile.scala 75:16:@50340.4]
  assign regs_43_io_reset = reset; // @[RegFile.scala 78:19:@50344.4]
  assign regs_43_io_enable = 1'h1; // @[RegFile.scala 74:20:@50338.4]
  assign regs_44_clock = clock; // @[:@50347.4]
  assign regs_44_reset = io_reset; // @[:@50348.4 RegFile.scala 76:16:@50355.4]
  assign regs_44_io_in = io_argOuts_42_bits; // @[RegFile.scala 75:16:@50354.4]
  assign regs_44_io_reset = reset; // @[RegFile.scala 78:19:@50358.4]
  assign regs_44_io_enable = 1'h1; // @[RegFile.scala 74:20:@50352.4]
  assign regs_45_clock = clock; // @[:@50361.4]
  assign regs_45_reset = io_reset; // @[:@50362.4 RegFile.scala 76:16:@50369.4]
  assign regs_45_io_in = io_argOuts_43_bits; // @[RegFile.scala 75:16:@50368.4]
  assign regs_45_io_reset = reset; // @[RegFile.scala 78:19:@50372.4]
  assign regs_45_io_enable = 1'h1; // @[RegFile.scala 74:20:@50366.4]
  assign regs_46_clock = clock; // @[:@50375.4]
  assign regs_46_reset = io_reset; // @[:@50376.4 RegFile.scala 76:16:@50383.4]
  assign regs_46_io_in = io_argOuts_44_bits; // @[RegFile.scala 75:16:@50382.4]
  assign regs_46_io_reset = reset; // @[RegFile.scala 78:19:@50386.4]
  assign regs_46_io_enable = 1'h1; // @[RegFile.scala 74:20:@50380.4]
  assign regs_47_clock = clock; // @[:@50389.4]
  assign regs_47_reset = io_reset; // @[:@50390.4 RegFile.scala 76:16:@50397.4]
  assign regs_47_io_in = io_argOuts_45_bits; // @[RegFile.scala 75:16:@50396.4]
  assign regs_47_io_reset = reset; // @[RegFile.scala 78:19:@50400.4]
  assign regs_47_io_enable = 1'h1; // @[RegFile.scala 74:20:@50394.4]
  assign regs_48_clock = clock; // @[:@50403.4]
  assign regs_48_reset = io_reset; // @[:@50404.4 RegFile.scala 76:16:@50411.4]
  assign regs_48_io_in = io_argOuts_46_bits; // @[RegFile.scala 75:16:@50410.4]
  assign regs_48_io_reset = reset; // @[RegFile.scala 78:19:@50414.4]
  assign regs_48_io_enable = 1'h1; // @[RegFile.scala 74:20:@50408.4]
  assign regs_49_clock = clock; // @[:@50417.4]
  assign regs_49_reset = io_reset; // @[:@50418.4 RegFile.scala 76:16:@50425.4]
  assign regs_49_io_in = 64'h0; // @[RegFile.scala 75:16:@50424.4]
  assign regs_49_io_reset = reset; // @[RegFile.scala 78:19:@50428.4]
  assign regs_49_io_enable = 1'h1; // @[RegFile.scala 74:20:@50422.4]
  assign regs_50_clock = clock; // @[:@50431.4]
  assign regs_50_reset = io_reset; // @[:@50432.4 RegFile.scala 76:16:@50439.4]
  assign regs_50_io_in = 64'h0; // @[RegFile.scala 75:16:@50438.4]
  assign regs_50_io_reset = reset; // @[RegFile.scala 78:19:@50442.4]
  assign regs_50_io_enable = 1'h1; // @[RegFile.scala 74:20:@50436.4]
  assign regs_51_clock = clock; // @[:@50445.4]
  assign regs_51_reset = io_reset; // @[:@50446.4 RegFile.scala 76:16:@50453.4]
  assign regs_51_io_in = 64'h0; // @[RegFile.scala 75:16:@50452.4]
  assign regs_51_io_reset = reset; // @[RegFile.scala 78:19:@50456.4]
  assign regs_51_io_enable = 1'h1; // @[RegFile.scala 74:20:@50450.4]
  assign regs_52_clock = clock; // @[:@50459.4]
  assign regs_52_reset = io_reset; // @[:@50460.4 RegFile.scala 76:16:@50467.4]
  assign regs_52_io_in = 64'h0; // @[RegFile.scala 75:16:@50466.4]
  assign regs_52_io_reset = reset; // @[RegFile.scala 78:19:@50470.4]
  assign regs_52_io_enable = 1'h1; // @[RegFile.scala 74:20:@50464.4]
  assign regs_53_clock = clock; // @[:@50473.4]
  assign regs_53_reset = io_reset; // @[:@50474.4 RegFile.scala 76:16:@50481.4]
  assign regs_53_io_in = 64'h0; // @[RegFile.scala 75:16:@50480.4]
  assign regs_53_io_reset = reset; // @[RegFile.scala 78:19:@50484.4]
  assign regs_53_io_enable = 1'h1; // @[RegFile.scala 74:20:@50478.4]
  assign regs_54_clock = clock; // @[:@50487.4]
  assign regs_54_reset = io_reset; // @[:@50488.4 RegFile.scala 76:16:@50495.4]
  assign regs_54_io_in = 64'h0; // @[RegFile.scala 75:16:@50494.4]
  assign regs_54_io_reset = reset; // @[RegFile.scala 78:19:@50498.4]
  assign regs_54_io_enable = 1'h1; // @[RegFile.scala 74:20:@50492.4]
  assign regs_55_clock = clock; // @[:@50501.4]
  assign regs_55_reset = io_reset; // @[:@50502.4 RegFile.scala 76:16:@50509.4]
  assign regs_55_io_in = 64'h0; // @[RegFile.scala 75:16:@50508.4]
  assign regs_55_io_reset = reset; // @[RegFile.scala 78:19:@50512.4]
  assign regs_55_io_enable = 1'h1; // @[RegFile.scala 74:20:@50506.4]
  assign regs_56_clock = clock; // @[:@50515.4]
  assign regs_56_reset = io_reset; // @[:@50516.4 RegFile.scala 76:16:@50523.4]
  assign regs_56_io_in = 64'h0; // @[RegFile.scala 75:16:@50522.4]
  assign regs_56_io_reset = reset; // @[RegFile.scala 78:19:@50526.4]
  assign regs_56_io_enable = 1'h1; // @[RegFile.scala 74:20:@50520.4]
  assign regs_57_clock = clock; // @[:@50529.4]
  assign regs_57_reset = io_reset; // @[:@50530.4 RegFile.scala 76:16:@50537.4]
  assign regs_57_io_in = 64'h0; // @[RegFile.scala 75:16:@50536.4]
  assign regs_57_io_reset = reset; // @[RegFile.scala 78:19:@50540.4]
  assign regs_57_io_enable = 1'h1; // @[RegFile.scala 74:20:@50534.4]
  assign regs_58_clock = clock; // @[:@50543.4]
  assign regs_58_reset = io_reset; // @[:@50544.4 RegFile.scala 76:16:@50551.4]
  assign regs_58_io_in = 64'h0; // @[RegFile.scala 75:16:@50550.4]
  assign regs_58_io_reset = reset; // @[RegFile.scala 78:19:@50554.4]
  assign regs_58_io_enable = 1'h1; // @[RegFile.scala 74:20:@50548.4]
  assign regs_59_clock = clock; // @[:@50557.4]
  assign regs_59_reset = io_reset; // @[:@50558.4 RegFile.scala 76:16:@50565.4]
  assign regs_59_io_in = io_argOuts_57_bits; // @[RegFile.scala 75:16:@50564.4]
  assign regs_59_io_reset = reset; // @[RegFile.scala 78:19:@50568.4]
  assign regs_59_io_enable = 1'h1; // @[RegFile.scala 74:20:@50562.4]
  assign regs_60_clock = clock; // @[:@50571.4]
  assign regs_60_reset = io_reset; // @[:@50572.4 RegFile.scala 76:16:@50579.4]
  assign regs_60_io_in = 64'h0; // @[RegFile.scala 75:16:@50578.4]
  assign regs_60_io_reset = reset; // @[RegFile.scala 78:19:@50582.4]
  assign regs_60_io_enable = 1'h1; // @[RegFile.scala 74:20:@50576.4]
  assign regs_61_clock = clock; // @[:@50585.4]
  assign regs_61_reset = io_reset; // @[:@50586.4 RegFile.scala 76:16:@50593.4]
  assign regs_61_io_in = 64'h0; // @[RegFile.scala 75:16:@50592.4]
  assign regs_61_io_reset = reset; // @[RegFile.scala 78:19:@50596.4]
  assign regs_61_io_enable = 1'h1; // @[RegFile.scala 74:20:@50590.4]
  assign regs_62_clock = clock; // @[:@50599.4]
  assign regs_62_reset = io_reset; // @[:@50600.4 RegFile.scala 76:16:@50607.4]
  assign regs_62_io_in = 64'h0; // @[RegFile.scala 75:16:@50606.4]
  assign regs_62_io_reset = reset; // @[RegFile.scala 78:19:@50610.4]
  assign regs_62_io_enable = 1'h1; // @[RegFile.scala 74:20:@50604.4]
  assign regs_63_clock = clock; // @[:@50613.4]
  assign regs_63_reset = io_reset; // @[:@50614.4 RegFile.scala 76:16:@50621.4]
  assign regs_63_io_in = 64'h0; // @[RegFile.scala 75:16:@50620.4]
  assign regs_63_io_reset = reset; // @[RegFile.scala 78:19:@50624.4]
  assign regs_63_io_enable = 1'h1; // @[RegFile.scala 74:20:@50618.4]
  assign regs_64_clock = clock; // @[:@50627.4]
  assign regs_64_reset = io_reset; // @[:@50628.4 RegFile.scala 76:16:@50635.4]
  assign regs_64_io_in = 64'h0; // @[RegFile.scala 75:16:@50634.4]
  assign regs_64_io_reset = reset; // @[RegFile.scala 78:19:@50638.4]
  assign regs_64_io_enable = 1'h1; // @[RegFile.scala 74:20:@50632.4]
  assign regs_65_clock = clock; // @[:@50641.4]
  assign regs_65_reset = io_reset; // @[:@50642.4 RegFile.scala 76:16:@50649.4]
  assign regs_65_io_in = 64'h0; // @[RegFile.scala 75:16:@50648.4]
  assign regs_65_io_reset = reset; // @[RegFile.scala 78:19:@50652.4]
  assign regs_65_io_enable = 1'h1; // @[RegFile.scala 74:20:@50646.4]
  assign regs_66_clock = clock; // @[:@50655.4]
  assign regs_66_reset = io_reset; // @[:@50656.4 RegFile.scala 76:16:@50663.4]
  assign regs_66_io_in = 64'h0; // @[RegFile.scala 75:16:@50662.4]
  assign regs_66_io_reset = reset; // @[RegFile.scala 78:19:@50666.4]
  assign regs_66_io_enable = 1'h1; // @[RegFile.scala 74:20:@50660.4]
  assign regs_67_clock = clock; // @[:@50669.4]
  assign regs_67_reset = io_reset; // @[:@50670.4 RegFile.scala 76:16:@50677.4]
  assign regs_67_io_in = 64'h0; // @[RegFile.scala 75:16:@50676.4]
  assign regs_67_io_reset = reset; // @[RegFile.scala 78:19:@50680.4]
  assign regs_67_io_enable = 1'h1; // @[RegFile.scala 74:20:@50674.4]
  assign regs_68_clock = clock; // @[:@50683.4]
  assign regs_68_reset = io_reset; // @[:@50684.4 RegFile.scala 76:16:@50691.4]
  assign regs_68_io_in = 64'h0; // @[RegFile.scala 75:16:@50690.4]
  assign regs_68_io_reset = reset; // @[RegFile.scala 78:19:@50694.4]
  assign regs_68_io_enable = 1'h1; // @[RegFile.scala 74:20:@50688.4]
  assign regs_69_clock = clock; // @[:@50697.4]
  assign regs_69_reset = io_reset; // @[:@50698.4 RegFile.scala 76:16:@50705.4]
  assign regs_69_io_in = 64'h0; // @[RegFile.scala 75:16:@50704.4]
  assign regs_69_io_reset = reset; // @[RegFile.scala 78:19:@50708.4]
  assign regs_69_io_enable = 1'h1; // @[RegFile.scala 74:20:@50702.4]
  assign regs_70_clock = clock; // @[:@50711.4]
  assign regs_70_reset = io_reset; // @[:@50712.4 RegFile.scala 76:16:@50719.4]
  assign regs_70_io_in = 64'h0; // @[RegFile.scala 75:16:@50718.4]
  assign regs_70_io_reset = reset; // @[RegFile.scala 78:19:@50722.4]
  assign regs_70_io_enable = 1'h1; // @[RegFile.scala 74:20:@50716.4]
  assign regs_71_clock = clock; // @[:@50725.4]
  assign regs_71_reset = io_reset; // @[:@50726.4 RegFile.scala 76:16:@50733.4]
  assign regs_71_io_in = 64'h0; // @[RegFile.scala 75:16:@50732.4]
  assign regs_71_io_reset = reset; // @[RegFile.scala 78:19:@50736.4]
  assign regs_71_io_enable = 1'h1; // @[RegFile.scala 74:20:@50730.4]
  assign regs_72_clock = clock; // @[:@50739.4]
  assign regs_72_reset = io_reset; // @[:@50740.4 RegFile.scala 76:16:@50747.4]
  assign regs_72_io_in = 64'h0; // @[RegFile.scala 75:16:@50746.4]
  assign regs_72_io_reset = reset; // @[RegFile.scala 78:19:@50750.4]
  assign regs_72_io_enable = 1'h1; // @[RegFile.scala 74:20:@50744.4]
  assign regs_73_clock = clock; // @[:@50753.4]
  assign regs_73_reset = io_reset; // @[:@50754.4 RegFile.scala 76:16:@50761.4]
  assign regs_73_io_in = 64'h0; // @[RegFile.scala 75:16:@50760.4]
  assign regs_73_io_reset = reset; // @[RegFile.scala 78:19:@50764.4]
  assign regs_73_io_enable = 1'h1; // @[RegFile.scala 74:20:@50758.4]
  assign regs_74_clock = clock; // @[:@50767.4]
  assign regs_74_reset = io_reset; // @[:@50768.4 RegFile.scala 76:16:@50775.4]
  assign regs_74_io_in = 64'h0; // @[RegFile.scala 75:16:@50774.4]
  assign regs_74_io_reset = reset; // @[RegFile.scala 78:19:@50778.4]
  assign regs_74_io_enable = 1'h1; // @[RegFile.scala 74:20:@50772.4]
  assign regs_75_clock = clock; // @[:@50781.4]
  assign regs_75_reset = io_reset; // @[:@50782.4 RegFile.scala 76:16:@50789.4]
  assign regs_75_io_in = 64'h0; // @[RegFile.scala 75:16:@50788.4]
  assign regs_75_io_reset = reset; // @[RegFile.scala 78:19:@50792.4]
  assign regs_75_io_enable = 1'h1; // @[RegFile.scala 74:20:@50786.4]
  assign regs_76_clock = clock; // @[:@50795.4]
  assign regs_76_reset = io_reset; // @[:@50796.4 RegFile.scala 76:16:@50803.4]
  assign regs_76_io_in = 64'h0; // @[RegFile.scala 75:16:@50802.4]
  assign regs_76_io_reset = reset; // @[RegFile.scala 78:19:@50806.4]
  assign regs_76_io_enable = 1'h1; // @[RegFile.scala 74:20:@50800.4]
  assign regs_77_clock = clock; // @[:@50809.4]
  assign regs_77_reset = io_reset; // @[:@50810.4 RegFile.scala 76:16:@50817.4]
  assign regs_77_io_in = 64'h0; // @[RegFile.scala 75:16:@50816.4]
  assign regs_77_io_reset = reset; // @[RegFile.scala 78:19:@50820.4]
  assign regs_77_io_enable = 1'h1; // @[RegFile.scala 74:20:@50814.4]
  assign regs_78_clock = clock; // @[:@50823.4]
  assign regs_78_reset = io_reset; // @[:@50824.4 RegFile.scala 76:16:@50831.4]
  assign regs_78_io_in = 64'h0; // @[RegFile.scala 75:16:@50830.4]
  assign regs_78_io_reset = reset; // @[RegFile.scala 78:19:@50834.4]
  assign regs_78_io_enable = 1'h1; // @[RegFile.scala 74:20:@50828.4]
  assign regs_79_clock = clock; // @[:@50837.4]
  assign regs_79_reset = io_reset; // @[:@50838.4 RegFile.scala 76:16:@50845.4]
  assign regs_79_io_in = 64'h0; // @[RegFile.scala 75:16:@50844.4]
  assign regs_79_io_reset = reset; // @[RegFile.scala 78:19:@50848.4]
  assign regs_79_io_enable = 1'h1; // @[RegFile.scala 74:20:@50842.4]
  assign regs_80_clock = clock; // @[:@50851.4]
  assign regs_80_reset = io_reset; // @[:@50852.4 RegFile.scala 76:16:@50859.4]
  assign regs_80_io_in = 64'h0; // @[RegFile.scala 75:16:@50858.4]
  assign regs_80_io_reset = reset; // @[RegFile.scala 78:19:@50862.4]
  assign regs_80_io_enable = 1'h1; // @[RegFile.scala 74:20:@50856.4]
  assign regs_81_clock = clock; // @[:@50865.4]
  assign regs_81_reset = io_reset; // @[:@50866.4 RegFile.scala 76:16:@50873.4]
  assign regs_81_io_in = 64'h0; // @[RegFile.scala 75:16:@50872.4]
  assign regs_81_io_reset = reset; // @[RegFile.scala 78:19:@50876.4]
  assign regs_81_io_enable = 1'h1; // @[RegFile.scala 74:20:@50870.4]
  assign regs_82_clock = clock; // @[:@50879.4]
  assign regs_82_reset = io_reset; // @[:@50880.4 RegFile.scala 76:16:@50887.4]
  assign regs_82_io_in = 64'h0; // @[RegFile.scala 75:16:@50886.4]
  assign regs_82_io_reset = reset; // @[RegFile.scala 78:19:@50890.4]
  assign regs_82_io_enable = 1'h1; // @[RegFile.scala 74:20:@50884.4]
  assign regs_83_clock = clock; // @[:@50893.4]
  assign regs_83_reset = io_reset; // @[:@50894.4 RegFile.scala 76:16:@50901.4]
  assign regs_83_io_in = 64'h0; // @[RegFile.scala 75:16:@50900.4]
  assign regs_83_io_reset = reset; // @[RegFile.scala 78:19:@50904.4]
  assign regs_83_io_enable = 1'h1; // @[RegFile.scala 74:20:@50898.4]
  assign regs_84_clock = clock; // @[:@50907.4]
  assign regs_84_reset = io_reset; // @[:@50908.4 RegFile.scala 76:16:@50915.4]
  assign regs_84_io_in = 64'h0; // @[RegFile.scala 75:16:@50914.4]
  assign regs_84_io_reset = reset; // @[RegFile.scala 78:19:@50918.4]
  assign regs_84_io_enable = 1'h1; // @[RegFile.scala 74:20:@50912.4]
  assign regs_85_clock = clock; // @[:@50921.4]
  assign regs_85_reset = io_reset; // @[:@50922.4 RegFile.scala 76:16:@50929.4]
  assign regs_85_io_in = 64'h0; // @[RegFile.scala 75:16:@50928.4]
  assign regs_85_io_reset = reset; // @[RegFile.scala 78:19:@50932.4]
  assign regs_85_io_enable = 1'h1; // @[RegFile.scala 74:20:@50926.4]
  assign regs_86_clock = clock; // @[:@50935.4]
  assign regs_86_reset = io_reset; // @[:@50936.4 RegFile.scala 76:16:@50943.4]
  assign regs_86_io_in = 64'h0; // @[RegFile.scala 75:16:@50942.4]
  assign regs_86_io_reset = reset; // @[RegFile.scala 78:19:@50946.4]
  assign regs_86_io_enable = 1'h1; // @[RegFile.scala 74:20:@50940.4]
  assign regs_87_clock = clock; // @[:@50949.4]
  assign regs_87_reset = io_reset; // @[:@50950.4 RegFile.scala 76:16:@50957.4]
  assign regs_87_io_in = 64'h0; // @[RegFile.scala 75:16:@50956.4]
  assign regs_87_io_reset = reset; // @[RegFile.scala 78:19:@50960.4]
  assign regs_87_io_enable = 1'h1; // @[RegFile.scala 74:20:@50954.4]
  assign regs_88_clock = clock; // @[:@50963.4]
  assign regs_88_reset = io_reset; // @[:@50964.4 RegFile.scala 76:16:@50971.4]
  assign regs_88_io_in = 64'h0; // @[RegFile.scala 75:16:@50970.4]
  assign regs_88_io_reset = reset; // @[RegFile.scala 78:19:@50974.4]
  assign regs_88_io_enable = 1'h1; // @[RegFile.scala 74:20:@50968.4]
  assign regs_89_clock = clock; // @[:@50977.4]
  assign regs_89_reset = io_reset; // @[:@50978.4 RegFile.scala 76:16:@50985.4]
  assign regs_89_io_in = 64'h0; // @[RegFile.scala 75:16:@50984.4]
  assign regs_89_io_reset = reset; // @[RegFile.scala 78:19:@50988.4]
  assign regs_89_io_enable = 1'h1; // @[RegFile.scala 74:20:@50982.4]
  assign regs_90_clock = clock; // @[:@50991.4]
  assign regs_90_reset = io_reset; // @[:@50992.4 RegFile.scala 76:16:@50999.4]
  assign regs_90_io_in = 64'h0; // @[RegFile.scala 75:16:@50998.4]
  assign regs_90_io_reset = reset; // @[RegFile.scala 78:19:@51002.4]
  assign regs_90_io_enable = 1'h1; // @[RegFile.scala 74:20:@50996.4]
  assign regs_91_clock = clock; // @[:@51005.4]
  assign regs_91_reset = io_reset; // @[:@51006.4 RegFile.scala 76:16:@51013.4]
  assign regs_91_io_in = 64'h0; // @[RegFile.scala 75:16:@51012.4]
  assign regs_91_io_reset = reset; // @[RegFile.scala 78:19:@51016.4]
  assign regs_91_io_enable = 1'h1; // @[RegFile.scala 74:20:@51010.4]
  assign regs_92_clock = clock; // @[:@51019.4]
  assign regs_92_reset = io_reset; // @[:@51020.4 RegFile.scala 76:16:@51027.4]
  assign regs_92_io_in = 64'h0; // @[RegFile.scala 75:16:@51026.4]
  assign regs_92_io_reset = reset; // @[RegFile.scala 78:19:@51030.4]
  assign regs_92_io_enable = 1'h1; // @[RegFile.scala 74:20:@51024.4]
  assign regs_93_clock = clock; // @[:@51033.4]
  assign regs_93_reset = io_reset; // @[:@51034.4 RegFile.scala 76:16:@51041.4]
  assign regs_93_io_in = 64'h0; // @[RegFile.scala 75:16:@51040.4]
  assign regs_93_io_reset = reset; // @[RegFile.scala 78:19:@51044.4]
  assign regs_93_io_enable = 1'h1; // @[RegFile.scala 74:20:@51038.4]
  assign regs_94_clock = clock; // @[:@51047.4]
  assign regs_94_reset = io_reset; // @[:@51048.4 RegFile.scala 76:16:@51055.4]
  assign regs_94_io_in = 64'h0; // @[RegFile.scala 75:16:@51054.4]
  assign regs_94_io_reset = reset; // @[RegFile.scala 78:19:@51058.4]
  assign regs_94_io_enable = 1'h1; // @[RegFile.scala 74:20:@51052.4]
  assign regs_95_clock = clock; // @[:@51061.4]
  assign regs_95_reset = io_reset; // @[:@51062.4 RegFile.scala 76:16:@51069.4]
  assign regs_95_io_in = 64'h0; // @[RegFile.scala 75:16:@51068.4]
  assign regs_95_io_reset = reset; // @[RegFile.scala 78:19:@51072.4]
  assign regs_95_io_enable = 1'h1; // @[RegFile.scala 74:20:@51066.4]
  assign regs_96_clock = clock; // @[:@51075.4]
  assign regs_96_reset = io_reset; // @[:@51076.4 RegFile.scala 76:16:@51083.4]
  assign regs_96_io_in = 64'h0; // @[RegFile.scala 75:16:@51082.4]
  assign regs_96_io_reset = reset; // @[RegFile.scala 78:19:@51086.4]
  assign regs_96_io_enable = 1'h1; // @[RegFile.scala 74:20:@51080.4]
  assign regs_97_clock = clock; // @[:@51089.4]
  assign regs_97_reset = io_reset; // @[:@51090.4 RegFile.scala 76:16:@51097.4]
  assign regs_97_io_in = 64'h0; // @[RegFile.scala 75:16:@51096.4]
  assign regs_97_io_reset = reset; // @[RegFile.scala 78:19:@51100.4]
  assign regs_97_io_enable = 1'h1; // @[RegFile.scala 74:20:@51094.4]
  assign regs_98_clock = clock; // @[:@51103.4]
  assign regs_98_reset = io_reset; // @[:@51104.4 RegFile.scala 76:16:@51111.4]
  assign regs_98_io_in = 64'h0; // @[RegFile.scala 75:16:@51110.4]
  assign regs_98_io_reset = reset; // @[RegFile.scala 78:19:@51114.4]
  assign regs_98_io_enable = 1'h1; // @[RegFile.scala 74:20:@51108.4]
  assign regs_99_clock = clock; // @[:@51117.4]
  assign regs_99_reset = io_reset; // @[:@51118.4 RegFile.scala 76:16:@51125.4]
  assign regs_99_io_in = 64'h0; // @[RegFile.scala 75:16:@51124.4]
  assign regs_99_io_reset = reset; // @[RegFile.scala 78:19:@51128.4]
  assign regs_99_io_enable = 1'h1; // @[RegFile.scala 74:20:@51122.4]
  assign regs_100_clock = clock; // @[:@51131.4]
  assign regs_100_reset = io_reset; // @[:@51132.4 RegFile.scala 76:16:@51139.4]
  assign regs_100_io_in = 64'h0; // @[RegFile.scala 75:16:@51138.4]
  assign regs_100_io_reset = reset; // @[RegFile.scala 78:19:@51142.4]
  assign regs_100_io_enable = 1'h1; // @[RegFile.scala 74:20:@51136.4]
  assign regs_101_clock = clock; // @[:@51145.4]
  assign regs_101_reset = io_reset; // @[:@51146.4 RegFile.scala 76:16:@51153.4]
  assign regs_101_io_in = 64'h0; // @[RegFile.scala 75:16:@51152.4]
  assign regs_101_io_reset = reset; // @[RegFile.scala 78:19:@51156.4]
  assign regs_101_io_enable = 1'h1; // @[RegFile.scala 74:20:@51150.4]
  assign regs_102_clock = clock; // @[:@51159.4]
  assign regs_102_reset = io_reset; // @[:@51160.4 RegFile.scala 76:16:@51167.4]
  assign regs_102_io_in = 64'h0; // @[RegFile.scala 75:16:@51166.4]
  assign regs_102_io_reset = reset; // @[RegFile.scala 78:19:@51170.4]
  assign regs_102_io_enable = 1'h1; // @[RegFile.scala 74:20:@51164.4]
  assign regs_103_clock = clock; // @[:@51173.4]
  assign regs_103_reset = io_reset; // @[:@51174.4 RegFile.scala 76:16:@51181.4]
  assign regs_103_io_in = 64'h0; // @[RegFile.scala 75:16:@51180.4]
  assign regs_103_io_reset = reset; // @[RegFile.scala 78:19:@51184.4]
  assign regs_103_io_enable = 1'h1; // @[RegFile.scala 74:20:@51178.4]
  assign regs_104_clock = clock; // @[:@51187.4]
  assign regs_104_reset = io_reset; // @[:@51188.4 RegFile.scala 76:16:@51195.4]
  assign regs_104_io_in = 64'h0; // @[RegFile.scala 75:16:@51194.4]
  assign regs_104_io_reset = reset; // @[RegFile.scala 78:19:@51198.4]
  assign regs_104_io_enable = 1'h1; // @[RegFile.scala 74:20:@51192.4]
  assign regs_105_clock = clock; // @[:@51201.4]
  assign regs_105_reset = io_reset; // @[:@51202.4 RegFile.scala 76:16:@51209.4]
  assign regs_105_io_in = 64'h0; // @[RegFile.scala 75:16:@51208.4]
  assign regs_105_io_reset = reset; // @[RegFile.scala 78:19:@51212.4]
  assign regs_105_io_enable = 1'h1; // @[RegFile.scala 74:20:@51206.4]
  assign regs_106_clock = clock; // @[:@51215.4]
  assign regs_106_reset = io_reset; // @[:@51216.4 RegFile.scala 76:16:@51223.4]
  assign regs_106_io_in = 64'h0; // @[RegFile.scala 75:16:@51222.4]
  assign regs_106_io_reset = reset; // @[RegFile.scala 78:19:@51226.4]
  assign regs_106_io_enable = 1'h1; // @[RegFile.scala 74:20:@51220.4]
  assign regs_107_clock = clock; // @[:@51229.4]
  assign regs_107_reset = io_reset; // @[:@51230.4 RegFile.scala 76:16:@51237.4]
  assign regs_107_io_in = 64'h0; // @[RegFile.scala 75:16:@51236.4]
  assign regs_107_io_reset = reset; // @[RegFile.scala 78:19:@51240.4]
  assign regs_107_io_enable = 1'h1; // @[RegFile.scala 74:20:@51234.4]
  assign regs_108_clock = clock; // @[:@51243.4]
  assign regs_108_reset = io_reset; // @[:@51244.4 RegFile.scala 76:16:@51251.4]
  assign regs_108_io_in = 64'h0; // @[RegFile.scala 75:16:@51250.4]
  assign regs_108_io_reset = reset; // @[RegFile.scala 78:19:@51254.4]
  assign regs_108_io_enable = 1'h1; // @[RegFile.scala 74:20:@51248.4]
  assign regs_109_clock = clock; // @[:@51257.4]
  assign regs_109_reset = io_reset; // @[:@51258.4 RegFile.scala 76:16:@51265.4]
  assign regs_109_io_in = 64'h0; // @[RegFile.scala 75:16:@51264.4]
  assign regs_109_io_reset = reset; // @[RegFile.scala 78:19:@51268.4]
  assign regs_109_io_enable = 1'h1; // @[RegFile.scala 74:20:@51262.4]
  assign regs_110_clock = clock; // @[:@51271.4]
  assign regs_110_reset = io_reset; // @[:@51272.4 RegFile.scala 76:16:@51279.4]
  assign regs_110_io_in = 64'h0; // @[RegFile.scala 75:16:@51278.4]
  assign regs_110_io_reset = reset; // @[RegFile.scala 78:19:@51282.4]
  assign regs_110_io_enable = 1'h1; // @[RegFile.scala 74:20:@51276.4]
  assign regs_111_clock = clock; // @[:@51285.4]
  assign regs_111_reset = io_reset; // @[:@51286.4 RegFile.scala 76:16:@51293.4]
  assign regs_111_io_in = 64'h0; // @[RegFile.scala 75:16:@51292.4]
  assign regs_111_io_reset = reset; // @[RegFile.scala 78:19:@51296.4]
  assign regs_111_io_enable = 1'h1; // @[RegFile.scala 74:20:@51290.4]
  assign regs_112_clock = clock; // @[:@51299.4]
  assign regs_112_reset = io_reset; // @[:@51300.4 RegFile.scala 76:16:@51307.4]
  assign regs_112_io_in = 64'h0; // @[RegFile.scala 75:16:@51306.4]
  assign regs_112_io_reset = reset; // @[RegFile.scala 78:19:@51310.4]
  assign regs_112_io_enable = 1'h1; // @[RegFile.scala 74:20:@51304.4]
  assign regs_113_clock = clock; // @[:@51313.4]
  assign regs_113_reset = io_reset; // @[:@51314.4 RegFile.scala 76:16:@51321.4]
  assign regs_113_io_in = 64'h0; // @[RegFile.scala 75:16:@51320.4]
  assign regs_113_io_reset = reset; // @[RegFile.scala 78:19:@51324.4]
  assign regs_113_io_enable = 1'h1; // @[RegFile.scala 74:20:@51318.4]
  assign regs_114_clock = clock; // @[:@51327.4]
  assign regs_114_reset = io_reset; // @[:@51328.4 RegFile.scala 76:16:@51335.4]
  assign regs_114_io_in = 64'h0; // @[RegFile.scala 75:16:@51334.4]
  assign regs_114_io_reset = reset; // @[RegFile.scala 78:19:@51338.4]
  assign regs_114_io_enable = 1'h1; // @[RegFile.scala 74:20:@51332.4]
  assign regs_115_clock = clock; // @[:@51341.4]
  assign regs_115_reset = io_reset; // @[:@51342.4 RegFile.scala 76:16:@51349.4]
  assign regs_115_io_in = 64'h0; // @[RegFile.scala 75:16:@51348.4]
  assign regs_115_io_reset = reset; // @[RegFile.scala 78:19:@51352.4]
  assign regs_115_io_enable = 1'h1; // @[RegFile.scala 74:20:@51346.4]
  assign regs_116_clock = clock; // @[:@51355.4]
  assign regs_116_reset = io_reset; // @[:@51356.4 RegFile.scala 76:16:@51363.4]
  assign regs_116_io_in = 64'h0; // @[RegFile.scala 75:16:@51362.4]
  assign regs_116_io_reset = reset; // @[RegFile.scala 78:19:@51366.4]
  assign regs_116_io_enable = 1'h1; // @[RegFile.scala 74:20:@51360.4]
  assign regs_117_clock = clock; // @[:@51369.4]
  assign regs_117_reset = io_reset; // @[:@51370.4 RegFile.scala 76:16:@51377.4]
  assign regs_117_io_in = 64'h0; // @[RegFile.scala 75:16:@51376.4]
  assign regs_117_io_reset = reset; // @[RegFile.scala 78:19:@51380.4]
  assign regs_117_io_enable = 1'h1; // @[RegFile.scala 74:20:@51374.4]
  assign regs_118_clock = clock; // @[:@51383.4]
  assign regs_118_reset = io_reset; // @[:@51384.4 RegFile.scala 76:16:@51391.4]
  assign regs_118_io_in = 64'h0; // @[RegFile.scala 75:16:@51390.4]
  assign regs_118_io_reset = reset; // @[RegFile.scala 78:19:@51394.4]
  assign regs_118_io_enable = 1'h1; // @[RegFile.scala 74:20:@51388.4]
  assign regs_119_clock = clock; // @[:@51397.4]
  assign regs_119_reset = io_reset; // @[:@51398.4 RegFile.scala 76:16:@51405.4]
  assign regs_119_io_in = 64'h0; // @[RegFile.scala 75:16:@51404.4]
  assign regs_119_io_reset = reset; // @[RegFile.scala 78:19:@51408.4]
  assign regs_119_io_enable = 1'h1; // @[RegFile.scala 74:20:@51402.4]
  assign regs_120_clock = clock; // @[:@51411.4]
  assign regs_120_reset = io_reset; // @[:@51412.4 RegFile.scala 76:16:@51419.4]
  assign regs_120_io_in = 64'h0; // @[RegFile.scala 75:16:@51418.4]
  assign regs_120_io_reset = reset; // @[RegFile.scala 78:19:@51422.4]
  assign regs_120_io_enable = 1'h1; // @[RegFile.scala 74:20:@51416.4]
  assign regs_121_clock = clock; // @[:@51425.4]
  assign regs_121_reset = io_reset; // @[:@51426.4 RegFile.scala 76:16:@51433.4]
  assign regs_121_io_in = 64'h0; // @[RegFile.scala 75:16:@51432.4]
  assign regs_121_io_reset = reset; // @[RegFile.scala 78:19:@51436.4]
  assign regs_121_io_enable = 1'h1; // @[RegFile.scala 74:20:@51430.4]
  assign regs_122_clock = clock; // @[:@51439.4]
  assign regs_122_reset = io_reset; // @[:@51440.4 RegFile.scala 76:16:@51447.4]
  assign regs_122_io_in = 64'h0; // @[RegFile.scala 75:16:@51446.4]
  assign regs_122_io_reset = reset; // @[RegFile.scala 78:19:@51450.4]
  assign regs_122_io_enable = 1'h1; // @[RegFile.scala 74:20:@51444.4]
  assign regs_123_clock = clock; // @[:@51453.4]
  assign regs_123_reset = io_reset; // @[:@51454.4 RegFile.scala 76:16:@51461.4]
  assign regs_123_io_in = 64'h0; // @[RegFile.scala 75:16:@51460.4]
  assign regs_123_io_reset = reset; // @[RegFile.scala 78:19:@51464.4]
  assign regs_123_io_enable = 1'h1; // @[RegFile.scala 74:20:@51458.4]
  assign regs_124_clock = clock; // @[:@51467.4]
  assign regs_124_reset = io_reset; // @[:@51468.4 RegFile.scala 76:16:@51475.4]
  assign regs_124_io_in = 64'h0; // @[RegFile.scala 75:16:@51474.4]
  assign regs_124_io_reset = reset; // @[RegFile.scala 78:19:@51478.4]
  assign regs_124_io_enable = 1'h1; // @[RegFile.scala 74:20:@51472.4]
  assign regs_125_clock = clock; // @[:@51481.4]
  assign regs_125_reset = io_reset; // @[:@51482.4 RegFile.scala 76:16:@51489.4]
  assign regs_125_io_in = 64'h0; // @[RegFile.scala 75:16:@51488.4]
  assign regs_125_io_reset = reset; // @[RegFile.scala 78:19:@51492.4]
  assign regs_125_io_enable = 1'h1; // @[RegFile.scala 74:20:@51486.4]
  assign regs_126_clock = clock; // @[:@51495.4]
  assign regs_126_reset = io_reset; // @[:@51496.4 RegFile.scala 76:16:@51503.4]
  assign regs_126_io_in = 64'h0; // @[RegFile.scala 75:16:@51502.4]
  assign regs_126_io_reset = reset; // @[RegFile.scala 78:19:@51506.4]
  assign regs_126_io_enable = 1'h1; // @[RegFile.scala 74:20:@51500.4]
  assign regs_127_clock = clock; // @[:@51509.4]
  assign regs_127_reset = io_reset; // @[:@51510.4 RegFile.scala 76:16:@51517.4]
  assign regs_127_io_in = 64'h0; // @[RegFile.scala 75:16:@51516.4]
  assign regs_127_io_reset = reset; // @[RegFile.scala 78:19:@51520.4]
  assign regs_127_io_enable = 1'h1; // @[RegFile.scala 74:20:@51514.4]
  assign regs_128_clock = clock; // @[:@51523.4]
  assign regs_128_reset = io_reset; // @[:@51524.4 RegFile.scala 76:16:@51531.4]
  assign regs_128_io_in = 64'h0; // @[RegFile.scala 75:16:@51530.4]
  assign regs_128_io_reset = reset; // @[RegFile.scala 78:19:@51534.4]
  assign regs_128_io_enable = 1'h1; // @[RegFile.scala 74:20:@51528.4]
  assign regs_129_clock = clock; // @[:@51537.4]
  assign regs_129_reset = io_reset; // @[:@51538.4 RegFile.scala 76:16:@51545.4]
  assign regs_129_io_in = 64'h0; // @[RegFile.scala 75:16:@51544.4]
  assign regs_129_io_reset = reset; // @[RegFile.scala 78:19:@51548.4]
  assign regs_129_io_enable = 1'h1; // @[RegFile.scala 74:20:@51542.4]
  assign regs_130_clock = clock; // @[:@51551.4]
  assign regs_130_reset = io_reset; // @[:@51552.4 RegFile.scala 76:16:@51559.4]
  assign regs_130_io_in = 64'h0; // @[RegFile.scala 75:16:@51558.4]
  assign regs_130_io_reset = reset; // @[RegFile.scala 78:19:@51562.4]
  assign regs_130_io_enable = 1'h1; // @[RegFile.scala 74:20:@51556.4]
  assign regs_131_clock = clock; // @[:@51565.4]
  assign regs_131_reset = io_reset; // @[:@51566.4 RegFile.scala 76:16:@51573.4]
  assign regs_131_io_in = 64'h0; // @[RegFile.scala 75:16:@51572.4]
  assign regs_131_io_reset = reset; // @[RegFile.scala 78:19:@51576.4]
  assign regs_131_io_enable = 1'h1; // @[RegFile.scala 74:20:@51570.4]
  assign regs_132_clock = clock; // @[:@51579.4]
  assign regs_132_reset = io_reset; // @[:@51580.4 RegFile.scala 76:16:@51587.4]
  assign regs_132_io_in = 64'h0; // @[RegFile.scala 75:16:@51586.4]
  assign regs_132_io_reset = reset; // @[RegFile.scala 78:19:@51590.4]
  assign regs_132_io_enable = 1'h1; // @[RegFile.scala 74:20:@51584.4]
  assign regs_133_clock = clock; // @[:@51593.4]
  assign regs_133_reset = io_reset; // @[:@51594.4 RegFile.scala 76:16:@51601.4]
  assign regs_133_io_in = 64'h0; // @[RegFile.scala 75:16:@51600.4]
  assign regs_133_io_reset = reset; // @[RegFile.scala 78:19:@51604.4]
  assign regs_133_io_enable = 1'h1; // @[RegFile.scala 74:20:@51598.4]
  assign regs_134_clock = clock; // @[:@51607.4]
  assign regs_134_reset = io_reset; // @[:@51608.4 RegFile.scala 76:16:@51615.4]
  assign regs_134_io_in = 64'h0; // @[RegFile.scala 75:16:@51614.4]
  assign regs_134_io_reset = reset; // @[RegFile.scala 78:19:@51618.4]
  assign regs_134_io_enable = 1'h1; // @[RegFile.scala 74:20:@51612.4]
  assign regs_135_clock = clock; // @[:@51621.4]
  assign regs_135_reset = io_reset; // @[:@51622.4 RegFile.scala 76:16:@51629.4]
  assign regs_135_io_in = 64'h0; // @[RegFile.scala 75:16:@51628.4]
  assign regs_135_io_reset = reset; // @[RegFile.scala 78:19:@51632.4]
  assign regs_135_io_enable = 1'h1; // @[RegFile.scala 74:20:@51626.4]
  assign regs_136_clock = clock; // @[:@51635.4]
  assign regs_136_reset = io_reset; // @[:@51636.4 RegFile.scala 76:16:@51643.4]
  assign regs_136_io_in = 64'h0; // @[RegFile.scala 75:16:@51642.4]
  assign regs_136_io_reset = reset; // @[RegFile.scala 78:19:@51646.4]
  assign regs_136_io_enable = 1'h1; // @[RegFile.scala 74:20:@51640.4]
  assign regs_137_clock = clock; // @[:@51649.4]
  assign regs_137_reset = io_reset; // @[:@51650.4 RegFile.scala 76:16:@51657.4]
  assign regs_137_io_in = 64'h0; // @[RegFile.scala 75:16:@51656.4]
  assign regs_137_io_reset = reset; // @[RegFile.scala 78:19:@51660.4]
  assign regs_137_io_enable = 1'h1; // @[RegFile.scala 74:20:@51654.4]
  assign regs_138_clock = clock; // @[:@51663.4]
  assign regs_138_reset = io_reset; // @[:@51664.4 RegFile.scala 76:16:@51671.4]
  assign regs_138_io_in = 64'h0; // @[RegFile.scala 75:16:@51670.4]
  assign regs_138_io_reset = reset; // @[RegFile.scala 78:19:@51674.4]
  assign regs_138_io_enable = 1'h1; // @[RegFile.scala 74:20:@51668.4]
  assign regs_139_clock = clock; // @[:@51677.4]
  assign regs_139_reset = io_reset; // @[:@51678.4 RegFile.scala 76:16:@51685.4]
  assign regs_139_io_in = 64'h0; // @[RegFile.scala 75:16:@51684.4]
  assign regs_139_io_reset = reset; // @[RegFile.scala 78:19:@51688.4]
  assign regs_139_io_enable = 1'h1; // @[RegFile.scala 74:20:@51682.4]
  assign regs_140_clock = clock; // @[:@51691.4]
  assign regs_140_reset = io_reset; // @[:@51692.4 RegFile.scala 76:16:@51699.4]
  assign regs_140_io_in = 64'h0; // @[RegFile.scala 75:16:@51698.4]
  assign regs_140_io_reset = reset; // @[RegFile.scala 78:19:@51702.4]
  assign regs_140_io_enable = 1'h1; // @[RegFile.scala 74:20:@51696.4]
  assign regs_141_clock = clock; // @[:@51705.4]
  assign regs_141_reset = io_reset; // @[:@51706.4 RegFile.scala 76:16:@51713.4]
  assign regs_141_io_in = 64'h0; // @[RegFile.scala 75:16:@51712.4]
  assign regs_141_io_reset = reset; // @[RegFile.scala 78:19:@51716.4]
  assign regs_141_io_enable = 1'h1; // @[RegFile.scala 74:20:@51710.4]
  assign regs_142_clock = clock; // @[:@51719.4]
  assign regs_142_reset = io_reset; // @[:@51720.4 RegFile.scala 76:16:@51727.4]
  assign regs_142_io_in = 64'h0; // @[RegFile.scala 75:16:@51726.4]
  assign regs_142_io_reset = reset; // @[RegFile.scala 78:19:@51730.4]
  assign regs_142_io_enable = 1'h1; // @[RegFile.scala 74:20:@51724.4]
  assign regs_143_clock = clock; // @[:@51733.4]
  assign regs_143_reset = io_reset; // @[:@51734.4 RegFile.scala 76:16:@51741.4]
  assign regs_143_io_in = 64'h0; // @[RegFile.scala 75:16:@51740.4]
  assign regs_143_io_reset = reset; // @[RegFile.scala 78:19:@51744.4]
  assign regs_143_io_enable = 1'h1; // @[RegFile.scala 74:20:@51738.4]
  assign regs_144_clock = clock; // @[:@51747.4]
  assign regs_144_reset = io_reset; // @[:@51748.4 RegFile.scala 76:16:@51755.4]
  assign regs_144_io_in = 64'h0; // @[RegFile.scala 75:16:@51754.4]
  assign regs_144_io_reset = reset; // @[RegFile.scala 78:19:@51758.4]
  assign regs_144_io_enable = 1'h1; // @[RegFile.scala 74:20:@51752.4]
  assign regs_145_clock = clock; // @[:@51761.4]
  assign regs_145_reset = io_reset; // @[:@51762.4 RegFile.scala 76:16:@51769.4]
  assign regs_145_io_in = 64'h0; // @[RegFile.scala 75:16:@51768.4]
  assign regs_145_io_reset = reset; // @[RegFile.scala 78:19:@51772.4]
  assign regs_145_io_enable = 1'h1; // @[RegFile.scala 74:20:@51766.4]
  assign regs_146_clock = clock; // @[:@51775.4]
  assign regs_146_reset = io_reset; // @[:@51776.4 RegFile.scala 76:16:@51783.4]
  assign regs_146_io_in = 64'h0; // @[RegFile.scala 75:16:@51782.4]
  assign regs_146_io_reset = reset; // @[RegFile.scala 78:19:@51786.4]
  assign regs_146_io_enable = 1'h1; // @[RegFile.scala 74:20:@51780.4]
  assign regs_147_clock = clock; // @[:@51789.4]
  assign regs_147_reset = io_reset; // @[:@51790.4 RegFile.scala 76:16:@51797.4]
  assign regs_147_io_in = 64'h0; // @[RegFile.scala 75:16:@51796.4]
  assign regs_147_io_reset = reset; // @[RegFile.scala 78:19:@51800.4]
  assign regs_147_io_enable = 1'h1; // @[RegFile.scala 74:20:@51794.4]
  assign regs_148_clock = clock; // @[:@51803.4]
  assign regs_148_reset = io_reset; // @[:@51804.4 RegFile.scala 76:16:@51811.4]
  assign regs_148_io_in = 64'h0; // @[RegFile.scala 75:16:@51810.4]
  assign regs_148_io_reset = reset; // @[RegFile.scala 78:19:@51814.4]
  assign regs_148_io_enable = 1'h1; // @[RegFile.scala 74:20:@51808.4]
  assign regs_149_clock = clock; // @[:@51817.4]
  assign regs_149_reset = io_reset; // @[:@51818.4 RegFile.scala 76:16:@51825.4]
  assign regs_149_io_in = 64'h0; // @[RegFile.scala 75:16:@51824.4]
  assign regs_149_io_reset = reset; // @[RegFile.scala 78:19:@51828.4]
  assign regs_149_io_enable = 1'h1; // @[RegFile.scala 74:20:@51822.4]
  assign regs_150_clock = clock; // @[:@51831.4]
  assign regs_150_reset = io_reset; // @[:@51832.4 RegFile.scala 76:16:@51839.4]
  assign regs_150_io_in = 64'h0; // @[RegFile.scala 75:16:@51838.4]
  assign regs_150_io_reset = reset; // @[RegFile.scala 78:19:@51842.4]
  assign regs_150_io_enable = 1'h1; // @[RegFile.scala 74:20:@51836.4]
  assign regs_151_clock = clock; // @[:@51845.4]
  assign regs_151_reset = io_reset; // @[:@51846.4 RegFile.scala 76:16:@51853.4]
  assign regs_151_io_in = 64'h0; // @[RegFile.scala 75:16:@51852.4]
  assign regs_151_io_reset = reset; // @[RegFile.scala 78:19:@51856.4]
  assign regs_151_io_enable = 1'h1; // @[RegFile.scala 74:20:@51850.4]
  assign regs_152_clock = clock; // @[:@51859.4]
  assign regs_152_reset = io_reset; // @[:@51860.4 RegFile.scala 76:16:@51867.4]
  assign regs_152_io_in = 64'h0; // @[RegFile.scala 75:16:@51866.4]
  assign regs_152_io_reset = reset; // @[RegFile.scala 78:19:@51870.4]
  assign regs_152_io_enable = 1'h1; // @[RegFile.scala 74:20:@51864.4]
  assign regs_153_clock = clock; // @[:@51873.4]
  assign regs_153_reset = io_reset; // @[:@51874.4 RegFile.scala 76:16:@51881.4]
  assign regs_153_io_in = 64'h0; // @[RegFile.scala 75:16:@51880.4]
  assign regs_153_io_reset = reset; // @[RegFile.scala 78:19:@51884.4]
  assign regs_153_io_enable = 1'h1; // @[RegFile.scala 74:20:@51878.4]
  assign regs_154_clock = clock; // @[:@51887.4]
  assign regs_154_reset = io_reset; // @[:@51888.4 RegFile.scala 76:16:@51895.4]
  assign regs_154_io_in = 64'h0; // @[RegFile.scala 75:16:@51894.4]
  assign regs_154_io_reset = reset; // @[RegFile.scala 78:19:@51898.4]
  assign regs_154_io_enable = 1'h1; // @[RegFile.scala 74:20:@51892.4]
  assign regs_155_clock = clock; // @[:@51901.4]
  assign regs_155_reset = io_reset; // @[:@51902.4 RegFile.scala 76:16:@51909.4]
  assign regs_155_io_in = 64'h0; // @[RegFile.scala 75:16:@51908.4]
  assign regs_155_io_reset = reset; // @[RegFile.scala 78:19:@51912.4]
  assign regs_155_io_enable = 1'h1; // @[RegFile.scala 74:20:@51906.4]
  assign regs_156_clock = clock; // @[:@51915.4]
  assign regs_156_reset = io_reset; // @[:@51916.4 RegFile.scala 76:16:@51923.4]
  assign regs_156_io_in = 64'h0; // @[RegFile.scala 75:16:@51922.4]
  assign regs_156_io_reset = reset; // @[RegFile.scala 78:19:@51926.4]
  assign regs_156_io_enable = 1'h1; // @[RegFile.scala 74:20:@51920.4]
  assign regs_157_clock = clock; // @[:@51929.4]
  assign regs_157_reset = io_reset; // @[:@51930.4 RegFile.scala 76:16:@51937.4]
  assign regs_157_io_in = 64'h0; // @[RegFile.scala 75:16:@51936.4]
  assign regs_157_io_reset = reset; // @[RegFile.scala 78:19:@51940.4]
  assign regs_157_io_enable = 1'h1; // @[RegFile.scala 74:20:@51934.4]
  assign regs_158_clock = clock; // @[:@51943.4]
  assign regs_158_reset = io_reset; // @[:@51944.4 RegFile.scala 76:16:@51951.4]
  assign regs_158_io_in = 64'h0; // @[RegFile.scala 75:16:@51950.4]
  assign regs_158_io_reset = reset; // @[RegFile.scala 78:19:@51954.4]
  assign regs_158_io_enable = 1'h1; // @[RegFile.scala 74:20:@51948.4]
  assign regs_159_clock = clock; // @[:@51957.4]
  assign regs_159_reset = io_reset; // @[:@51958.4 RegFile.scala 76:16:@51965.4]
  assign regs_159_io_in = 64'h0; // @[RegFile.scala 75:16:@51964.4]
  assign regs_159_io_reset = reset; // @[RegFile.scala 78:19:@51968.4]
  assign regs_159_io_enable = 1'h1; // @[RegFile.scala 74:20:@51962.4]
  assign regs_160_clock = clock; // @[:@51971.4]
  assign regs_160_reset = io_reset; // @[:@51972.4 RegFile.scala 76:16:@51979.4]
  assign regs_160_io_in = 64'h0; // @[RegFile.scala 75:16:@51978.4]
  assign regs_160_io_reset = reset; // @[RegFile.scala 78:19:@51982.4]
  assign regs_160_io_enable = 1'h1; // @[RegFile.scala 74:20:@51976.4]
  assign regs_161_clock = clock; // @[:@51985.4]
  assign regs_161_reset = io_reset; // @[:@51986.4 RegFile.scala 76:16:@51993.4]
  assign regs_161_io_in = 64'h0; // @[RegFile.scala 75:16:@51992.4]
  assign regs_161_io_reset = reset; // @[RegFile.scala 78:19:@51996.4]
  assign regs_161_io_enable = 1'h1; // @[RegFile.scala 74:20:@51990.4]
  assign regs_162_clock = clock; // @[:@51999.4]
  assign regs_162_reset = io_reset; // @[:@52000.4 RegFile.scala 76:16:@52007.4]
  assign regs_162_io_in = 64'h0; // @[RegFile.scala 75:16:@52006.4]
  assign regs_162_io_reset = reset; // @[RegFile.scala 78:19:@52010.4]
  assign regs_162_io_enable = 1'h1; // @[RegFile.scala 74:20:@52004.4]
  assign regs_163_clock = clock; // @[:@52013.4]
  assign regs_163_reset = io_reset; // @[:@52014.4 RegFile.scala 76:16:@52021.4]
  assign regs_163_io_in = 64'h0; // @[RegFile.scala 75:16:@52020.4]
  assign regs_163_io_reset = reset; // @[RegFile.scala 78:19:@52024.4]
  assign regs_163_io_enable = 1'h1; // @[RegFile.scala 74:20:@52018.4]
  assign regs_164_clock = clock; // @[:@52027.4]
  assign regs_164_reset = io_reset; // @[:@52028.4 RegFile.scala 76:16:@52035.4]
  assign regs_164_io_in = 64'h0; // @[RegFile.scala 75:16:@52034.4]
  assign regs_164_io_reset = reset; // @[RegFile.scala 78:19:@52038.4]
  assign regs_164_io_enable = 1'h1; // @[RegFile.scala 74:20:@52032.4]
  assign regs_165_clock = clock; // @[:@52041.4]
  assign regs_165_reset = io_reset; // @[:@52042.4 RegFile.scala 76:16:@52049.4]
  assign regs_165_io_in = 64'h0; // @[RegFile.scala 75:16:@52048.4]
  assign regs_165_io_reset = reset; // @[RegFile.scala 78:19:@52052.4]
  assign regs_165_io_enable = 1'h1; // @[RegFile.scala 74:20:@52046.4]
  assign regs_166_clock = clock; // @[:@52055.4]
  assign regs_166_reset = io_reset; // @[:@52056.4 RegFile.scala 76:16:@52063.4]
  assign regs_166_io_in = 64'h0; // @[RegFile.scala 75:16:@52062.4]
  assign regs_166_io_reset = reset; // @[RegFile.scala 78:19:@52066.4]
  assign regs_166_io_enable = 1'h1; // @[RegFile.scala 74:20:@52060.4]
  assign regs_167_clock = clock; // @[:@52069.4]
  assign regs_167_reset = io_reset; // @[:@52070.4 RegFile.scala 76:16:@52077.4]
  assign regs_167_io_in = 64'h0; // @[RegFile.scala 75:16:@52076.4]
  assign regs_167_io_reset = reset; // @[RegFile.scala 78:19:@52080.4]
  assign regs_167_io_enable = 1'h1; // @[RegFile.scala 74:20:@52074.4]
  assign regs_168_clock = clock; // @[:@52083.4]
  assign regs_168_reset = io_reset; // @[:@52084.4 RegFile.scala 76:16:@52091.4]
  assign regs_168_io_in = 64'h0; // @[RegFile.scala 75:16:@52090.4]
  assign regs_168_io_reset = reset; // @[RegFile.scala 78:19:@52094.4]
  assign regs_168_io_enable = 1'h1; // @[RegFile.scala 74:20:@52088.4]
  assign regs_169_clock = clock; // @[:@52097.4]
  assign regs_169_reset = io_reset; // @[:@52098.4 RegFile.scala 76:16:@52105.4]
  assign regs_169_io_in = 64'h0; // @[RegFile.scala 75:16:@52104.4]
  assign regs_169_io_reset = reset; // @[RegFile.scala 78:19:@52108.4]
  assign regs_169_io_enable = 1'h1; // @[RegFile.scala 74:20:@52102.4]
  assign regs_170_clock = clock; // @[:@52111.4]
  assign regs_170_reset = io_reset; // @[:@52112.4 RegFile.scala 76:16:@52119.4]
  assign regs_170_io_in = 64'h0; // @[RegFile.scala 75:16:@52118.4]
  assign regs_170_io_reset = reset; // @[RegFile.scala 78:19:@52122.4]
  assign regs_170_io_enable = 1'h1; // @[RegFile.scala 74:20:@52116.4]
  assign regs_171_clock = clock; // @[:@52125.4]
  assign regs_171_reset = io_reset; // @[:@52126.4 RegFile.scala 76:16:@52133.4]
  assign regs_171_io_in = 64'h0; // @[RegFile.scala 75:16:@52132.4]
  assign regs_171_io_reset = reset; // @[RegFile.scala 78:19:@52136.4]
  assign regs_171_io_enable = 1'h1; // @[RegFile.scala 74:20:@52130.4]
  assign regs_172_clock = clock; // @[:@52139.4]
  assign regs_172_reset = io_reset; // @[:@52140.4 RegFile.scala 76:16:@52147.4]
  assign regs_172_io_in = 64'h0; // @[RegFile.scala 75:16:@52146.4]
  assign regs_172_io_reset = reset; // @[RegFile.scala 78:19:@52150.4]
  assign regs_172_io_enable = 1'h1; // @[RegFile.scala 74:20:@52144.4]
  assign regs_173_clock = clock; // @[:@52153.4]
  assign regs_173_reset = io_reset; // @[:@52154.4 RegFile.scala 76:16:@52161.4]
  assign regs_173_io_in = 64'h0; // @[RegFile.scala 75:16:@52160.4]
  assign regs_173_io_reset = reset; // @[RegFile.scala 78:19:@52164.4]
  assign regs_173_io_enable = 1'h1; // @[RegFile.scala 74:20:@52158.4]
  assign regs_174_clock = clock; // @[:@52167.4]
  assign regs_174_reset = io_reset; // @[:@52168.4 RegFile.scala 76:16:@52175.4]
  assign regs_174_io_in = 64'h0; // @[RegFile.scala 75:16:@52174.4]
  assign regs_174_io_reset = reset; // @[RegFile.scala 78:19:@52178.4]
  assign regs_174_io_enable = 1'h1; // @[RegFile.scala 74:20:@52172.4]
  assign regs_175_clock = clock; // @[:@52181.4]
  assign regs_175_reset = io_reset; // @[:@52182.4 RegFile.scala 76:16:@52189.4]
  assign regs_175_io_in = 64'h0; // @[RegFile.scala 75:16:@52188.4]
  assign regs_175_io_reset = reset; // @[RegFile.scala 78:19:@52192.4]
  assign regs_175_io_enable = 1'h1; // @[RegFile.scala 74:20:@52186.4]
  assign regs_176_clock = clock; // @[:@52195.4]
  assign regs_176_reset = io_reset; // @[:@52196.4 RegFile.scala 76:16:@52203.4]
  assign regs_176_io_in = 64'h0; // @[RegFile.scala 75:16:@52202.4]
  assign regs_176_io_reset = reset; // @[RegFile.scala 78:19:@52206.4]
  assign regs_176_io_enable = 1'h1; // @[RegFile.scala 74:20:@52200.4]
  assign regs_177_clock = clock; // @[:@52209.4]
  assign regs_177_reset = io_reset; // @[:@52210.4 RegFile.scala 76:16:@52217.4]
  assign regs_177_io_in = 64'h0; // @[RegFile.scala 75:16:@52216.4]
  assign regs_177_io_reset = reset; // @[RegFile.scala 78:19:@52220.4]
  assign regs_177_io_enable = 1'h1; // @[RegFile.scala 74:20:@52214.4]
  assign regs_178_clock = clock; // @[:@52223.4]
  assign regs_178_reset = io_reset; // @[:@52224.4 RegFile.scala 76:16:@52231.4]
  assign regs_178_io_in = 64'h0; // @[RegFile.scala 75:16:@52230.4]
  assign regs_178_io_reset = reset; // @[RegFile.scala 78:19:@52234.4]
  assign regs_178_io_enable = 1'h1; // @[RegFile.scala 74:20:@52228.4]
  assign regs_179_clock = clock; // @[:@52237.4]
  assign regs_179_reset = io_reset; // @[:@52238.4 RegFile.scala 76:16:@52245.4]
  assign regs_179_io_in = 64'h0; // @[RegFile.scala 75:16:@52244.4]
  assign regs_179_io_reset = reset; // @[RegFile.scala 78:19:@52248.4]
  assign regs_179_io_enable = 1'h1; // @[RegFile.scala 74:20:@52242.4]
  assign regs_180_clock = clock; // @[:@52251.4]
  assign regs_180_reset = io_reset; // @[:@52252.4 RegFile.scala 76:16:@52259.4]
  assign regs_180_io_in = 64'h0; // @[RegFile.scala 75:16:@52258.4]
  assign regs_180_io_reset = reset; // @[RegFile.scala 78:19:@52262.4]
  assign regs_180_io_enable = 1'h1; // @[RegFile.scala 74:20:@52256.4]
  assign regs_181_clock = clock; // @[:@52265.4]
  assign regs_181_reset = io_reset; // @[:@52266.4 RegFile.scala 76:16:@52273.4]
  assign regs_181_io_in = 64'h0; // @[RegFile.scala 75:16:@52272.4]
  assign regs_181_io_reset = reset; // @[RegFile.scala 78:19:@52276.4]
  assign regs_181_io_enable = 1'h1; // @[RegFile.scala 74:20:@52270.4]
  assign regs_182_clock = clock; // @[:@52279.4]
  assign regs_182_reset = io_reset; // @[:@52280.4 RegFile.scala 76:16:@52287.4]
  assign regs_182_io_in = 64'h0; // @[RegFile.scala 75:16:@52286.4]
  assign regs_182_io_reset = reset; // @[RegFile.scala 78:19:@52290.4]
  assign regs_182_io_enable = 1'h1; // @[RegFile.scala 74:20:@52284.4]
  assign regs_183_clock = clock; // @[:@52293.4]
  assign regs_183_reset = io_reset; // @[:@52294.4 RegFile.scala 76:16:@52301.4]
  assign regs_183_io_in = 64'h0; // @[RegFile.scala 75:16:@52300.4]
  assign regs_183_io_reset = reset; // @[RegFile.scala 78:19:@52304.4]
  assign regs_183_io_enable = 1'h1; // @[RegFile.scala 74:20:@52298.4]
  assign regs_184_clock = clock; // @[:@52307.4]
  assign regs_184_reset = io_reset; // @[:@52308.4 RegFile.scala 76:16:@52315.4]
  assign regs_184_io_in = 64'h0; // @[RegFile.scala 75:16:@52314.4]
  assign regs_184_io_reset = reset; // @[RegFile.scala 78:19:@52318.4]
  assign regs_184_io_enable = 1'h1; // @[RegFile.scala 74:20:@52312.4]
  assign regs_185_clock = clock; // @[:@52321.4]
  assign regs_185_reset = io_reset; // @[:@52322.4 RegFile.scala 76:16:@52329.4]
  assign regs_185_io_in = 64'h0; // @[RegFile.scala 75:16:@52328.4]
  assign regs_185_io_reset = reset; // @[RegFile.scala 78:19:@52332.4]
  assign regs_185_io_enable = 1'h1; // @[RegFile.scala 74:20:@52326.4]
  assign regs_186_clock = clock; // @[:@52335.4]
  assign regs_186_reset = io_reset; // @[:@52336.4 RegFile.scala 76:16:@52343.4]
  assign regs_186_io_in = 64'h0; // @[RegFile.scala 75:16:@52342.4]
  assign regs_186_io_reset = reset; // @[RegFile.scala 78:19:@52346.4]
  assign regs_186_io_enable = 1'h1; // @[RegFile.scala 74:20:@52340.4]
  assign regs_187_clock = clock; // @[:@52349.4]
  assign regs_187_reset = io_reset; // @[:@52350.4 RegFile.scala 76:16:@52357.4]
  assign regs_187_io_in = 64'h0; // @[RegFile.scala 75:16:@52356.4]
  assign regs_187_io_reset = reset; // @[RegFile.scala 78:19:@52360.4]
  assign regs_187_io_enable = 1'h1; // @[RegFile.scala 74:20:@52354.4]
  assign regs_188_clock = clock; // @[:@52363.4]
  assign regs_188_reset = io_reset; // @[:@52364.4 RegFile.scala 76:16:@52371.4]
  assign regs_188_io_in = 64'h0; // @[RegFile.scala 75:16:@52370.4]
  assign regs_188_io_reset = reset; // @[RegFile.scala 78:19:@52374.4]
  assign regs_188_io_enable = 1'h1; // @[RegFile.scala 74:20:@52368.4]
  assign regs_189_clock = clock; // @[:@52377.4]
  assign regs_189_reset = io_reset; // @[:@52378.4 RegFile.scala 76:16:@52385.4]
  assign regs_189_io_in = 64'h0; // @[RegFile.scala 75:16:@52384.4]
  assign regs_189_io_reset = reset; // @[RegFile.scala 78:19:@52388.4]
  assign regs_189_io_enable = 1'h1; // @[RegFile.scala 74:20:@52382.4]
  assign regs_190_clock = clock; // @[:@52391.4]
  assign regs_190_reset = io_reset; // @[:@52392.4 RegFile.scala 76:16:@52399.4]
  assign regs_190_io_in = 64'h0; // @[RegFile.scala 75:16:@52398.4]
  assign regs_190_io_reset = reset; // @[RegFile.scala 78:19:@52402.4]
  assign regs_190_io_enable = 1'h1; // @[RegFile.scala 74:20:@52396.4]
  assign regs_191_clock = clock; // @[:@52405.4]
  assign regs_191_reset = io_reset; // @[:@52406.4 RegFile.scala 76:16:@52413.4]
  assign regs_191_io_in = 64'h0; // @[RegFile.scala 75:16:@52412.4]
  assign regs_191_io_reset = reset; // @[RegFile.scala 78:19:@52416.4]
  assign regs_191_io_enable = 1'h1; // @[RegFile.scala 74:20:@52410.4]
  assign regs_192_clock = clock; // @[:@52419.4]
  assign regs_192_reset = io_reset; // @[:@52420.4 RegFile.scala 76:16:@52427.4]
  assign regs_192_io_in = 64'h0; // @[RegFile.scala 75:16:@52426.4]
  assign regs_192_io_reset = reset; // @[RegFile.scala 78:19:@52430.4]
  assign regs_192_io_enable = 1'h1; // @[RegFile.scala 74:20:@52424.4]
  assign regs_193_clock = clock; // @[:@52433.4]
  assign regs_193_reset = io_reset; // @[:@52434.4 RegFile.scala 76:16:@52441.4]
  assign regs_193_io_in = 64'h0; // @[RegFile.scala 75:16:@52440.4]
  assign regs_193_io_reset = reset; // @[RegFile.scala 78:19:@52444.4]
  assign regs_193_io_enable = 1'h1; // @[RegFile.scala 74:20:@52438.4]
  assign regs_194_clock = clock; // @[:@52447.4]
  assign regs_194_reset = io_reset; // @[:@52448.4 RegFile.scala 76:16:@52455.4]
  assign regs_194_io_in = 64'h0; // @[RegFile.scala 75:16:@52454.4]
  assign regs_194_io_reset = reset; // @[RegFile.scala 78:19:@52458.4]
  assign regs_194_io_enable = 1'h1; // @[RegFile.scala 74:20:@52452.4]
  assign regs_195_clock = clock; // @[:@52461.4]
  assign regs_195_reset = io_reset; // @[:@52462.4 RegFile.scala 76:16:@52469.4]
  assign regs_195_io_in = 64'h0; // @[RegFile.scala 75:16:@52468.4]
  assign regs_195_io_reset = reset; // @[RegFile.scala 78:19:@52472.4]
  assign regs_195_io_enable = 1'h1; // @[RegFile.scala 74:20:@52466.4]
  assign regs_196_clock = clock; // @[:@52475.4]
  assign regs_196_reset = io_reset; // @[:@52476.4 RegFile.scala 76:16:@52483.4]
  assign regs_196_io_in = 64'h0; // @[RegFile.scala 75:16:@52482.4]
  assign regs_196_io_reset = reset; // @[RegFile.scala 78:19:@52486.4]
  assign regs_196_io_enable = 1'h1; // @[RegFile.scala 74:20:@52480.4]
  assign regs_197_clock = clock; // @[:@52489.4]
  assign regs_197_reset = io_reset; // @[:@52490.4 RegFile.scala 76:16:@52497.4]
  assign regs_197_io_in = 64'h0; // @[RegFile.scala 75:16:@52496.4]
  assign regs_197_io_reset = reset; // @[RegFile.scala 78:19:@52500.4]
  assign regs_197_io_enable = 1'h1; // @[RegFile.scala 74:20:@52494.4]
  assign regs_198_clock = clock; // @[:@52503.4]
  assign regs_198_reset = io_reset; // @[:@52504.4 RegFile.scala 76:16:@52511.4]
  assign regs_198_io_in = 64'h0; // @[RegFile.scala 75:16:@52510.4]
  assign regs_198_io_reset = reset; // @[RegFile.scala 78:19:@52514.4]
  assign regs_198_io_enable = 1'h1; // @[RegFile.scala 74:20:@52508.4]
  assign regs_199_clock = clock; // @[:@52517.4]
  assign regs_199_reset = io_reset; // @[:@52518.4 RegFile.scala 76:16:@52525.4]
  assign regs_199_io_in = 64'h0; // @[RegFile.scala 75:16:@52524.4]
  assign regs_199_io_reset = reset; // @[RegFile.scala 78:19:@52528.4]
  assign regs_199_io_enable = 1'h1; // @[RegFile.scala 74:20:@52522.4]
  assign regs_200_clock = clock; // @[:@52531.4]
  assign regs_200_reset = io_reset; // @[:@52532.4 RegFile.scala 76:16:@52539.4]
  assign regs_200_io_in = 64'h0; // @[RegFile.scala 75:16:@52538.4]
  assign regs_200_io_reset = reset; // @[RegFile.scala 78:19:@52542.4]
  assign regs_200_io_enable = 1'h1; // @[RegFile.scala 74:20:@52536.4]
  assign regs_201_clock = clock; // @[:@52545.4]
  assign regs_201_reset = io_reset; // @[:@52546.4 RegFile.scala 76:16:@52553.4]
  assign regs_201_io_in = 64'h0; // @[RegFile.scala 75:16:@52552.4]
  assign regs_201_io_reset = reset; // @[RegFile.scala 78:19:@52556.4]
  assign regs_201_io_enable = 1'h1; // @[RegFile.scala 74:20:@52550.4]
  assign regs_202_clock = clock; // @[:@52559.4]
  assign regs_202_reset = io_reset; // @[:@52560.4 RegFile.scala 76:16:@52567.4]
  assign regs_202_io_in = 64'h0; // @[RegFile.scala 75:16:@52566.4]
  assign regs_202_io_reset = reset; // @[RegFile.scala 78:19:@52570.4]
  assign regs_202_io_enable = 1'h1; // @[RegFile.scala 74:20:@52564.4]
  assign regs_203_clock = clock; // @[:@52573.4]
  assign regs_203_reset = io_reset; // @[:@52574.4 RegFile.scala 76:16:@52581.4]
  assign regs_203_io_in = 64'h0; // @[RegFile.scala 75:16:@52580.4]
  assign regs_203_io_reset = reset; // @[RegFile.scala 78:19:@52584.4]
  assign regs_203_io_enable = 1'h1; // @[RegFile.scala 74:20:@52578.4]
  assign regs_204_clock = clock; // @[:@52587.4]
  assign regs_204_reset = io_reset; // @[:@52588.4 RegFile.scala 76:16:@52595.4]
  assign regs_204_io_in = 64'h0; // @[RegFile.scala 75:16:@52594.4]
  assign regs_204_io_reset = reset; // @[RegFile.scala 78:19:@52598.4]
  assign regs_204_io_enable = 1'h1; // @[RegFile.scala 74:20:@52592.4]
  assign regs_205_clock = clock; // @[:@52601.4]
  assign regs_205_reset = io_reset; // @[:@52602.4 RegFile.scala 76:16:@52609.4]
  assign regs_205_io_in = 64'h0; // @[RegFile.scala 75:16:@52608.4]
  assign regs_205_io_reset = reset; // @[RegFile.scala 78:19:@52612.4]
  assign regs_205_io_enable = 1'h1; // @[RegFile.scala 74:20:@52606.4]
  assign regs_206_clock = clock; // @[:@52615.4]
  assign regs_206_reset = io_reset; // @[:@52616.4 RegFile.scala 76:16:@52623.4]
  assign regs_206_io_in = 64'h0; // @[RegFile.scala 75:16:@52622.4]
  assign regs_206_io_reset = reset; // @[RegFile.scala 78:19:@52626.4]
  assign regs_206_io_enable = 1'h1; // @[RegFile.scala 74:20:@52620.4]
  assign regs_207_clock = clock; // @[:@52629.4]
  assign regs_207_reset = io_reset; // @[:@52630.4 RegFile.scala 76:16:@52637.4]
  assign regs_207_io_in = 64'h0; // @[RegFile.scala 75:16:@52636.4]
  assign regs_207_io_reset = reset; // @[RegFile.scala 78:19:@52640.4]
  assign regs_207_io_enable = 1'h1; // @[RegFile.scala 74:20:@52634.4]
  assign regs_208_clock = clock; // @[:@52643.4]
  assign regs_208_reset = io_reset; // @[:@52644.4 RegFile.scala 76:16:@52651.4]
  assign regs_208_io_in = 64'h0; // @[RegFile.scala 75:16:@52650.4]
  assign regs_208_io_reset = reset; // @[RegFile.scala 78:19:@52654.4]
  assign regs_208_io_enable = 1'h1; // @[RegFile.scala 74:20:@52648.4]
  assign regs_209_clock = clock; // @[:@52657.4]
  assign regs_209_reset = io_reset; // @[:@52658.4 RegFile.scala 76:16:@52665.4]
  assign regs_209_io_in = 64'h0; // @[RegFile.scala 75:16:@52664.4]
  assign regs_209_io_reset = reset; // @[RegFile.scala 78:19:@52668.4]
  assign regs_209_io_enable = 1'h1; // @[RegFile.scala 74:20:@52662.4]
  assign regs_210_clock = clock; // @[:@52671.4]
  assign regs_210_reset = io_reset; // @[:@52672.4 RegFile.scala 76:16:@52679.4]
  assign regs_210_io_in = 64'h0; // @[RegFile.scala 75:16:@52678.4]
  assign regs_210_io_reset = reset; // @[RegFile.scala 78:19:@52682.4]
  assign regs_210_io_enable = 1'h1; // @[RegFile.scala 74:20:@52676.4]
  assign regs_211_clock = clock; // @[:@52685.4]
  assign regs_211_reset = io_reset; // @[:@52686.4 RegFile.scala 76:16:@52693.4]
  assign regs_211_io_in = 64'h0; // @[RegFile.scala 75:16:@52692.4]
  assign regs_211_io_reset = reset; // @[RegFile.scala 78:19:@52696.4]
  assign regs_211_io_enable = 1'h1; // @[RegFile.scala 74:20:@52690.4]
  assign regs_212_clock = clock; // @[:@52699.4]
  assign regs_212_reset = io_reset; // @[:@52700.4 RegFile.scala 76:16:@52707.4]
  assign regs_212_io_in = 64'h0; // @[RegFile.scala 75:16:@52706.4]
  assign regs_212_io_reset = reset; // @[RegFile.scala 78:19:@52710.4]
  assign regs_212_io_enable = 1'h1; // @[RegFile.scala 74:20:@52704.4]
  assign regs_213_clock = clock; // @[:@52713.4]
  assign regs_213_reset = io_reset; // @[:@52714.4 RegFile.scala 76:16:@52721.4]
  assign regs_213_io_in = 64'h0; // @[RegFile.scala 75:16:@52720.4]
  assign regs_213_io_reset = reset; // @[RegFile.scala 78:19:@52724.4]
  assign regs_213_io_enable = 1'h1; // @[RegFile.scala 74:20:@52718.4]
  assign regs_214_clock = clock; // @[:@52727.4]
  assign regs_214_reset = io_reset; // @[:@52728.4 RegFile.scala 76:16:@52735.4]
  assign regs_214_io_in = 64'h0; // @[RegFile.scala 75:16:@52734.4]
  assign regs_214_io_reset = reset; // @[RegFile.scala 78:19:@52738.4]
  assign regs_214_io_enable = 1'h1; // @[RegFile.scala 74:20:@52732.4]
  assign regs_215_clock = clock; // @[:@52741.4]
  assign regs_215_reset = io_reset; // @[:@52742.4 RegFile.scala 76:16:@52749.4]
  assign regs_215_io_in = 64'h0; // @[RegFile.scala 75:16:@52748.4]
  assign regs_215_io_reset = reset; // @[RegFile.scala 78:19:@52752.4]
  assign regs_215_io_enable = 1'h1; // @[RegFile.scala 74:20:@52746.4]
  assign regs_216_clock = clock; // @[:@52755.4]
  assign regs_216_reset = io_reset; // @[:@52756.4 RegFile.scala 76:16:@52763.4]
  assign regs_216_io_in = 64'h0; // @[RegFile.scala 75:16:@52762.4]
  assign regs_216_io_reset = reset; // @[RegFile.scala 78:19:@52766.4]
  assign regs_216_io_enable = 1'h1; // @[RegFile.scala 74:20:@52760.4]
  assign regs_217_clock = clock; // @[:@52769.4]
  assign regs_217_reset = io_reset; // @[:@52770.4 RegFile.scala 76:16:@52777.4]
  assign regs_217_io_in = 64'h0; // @[RegFile.scala 75:16:@52776.4]
  assign regs_217_io_reset = reset; // @[RegFile.scala 78:19:@52780.4]
  assign regs_217_io_enable = 1'h1; // @[RegFile.scala 74:20:@52774.4]
  assign regs_218_clock = clock; // @[:@52783.4]
  assign regs_218_reset = io_reset; // @[:@52784.4 RegFile.scala 76:16:@52791.4]
  assign regs_218_io_in = 64'h0; // @[RegFile.scala 75:16:@52790.4]
  assign regs_218_io_reset = reset; // @[RegFile.scala 78:19:@52794.4]
  assign regs_218_io_enable = 1'h1; // @[RegFile.scala 74:20:@52788.4]
  assign regs_219_clock = clock; // @[:@52797.4]
  assign regs_219_reset = io_reset; // @[:@52798.4 RegFile.scala 76:16:@52805.4]
  assign regs_219_io_in = 64'h0; // @[RegFile.scala 75:16:@52804.4]
  assign regs_219_io_reset = reset; // @[RegFile.scala 78:19:@52808.4]
  assign regs_219_io_enable = 1'h1; // @[RegFile.scala 74:20:@52802.4]
  assign regs_220_clock = clock; // @[:@52811.4]
  assign regs_220_reset = io_reset; // @[:@52812.4 RegFile.scala 76:16:@52819.4]
  assign regs_220_io_in = 64'h0; // @[RegFile.scala 75:16:@52818.4]
  assign regs_220_io_reset = reset; // @[RegFile.scala 78:19:@52822.4]
  assign regs_220_io_enable = 1'h1; // @[RegFile.scala 74:20:@52816.4]
  assign regs_221_clock = clock; // @[:@52825.4]
  assign regs_221_reset = io_reset; // @[:@52826.4 RegFile.scala 76:16:@52833.4]
  assign regs_221_io_in = 64'h0; // @[RegFile.scala 75:16:@52832.4]
  assign regs_221_io_reset = reset; // @[RegFile.scala 78:19:@52836.4]
  assign regs_221_io_enable = 1'h1; // @[RegFile.scala 74:20:@52830.4]
  assign regs_222_clock = clock; // @[:@52839.4]
  assign regs_222_reset = io_reset; // @[:@52840.4 RegFile.scala 76:16:@52847.4]
  assign regs_222_io_in = 64'h0; // @[RegFile.scala 75:16:@52846.4]
  assign regs_222_io_reset = reset; // @[RegFile.scala 78:19:@52850.4]
  assign regs_222_io_enable = 1'h1; // @[RegFile.scala 74:20:@52844.4]
  assign regs_223_clock = clock; // @[:@52853.4]
  assign regs_223_reset = io_reset; // @[:@52854.4 RegFile.scala 76:16:@52861.4]
  assign regs_223_io_in = 64'h0; // @[RegFile.scala 75:16:@52860.4]
  assign regs_223_io_reset = reset; // @[RegFile.scala 78:19:@52864.4]
  assign regs_223_io_enable = 1'h1; // @[RegFile.scala 74:20:@52858.4]
  assign regs_224_clock = clock; // @[:@52867.4]
  assign regs_224_reset = io_reset; // @[:@52868.4 RegFile.scala 76:16:@52875.4]
  assign regs_224_io_in = 64'h0; // @[RegFile.scala 75:16:@52874.4]
  assign regs_224_io_reset = reset; // @[RegFile.scala 78:19:@52878.4]
  assign regs_224_io_enable = 1'h1; // @[RegFile.scala 74:20:@52872.4]
  assign regs_225_clock = clock; // @[:@52881.4]
  assign regs_225_reset = io_reset; // @[:@52882.4 RegFile.scala 76:16:@52889.4]
  assign regs_225_io_in = 64'h0; // @[RegFile.scala 75:16:@52888.4]
  assign regs_225_io_reset = reset; // @[RegFile.scala 78:19:@52892.4]
  assign regs_225_io_enable = 1'h1; // @[RegFile.scala 74:20:@52886.4]
  assign regs_226_clock = clock; // @[:@52895.4]
  assign regs_226_reset = io_reset; // @[:@52896.4 RegFile.scala 76:16:@52903.4]
  assign regs_226_io_in = 64'h0; // @[RegFile.scala 75:16:@52902.4]
  assign regs_226_io_reset = reset; // @[RegFile.scala 78:19:@52906.4]
  assign regs_226_io_enable = 1'h1; // @[RegFile.scala 74:20:@52900.4]
  assign regs_227_clock = clock; // @[:@52909.4]
  assign regs_227_reset = io_reset; // @[:@52910.4 RegFile.scala 76:16:@52917.4]
  assign regs_227_io_in = 64'h0; // @[RegFile.scala 75:16:@52916.4]
  assign regs_227_io_reset = reset; // @[RegFile.scala 78:19:@52920.4]
  assign regs_227_io_enable = 1'h1; // @[RegFile.scala 74:20:@52914.4]
  assign regs_228_clock = clock; // @[:@52923.4]
  assign regs_228_reset = io_reset; // @[:@52924.4 RegFile.scala 76:16:@52931.4]
  assign regs_228_io_in = 64'h0; // @[RegFile.scala 75:16:@52930.4]
  assign regs_228_io_reset = reset; // @[RegFile.scala 78:19:@52934.4]
  assign regs_228_io_enable = 1'h1; // @[RegFile.scala 74:20:@52928.4]
  assign regs_229_clock = clock; // @[:@52937.4]
  assign regs_229_reset = io_reset; // @[:@52938.4 RegFile.scala 76:16:@52945.4]
  assign regs_229_io_in = 64'h0; // @[RegFile.scala 75:16:@52944.4]
  assign regs_229_io_reset = reset; // @[RegFile.scala 78:19:@52948.4]
  assign regs_229_io_enable = 1'h1; // @[RegFile.scala 74:20:@52942.4]
  assign regs_230_clock = clock; // @[:@52951.4]
  assign regs_230_reset = io_reset; // @[:@52952.4 RegFile.scala 76:16:@52959.4]
  assign regs_230_io_in = 64'h0; // @[RegFile.scala 75:16:@52958.4]
  assign regs_230_io_reset = reset; // @[RegFile.scala 78:19:@52962.4]
  assign regs_230_io_enable = 1'h1; // @[RegFile.scala 74:20:@52956.4]
  assign regs_231_clock = clock; // @[:@52965.4]
  assign regs_231_reset = io_reset; // @[:@52966.4 RegFile.scala 76:16:@52973.4]
  assign regs_231_io_in = 64'h0; // @[RegFile.scala 75:16:@52972.4]
  assign regs_231_io_reset = reset; // @[RegFile.scala 78:19:@52976.4]
  assign regs_231_io_enable = 1'h1; // @[RegFile.scala 74:20:@52970.4]
  assign regs_232_clock = clock; // @[:@52979.4]
  assign regs_232_reset = io_reset; // @[:@52980.4 RegFile.scala 76:16:@52987.4]
  assign regs_232_io_in = 64'h0; // @[RegFile.scala 75:16:@52986.4]
  assign regs_232_io_reset = reset; // @[RegFile.scala 78:19:@52990.4]
  assign regs_232_io_enable = 1'h1; // @[RegFile.scala 74:20:@52984.4]
  assign regs_233_clock = clock; // @[:@52993.4]
  assign regs_233_reset = io_reset; // @[:@52994.4 RegFile.scala 76:16:@53001.4]
  assign regs_233_io_in = 64'h0; // @[RegFile.scala 75:16:@53000.4]
  assign regs_233_io_reset = reset; // @[RegFile.scala 78:19:@53004.4]
  assign regs_233_io_enable = 1'h1; // @[RegFile.scala 74:20:@52998.4]
  assign regs_234_clock = clock; // @[:@53007.4]
  assign regs_234_reset = io_reset; // @[:@53008.4 RegFile.scala 76:16:@53015.4]
  assign regs_234_io_in = 64'h0; // @[RegFile.scala 75:16:@53014.4]
  assign regs_234_io_reset = reset; // @[RegFile.scala 78:19:@53018.4]
  assign regs_234_io_enable = 1'h1; // @[RegFile.scala 74:20:@53012.4]
  assign regs_235_clock = clock; // @[:@53021.4]
  assign regs_235_reset = io_reset; // @[:@53022.4 RegFile.scala 76:16:@53029.4]
  assign regs_235_io_in = 64'h0; // @[RegFile.scala 75:16:@53028.4]
  assign regs_235_io_reset = reset; // @[RegFile.scala 78:19:@53032.4]
  assign regs_235_io_enable = 1'h1; // @[RegFile.scala 74:20:@53026.4]
  assign regs_236_clock = clock; // @[:@53035.4]
  assign regs_236_reset = io_reset; // @[:@53036.4 RegFile.scala 76:16:@53043.4]
  assign regs_236_io_in = 64'h0; // @[RegFile.scala 75:16:@53042.4]
  assign regs_236_io_reset = reset; // @[RegFile.scala 78:19:@53046.4]
  assign regs_236_io_enable = 1'h1; // @[RegFile.scala 74:20:@53040.4]
  assign regs_237_clock = clock; // @[:@53049.4]
  assign regs_237_reset = io_reset; // @[:@53050.4 RegFile.scala 76:16:@53057.4]
  assign regs_237_io_in = 64'h0; // @[RegFile.scala 75:16:@53056.4]
  assign regs_237_io_reset = reset; // @[RegFile.scala 78:19:@53060.4]
  assign regs_237_io_enable = 1'h1; // @[RegFile.scala 74:20:@53054.4]
  assign regs_238_clock = clock; // @[:@53063.4]
  assign regs_238_reset = io_reset; // @[:@53064.4 RegFile.scala 76:16:@53071.4]
  assign regs_238_io_in = 64'h0; // @[RegFile.scala 75:16:@53070.4]
  assign regs_238_io_reset = reset; // @[RegFile.scala 78:19:@53074.4]
  assign regs_238_io_enable = 1'h1; // @[RegFile.scala 74:20:@53068.4]
  assign regs_239_clock = clock; // @[:@53077.4]
  assign regs_239_reset = io_reset; // @[:@53078.4 RegFile.scala 76:16:@53085.4]
  assign regs_239_io_in = 64'h0; // @[RegFile.scala 75:16:@53084.4]
  assign regs_239_io_reset = reset; // @[RegFile.scala 78:19:@53088.4]
  assign regs_239_io_enable = 1'h1; // @[RegFile.scala 74:20:@53082.4]
  assign regs_240_clock = clock; // @[:@53091.4]
  assign regs_240_reset = io_reset; // @[:@53092.4 RegFile.scala 76:16:@53099.4]
  assign regs_240_io_in = 64'h0; // @[RegFile.scala 75:16:@53098.4]
  assign regs_240_io_reset = reset; // @[RegFile.scala 78:19:@53102.4]
  assign regs_240_io_enable = 1'h1; // @[RegFile.scala 74:20:@53096.4]
  assign regs_241_clock = clock; // @[:@53105.4]
  assign regs_241_reset = io_reset; // @[:@53106.4 RegFile.scala 76:16:@53113.4]
  assign regs_241_io_in = 64'h0; // @[RegFile.scala 75:16:@53112.4]
  assign regs_241_io_reset = reset; // @[RegFile.scala 78:19:@53116.4]
  assign regs_241_io_enable = 1'h1; // @[RegFile.scala 74:20:@53110.4]
  assign regs_242_clock = clock; // @[:@53119.4]
  assign regs_242_reset = io_reset; // @[:@53120.4 RegFile.scala 76:16:@53127.4]
  assign regs_242_io_in = 64'h0; // @[RegFile.scala 75:16:@53126.4]
  assign regs_242_io_reset = reset; // @[RegFile.scala 78:19:@53130.4]
  assign regs_242_io_enable = 1'h1; // @[RegFile.scala 74:20:@53124.4]
  assign regs_243_clock = clock; // @[:@53133.4]
  assign regs_243_reset = io_reset; // @[:@53134.4 RegFile.scala 76:16:@53141.4]
  assign regs_243_io_in = 64'h0; // @[RegFile.scala 75:16:@53140.4]
  assign regs_243_io_reset = reset; // @[RegFile.scala 78:19:@53144.4]
  assign regs_243_io_enable = 1'h1; // @[RegFile.scala 74:20:@53138.4]
  assign regs_244_clock = clock; // @[:@53147.4]
  assign regs_244_reset = io_reset; // @[:@53148.4 RegFile.scala 76:16:@53155.4]
  assign regs_244_io_in = 64'h0; // @[RegFile.scala 75:16:@53154.4]
  assign regs_244_io_reset = reset; // @[RegFile.scala 78:19:@53158.4]
  assign regs_244_io_enable = 1'h1; // @[RegFile.scala 74:20:@53152.4]
  assign regs_245_clock = clock; // @[:@53161.4]
  assign regs_245_reset = io_reset; // @[:@53162.4 RegFile.scala 76:16:@53169.4]
  assign regs_245_io_in = 64'h0; // @[RegFile.scala 75:16:@53168.4]
  assign regs_245_io_reset = reset; // @[RegFile.scala 78:19:@53172.4]
  assign regs_245_io_enable = 1'h1; // @[RegFile.scala 74:20:@53166.4]
  assign regs_246_clock = clock; // @[:@53175.4]
  assign regs_246_reset = io_reset; // @[:@53176.4 RegFile.scala 76:16:@53183.4]
  assign regs_246_io_in = 64'h0; // @[RegFile.scala 75:16:@53182.4]
  assign regs_246_io_reset = reset; // @[RegFile.scala 78:19:@53186.4]
  assign regs_246_io_enable = 1'h1; // @[RegFile.scala 74:20:@53180.4]
  assign regs_247_clock = clock; // @[:@53189.4]
  assign regs_247_reset = io_reset; // @[:@53190.4 RegFile.scala 76:16:@53197.4]
  assign regs_247_io_in = 64'h0; // @[RegFile.scala 75:16:@53196.4]
  assign regs_247_io_reset = reset; // @[RegFile.scala 78:19:@53200.4]
  assign regs_247_io_enable = 1'h1; // @[RegFile.scala 74:20:@53194.4]
  assign regs_248_clock = clock; // @[:@53203.4]
  assign regs_248_reset = io_reset; // @[:@53204.4 RegFile.scala 76:16:@53211.4]
  assign regs_248_io_in = 64'h0; // @[RegFile.scala 75:16:@53210.4]
  assign regs_248_io_reset = reset; // @[RegFile.scala 78:19:@53214.4]
  assign regs_248_io_enable = 1'h1; // @[RegFile.scala 74:20:@53208.4]
  assign regs_249_clock = clock; // @[:@53217.4]
  assign regs_249_reset = io_reset; // @[:@53218.4 RegFile.scala 76:16:@53225.4]
  assign regs_249_io_in = 64'h0; // @[RegFile.scala 75:16:@53224.4]
  assign regs_249_io_reset = reset; // @[RegFile.scala 78:19:@53228.4]
  assign regs_249_io_enable = 1'h1; // @[RegFile.scala 74:20:@53222.4]
  assign regs_250_clock = clock; // @[:@53231.4]
  assign regs_250_reset = io_reset; // @[:@53232.4 RegFile.scala 76:16:@53239.4]
  assign regs_250_io_in = 64'h0; // @[RegFile.scala 75:16:@53238.4]
  assign regs_250_io_reset = reset; // @[RegFile.scala 78:19:@53242.4]
  assign regs_250_io_enable = 1'h1; // @[RegFile.scala 74:20:@53236.4]
  assign regs_251_clock = clock; // @[:@53245.4]
  assign regs_251_reset = io_reset; // @[:@53246.4 RegFile.scala 76:16:@53253.4]
  assign regs_251_io_in = 64'h0; // @[RegFile.scala 75:16:@53252.4]
  assign regs_251_io_reset = reset; // @[RegFile.scala 78:19:@53256.4]
  assign regs_251_io_enable = 1'h1; // @[RegFile.scala 74:20:@53250.4]
  assign regs_252_clock = clock; // @[:@53259.4]
  assign regs_252_reset = io_reset; // @[:@53260.4 RegFile.scala 76:16:@53267.4]
  assign regs_252_io_in = 64'h0; // @[RegFile.scala 75:16:@53266.4]
  assign regs_252_io_reset = reset; // @[RegFile.scala 78:19:@53270.4]
  assign regs_252_io_enable = 1'h1; // @[RegFile.scala 74:20:@53264.4]
  assign regs_253_clock = clock; // @[:@53273.4]
  assign regs_253_reset = io_reset; // @[:@53274.4 RegFile.scala 76:16:@53281.4]
  assign regs_253_io_in = 64'h0; // @[RegFile.scala 75:16:@53280.4]
  assign regs_253_io_reset = reset; // @[RegFile.scala 78:19:@53284.4]
  assign regs_253_io_enable = 1'h1; // @[RegFile.scala 74:20:@53278.4]
  assign regs_254_clock = clock; // @[:@53287.4]
  assign regs_254_reset = io_reset; // @[:@53288.4 RegFile.scala 76:16:@53295.4]
  assign regs_254_io_in = 64'h0; // @[RegFile.scala 75:16:@53294.4]
  assign regs_254_io_reset = reset; // @[RegFile.scala 78:19:@53298.4]
  assign regs_254_io_enable = 1'h1; // @[RegFile.scala 74:20:@53292.4]
  assign regs_255_clock = clock; // @[:@53301.4]
  assign regs_255_reset = io_reset; // @[:@53302.4 RegFile.scala 76:16:@53309.4]
  assign regs_255_io_in = 64'h0; // @[RegFile.scala 75:16:@53308.4]
  assign regs_255_io_reset = reset; // @[RegFile.scala 78:19:@53312.4]
  assign regs_255_io_enable = 1'h1; // @[RegFile.scala 74:20:@53306.4]
  assign regs_256_clock = clock; // @[:@53315.4]
  assign regs_256_reset = io_reset; // @[:@53316.4 RegFile.scala 76:16:@53323.4]
  assign regs_256_io_in = 64'h0; // @[RegFile.scala 75:16:@53322.4]
  assign regs_256_io_reset = reset; // @[RegFile.scala 78:19:@53326.4]
  assign regs_256_io_enable = 1'h1; // @[RegFile.scala 74:20:@53320.4]
  assign regs_257_clock = clock; // @[:@53329.4]
  assign regs_257_reset = io_reset; // @[:@53330.4 RegFile.scala 76:16:@53337.4]
  assign regs_257_io_in = 64'h0; // @[RegFile.scala 75:16:@53336.4]
  assign regs_257_io_reset = reset; // @[RegFile.scala 78:19:@53340.4]
  assign regs_257_io_enable = 1'h1; // @[RegFile.scala 74:20:@53334.4]
  assign regs_258_clock = clock; // @[:@53343.4]
  assign regs_258_reset = io_reset; // @[:@53344.4 RegFile.scala 76:16:@53351.4]
  assign regs_258_io_in = 64'h0; // @[RegFile.scala 75:16:@53350.4]
  assign regs_258_io_reset = reset; // @[RegFile.scala 78:19:@53354.4]
  assign regs_258_io_enable = 1'h1; // @[RegFile.scala 74:20:@53348.4]
  assign regs_259_clock = clock; // @[:@53357.4]
  assign regs_259_reset = io_reset; // @[:@53358.4 RegFile.scala 76:16:@53365.4]
  assign regs_259_io_in = 64'h0; // @[RegFile.scala 75:16:@53364.4]
  assign regs_259_io_reset = reset; // @[RegFile.scala 78:19:@53368.4]
  assign regs_259_io_enable = 1'h1; // @[RegFile.scala 74:20:@53362.4]
  assign regs_260_clock = clock; // @[:@53371.4]
  assign regs_260_reset = io_reset; // @[:@53372.4 RegFile.scala 76:16:@53379.4]
  assign regs_260_io_in = 64'h0; // @[RegFile.scala 75:16:@53378.4]
  assign regs_260_io_reset = reset; // @[RegFile.scala 78:19:@53382.4]
  assign regs_260_io_enable = 1'h1; // @[RegFile.scala 74:20:@53376.4]
  assign regs_261_clock = clock; // @[:@53385.4]
  assign regs_261_reset = io_reset; // @[:@53386.4 RegFile.scala 76:16:@53393.4]
  assign regs_261_io_in = 64'h0; // @[RegFile.scala 75:16:@53392.4]
  assign regs_261_io_reset = reset; // @[RegFile.scala 78:19:@53396.4]
  assign regs_261_io_enable = 1'h1; // @[RegFile.scala 74:20:@53390.4]
  assign regs_262_clock = clock; // @[:@53399.4]
  assign regs_262_reset = io_reset; // @[:@53400.4 RegFile.scala 76:16:@53407.4]
  assign regs_262_io_in = 64'h0; // @[RegFile.scala 75:16:@53406.4]
  assign regs_262_io_reset = reset; // @[RegFile.scala 78:19:@53410.4]
  assign regs_262_io_enable = 1'h1; // @[RegFile.scala 74:20:@53404.4]
  assign regs_263_clock = clock; // @[:@53413.4]
  assign regs_263_reset = io_reset; // @[:@53414.4 RegFile.scala 76:16:@53421.4]
  assign regs_263_io_in = 64'h0; // @[RegFile.scala 75:16:@53420.4]
  assign regs_263_io_reset = reset; // @[RegFile.scala 78:19:@53424.4]
  assign regs_263_io_enable = 1'h1; // @[RegFile.scala 74:20:@53418.4]
  assign regs_264_clock = clock; // @[:@53427.4]
  assign regs_264_reset = io_reset; // @[:@53428.4 RegFile.scala 76:16:@53435.4]
  assign regs_264_io_in = 64'h0; // @[RegFile.scala 75:16:@53434.4]
  assign regs_264_io_reset = reset; // @[RegFile.scala 78:19:@53438.4]
  assign regs_264_io_enable = 1'h1; // @[RegFile.scala 74:20:@53432.4]
  assign regs_265_clock = clock; // @[:@53441.4]
  assign regs_265_reset = io_reset; // @[:@53442.4 RegFile.scala 76:16:@53449.4]
  assign regs_265_io_in = 64'h0; // @[RegFile.scala 75:16:@53448.4]
  assign regs_265_io_reset = reset; // @[RegFile.scala 78:19:@53452.4]
  assign regs_265_io_enable = 1'h1; // @[RegFile.scala 74:20:@53446.4]
  assign regs_266_clock = clock; // @[:@53455.4]
  assign regs_266_reset = io_reset; // @[:@53456.4 RegFile.scala 76:16:@53463.4]
  assign regs_266_io_in = 64'h0; // @[RegFile.scala 75:16:@53462.4]
  assign regs_266_io_reset = reset; // @[RegFile.scala 78:19:@53466.4]
  assign regs_266_io_enable = 1'h1; // @[RegFile.scala 74:20:@53460.4]
  assign regs_267_clock = clock; // @[:@53469.4]
  assign regs_267_reset = io_reset; // @[:@53470.4 RegFile.scala 76:16:@53477.4]
  assign regs_267_io_in = 64'h0; // @[RegFile.scala 75:16:@53476.4]
  assign regs_267_io_reset = reset; // @[RegFile.scala 78:19:@53480.4]
  assign regs_267_io_enable = 1'h1; // @[RegFile.scala 74:20:@53474.4]
  assign regs_268_clock = clock; // @[:@53483.4]
  assign regs_268_reset = io_reset; // @[:@53484.4 RegFile.scala 76:16:@53491.4]
  assign regs_268_io_in = 64'h0; // @[RegFile.scala 75:16:@53490.4]
  assign regs_268_io_reset = reset; // @[RegFile.scala 78:19:@53494.4]
  assign regs_268_io_enable = 1'h1; // @[RegFile.scala 74:20:@53488.4]
  assign regs_269_clock = clock; // @[:@53497.4]
  assign regs_269_reset = io_reset; // @[:@53498.4 RegFile.scala 76:16:@53505.4]
  assign regs_269_io_in = 64'h0; // @[RegFile.scala 75:16:@53504.4]
  assign regs_269_io_reset = reset; // @[RegFile.scala 78:19:@53508.4]
  assign regs_269_io_enable = 1'h1; // @[RegFile.scala 74:20:@53502.4]
  assign regs_270_clock = clock; // @[:@53511.4]
  assign regs_270_reset = io_reset; // @[:@53512.4 RegFile.scala 76:16:@53519.4]
  assign regs_270_io_in = 64'h0; // @[RegFile.scala 75:16:@53518.4]
  assign regs_270_io_reset = reset; // @[RegFile.scala 78:19:@53522.4]
  assign regs_270_io_enable = 1'h1; // @[RegFile.scala 74:20:@53516.4]
  assign regs_271_clock = clock; // @[:@53525.4]
  assign regs_271_reset = io_reset; // @[:@53526.4 RegFile.scala 76:16:@53533.4]
  assign regs_271_io_in = 64'h0; // @[RegFile.scala 75:16:@53532.4]
  assign regs_271_io_reset = reset; // @[RegFile.scala 78:19:@53536.4]
  assign regs_271_io_enable = 1'h1; // @[RegFile.scala 74:20:@53530.4]
  assign regs_272_clock = clock; // @[:@53539.4]
  assign regs_272_reset = io_reset; // @[:@53540.4 RegFile.scala 76:16:@53547.4]
  assign regs_272_io_in = 64'h0; // @[RegFile.scala 75:16:@53546.4]
  assign regs_272_io_reset = reset; // @[RegFile.scala 78:19:@53550.4]
  assign regs_272_io_enable = 1'h1; // @[RegFile.scala 74:20:@53544.4]
  assign regs_273_clock = clock; // @[:@53553.4]
  assign regs_273_reset = io_reset; // @[:@53554.4 RegFile.scala 76:16:@53561.4]
  assign regs_273_io_in = 64'h0; // @[RegFile.scala 75:16:@53560.4]
  assign regs_273_io_reset = reset; // @[RegFile.scala 78:19:@53564.4]
  assign regs_273_io_enable = 1'h1; // @[RegFile.scala 74:20:@53558.4]
  assign regs_274_clock = clock; // @[:@53567.4]
  assign regs_274_reset = io_reset; // @[:@53568.4 RegFile.scala 76:16:@53575.4]
  assign regs_274_io_in = 64'h0; // @[RegFile.scala 75:16:@53574.4]
  assign regs_274_io_reset = reset; // @[RegFile.scala 78:19:@53578.4]
  assign regs_274_io_enable = 1'h1; // @[RegFile.scala 74:20:@53572.4]
  assign regs_275_clock = clock; // @[:@53581.4]
  assign regs_275_reset = io_reset; // @[:@53582.4 RegFile.scala 76:16:@53589.4]
  assign regs_275_io_in = 64'h0; // @[RegFile.scala 75:16:@53588.4]
  assign regs_275_io_reset = reset; // @[RegFile.scala 78:19:@53592.4]
  assign regs_275_io_enable = 1'h1; // @[RegFile.scala 74:20:@53586.4]
  assign regs_276_clock = clock; // @[:@53595.4]
  assign regs_276_reset = io_reset; // @[:@53596.4 RegFile.scala 76:16:@53603.4]
  assign regs_276_io_in = 64'h0; // @[RegFile.scala 75:16:@53602.4]
  assign regs_276_io_reset = reset; // @[RegFile.scala 78:19:@53606.4]
  assign regs_276_io_enable = 1'h1; // @[RegFile.scala 74:20:@53600.4]
  assign regs_277_clock = clock; // @[:@53609.4]
  assign regs_277_reset = io_reset; // @[:@53610.4 RegFile.scala 76:16:@53617.4]
  assign regs_277_io_in = 64'h0; // @[RegFile.scala 75:16:@53616.4]
  assign regs_277_io_reset = reset; // @[RegFile.scala 78:19:@53620.4]
  assign regs_277_io_enable = 1'h1; // @[RegFile.scala 74:20:@53614.4]
  assign regs_278_clock = clock; // @[:@53623.4]
  assign regs_278_reset = io_reset; // @[:@53624.4 RegFile.scala 76:16:@53631.4]
  assign regs_278_io_in = 64'h0; // @[RegFile.scala 75:16:@53630.4]
  assign regs_278_io_reset = reset; // @[RegFile.scala 78:19:@53634.4]
  assign regs_278_io_enable = 1'h1; // @[RegFile.scala 74:20:@53628.4]
  assign regs_279_clock = clock; // @[:@53637.4]
  assign regs_279_reset = io_reset; // @[:@53638.4 RegFile.scala 76:16:@53645.4]
  assign regs_279_io_in = 64'h0; // @[RegFile.scala 75:16:@53644.4]
  assign regs_279_io_reset = reset; // @[RegFile.scala 78:19:@53648.4]
  assign regs_279_io_enable = 1'h1; // @[RegFile.scala 74:20:@53642.4]
  assign regs_280_clock = clock; // @[:@53651.4]
  assign regs_280_reset = io_reset; // @[:@53652.4 RegFile.scala 76:16:@53659.4]
  assign regs_280_io_in = 64'h0; // @[RegFile.scala 75:16:@53658.4]
  assign regs_280_io_reset = reset; // @[RegFile.scala 78:19:@53662.4]
  assign regs_280_io_enable = 1'h1; // @[RegFile.scala 74:20:@53656.4]
  assign regs_281_clock = clock; // @[:@53665.4]
  assign regs_281_reset = io_reset; // @[:@53666.4 RegFile.scala 76:16:@53673.4]
  assign regs_281_io_in = 64'h0; // @[RegFile.scala 75:16:@53672.4]
  assign regs_281_io_reset = reset; // @[RegFile.scala 78:19:@53676.4]
  assign regs_281_io_enable = 1'h1; // @[RegFile.scala 74:20:@53670.4]
  assign regs_282_clock = clock; // @[:@53679.4]
  assign regs_282_reset = io_reset; // @[:@53680.4 RegFile.scala 76:16:@53687.4]
  assign regs_282_io_in = 64'h0; // @[RegFile.scala 75:16:@53686.4]
  assign regs_282_io_reset = reset; // @[RegFile.scala 78:19:@53690.4]
  assign regs_282_io_enable = 1'h1; // @[RegFile.scala 74:20:@53684.4]
  assign regs_283_clock = clock; // @[:@53693.4]
  assign regs_283_reset = io_reset; // @[:@53694.4 RegFile.scala 76:16:@53701.4]
  assign regs_283_io_in = 64'h0; // @[RegFile.scala 75:16:@53700.4]
  assign regs_283_io_reset = reset; // @[RegFile.scala 78:19:@53704.4]
  assign regs_283_io_enable = 1'h1; // @[RegFile.scala 74:20:@53698.4]
  assign regs_284_clock = clock; // @[:@53707.4]
  assign regs_284_reset = io_reset; // @[:@53708.4 RegFile.scala 76:16:@53715.4]
  assign regs_284_io_in = 64'h0; // @[RegFile.scala 75:16:@53714.4]
  assign regs_284_io_reset = reset; // @[RegFile.scala 78:19:@53718.4]
  assign regs_284_io_enable = 1'h1; // @[RegFile.scala 74:20:@53712.4]
  assign regs_285_clock = clock; // @[:@53721.4]
  assign regs_285_reset = io_reset; // @[:@53722.4 RegFile.scala 76:16:@53729.4]
  assign regs_285_io_in = 64'h0; // @[RegFile.scala 75:16:@53728.4]
  assign regs_285_io_reset = reset; // @[RegFile.scala 78:19:@53732.4]
  assign regs_285_io_enable = 1'h1; // @[RegFile.scala 74:20:@53726.4]
  assign regs_286_clock = clock; // @[:@53735.4]
  assign regs_286_reset = io_reset; // @[:@53736.4 RegFile.scala 76:16:@53743.4]
  assign regs_286_io_in = 64'h0; // @[RegFile.scala 75:16:@53742.4]
  assign regs_286_io_reset = reset; // @[RegFile.scala 78:19:@53746.4]
  assign regs_286_io_enable = 1'h1; // @[RegFile.scala 74:20:@53740.4]
  assign regs_287_clock = clock; // @[:@53749.4]
  assign regs_287_reset = io_reset; // @[:@53750.4 RegFile.scala 76:16:@53757.4]
  assign regs_287_io_in = 64'h0; // @[RegFile.scala 75:16:@53756.4]
  assign regs_287_io_reset = reset; // @[RegFile.scala 78:19:@53760.4]
  assign regs_287_io_enable = 1'h1; // @[RegFile.scala 74:20:@53754.4]
  assign regs_288_clock = clock; // @[:@53763.4]
  assign regs_288_reset = io_reset; // @[:@53764.4 RegFile.scala 76:16:@53771.4]
  assign regs_288_io_in = 64'h0; // @[RegFile.scala 75:16:@53770.4]
  assign regs_288_io_reset = reset; // @[RegFile.scala 78:19:@53774.4]
  assign regs_288_io_enable = 1'h1; // @[RegFile.scala 74:20:@53768.4]
  assign regs_289_clock = clock; // @[:@53777.4]
  assign regs_289_reset = io_reset; // @[:@53778.4 RegFile.scala 76:16:@53785.4]
  assign regs_289_io_in = 64'h0; // @[RegFile.scala 75:16:@53784.4]
  assign regs_289_io_reset = reset; // @[RegFile.scala 78:19:@53788.4]
  assign regs_289_io_enable = 1'h1; // @[RegFile.scala 74:20:@53782.4]
  assign regs_290_clock = clock; // @[:@53791.4]
  assign regs_290_reset = io_reset; // @[:@53792.4 RegFile.scala 76:16:@53799.4]
  assign regs_290_io_in = 64'h0; // @[RegFile.scala 75:16:@53798.4]
  assign regs_290_io_reset = reset; // @[RegFile.scala 78:19:@53802.4]
  assign regs_290_io_enable = 1'h1; // @[RegFile.scala 74:20:@53796.4]
  assign regs_291_clock = clock; // @[:@53805.4]
  assign regs_291_reset = io_reset; // @[:@53806.4 RegFile.scala 76:16:@53813.4]
  assign regs_291_io_in = 64'h0; // @[RegFile.scala 75:16:@53812.4]
  assign regs_291_io_reset = reset; // @[RegFile.scala 78:19:@53816.4]
  assign regs_291_io_enable = 1'h1; // @[RegFile.scala 74:20:@53810.4]
  assign regs_292_clock = clock; // @[:@53819.4]
  assign regs_292_reset = io_reset; // @[:@53820.4 RegFile.scala 76:16:@53827.4]
  assign regs_292_io_in = 64'h0; // @[RegFile.scala 75:16:@53826.4]
  assign regs_292_io_reset = reset; // @[RegFile.scala 78:19:@53830.4]
  assign regs_292_io_enable = 1'h1; // @[RegFile.scala 74:20:@53824.4]
  assign regs_293_clock = clock; // @[:@53833.4]
  assign regs_293_reset = io_reset; // @[:@53834.4 RegFile.scala 76:16:@53841.4]
  assign regs_293_io_in = 64'h0; // @[RegFile.scala 75:16:@53840.4]
  assign regs_293_io_reset = reset; // @[RegFile.scala 78:19:@53844.4]
  assign regs_293_io_enable = 1'h1; // @[RegFile.scala 74:20:@53838.4]
  assign regs_294_clock = clock; // @[:@53847.4]
  assign regs_294_reset = io_reset; // @[:@53848.4 RegFile.scala 76:16:@53855.4]
  assign regs_294_io_in = 64'h0; // @[RegFile.scala 75:16:@53854.4]
  assign regs_294_io_reset = reset; // @[RegFile.scala 78:19:@53858.4]
  assign regs_294_io_enable = 1'h1; // @[RegFile.scala 74:20:@53852.4]
  assign regs_295_clock = clock; // @[:@53861.4]
  assign regs_295_reset = io_reset; // @[:@53862.4 RegFile.scala 76:16:@53869.4]
  assign regs_295_io_in = 64'h0; // @[RegFile.scala 75:16:@53868.4]
  assign regs_295_io_reset = reset; // @[RegFile.scala 78:19:@53872.4]
  assign regs_295_io_enable = 1'h1; // @[RegFile.scala 74:20:@53866.4]
  assign regs_296_clock = clock; // @[:@53875.4]
  assign regs_296_reset = io_reset; // @[:@53876.4 RegFile.scala 76:16:@53883.4]
  assign regs_296_io_in = 64'h0; // @[RegFile.scala 75:16:@53882.4]
  assign regs_296_io_reset = reset; // @[RegFile.scala 78:19:@53886.4]
  assign regs_296_io_enable = 1'h1; // @[RegFile.scala 74:20:@53880.4]
  assign regs_297_clock = clock; // @[:@53889.4]
  assign regs_297_reset = io_reset; // @[:@53890.4 RegFile.scala 76:16:@53897.4]
  assign regs_297_io_in = 64'h0; // @[RegFile.scala 75:16:@53896.4]
  assign regs_297_io_reset = reset; // @[RegFile.scala 78:19:@53900.4]
  assign regs_297_io_enable = 1'h1; // @[RegFile.scala 74:20:@53894.4]
  assign regs_298_clock = clock; // @[:@53903.4]
  assign regs_298_reset = io_reset; // @[:@53904.4 RegFile.scala 76:16:@53911.4]
  assign regs_298_io_in = 64'h0; // @[RegFile.scala 75:16:@53910.4]
  assign regs_298_io_reset = reset; // @[RegFile.scala 78:19:@53914.4]
  assign regs_298_io_enable = 1'h1; // @[RegFile.scala 74:20:@53908.4]
  assign regs_299_clock = clock; // @[:@53917.4]
  assign regs_299_reset = io_reset; // @[:@53918.4 RegFile.scala 76:16:@53925.4]
  assign regs_299_io_in = 64'h0; // @[RegFile.scala 75:16:@53924.4]
  assign regs_299_io_reset = reset; // @[RegFile.scala 78:19:@53928.4]
  assign regs_299_io_enable = 1'h1; // @[RegFile.scala 74:20:@53922.4]
  assign regs_300_clock = clock; // @[:@53931.4]
  assign regs_300_reset = io_reset; // @[:@53932.4 RegFile.scala 76:16:@53939.4]
  assign regs_300_io_in = 64'h0; // @[RegFile.scala 75:16:@53938.4]
  assign regs_300_io_reset = reset; // @[RegFile.scala 78:19:@53942.4]
  assign regs_300_io_enable = 1'h1; // @[RegFile.scala 74:20:@53936.4]
  assign regs_301_clock = clock; // @[:@53945.4]
  assign regs_301_reset = io_reset; // @[:@53946.4 RegFile.scala 76:16:@53953.4]
  assign regs_301_io_in = 64'h0; // @[RegFile.scala 75:16:@53952.4]
  assign regs_301_io_reset = reset; // @[RegFile.scala 78:19:@53956.4]
  assign regs_301_io_enable = 1'h1; // @[RegFile.scala 74:20:@53950.4]
  assign regs_302_clock = clock; // @[:@53959.4]
  assign regs_302_reset = io_reset; // @[:@53960.4 RegFile.scala 76:16:@53967.4]
  assign regs_302_io_in = 64'h0; // @[RegFile.scala 75:16:@53966.4]
  assign regs_302_io_reset = reset; // @[RegFile.scala 78:19:@53970.4]
  assign regs_302_io_enable = 1'h1; // @[RegFile.scala 74:20:@53964.4]
  assign regs_303_clock = clock; // @[:@53973.4]
  assign regs_303_reset = io_reset; // @[:@53974.4 RegFile.scala 76:16:@53981.4]
  assign regs_303_io_in = 64'h0; // @[RegFile.scala 75:16:@53980.4]
  assign regs_303_io_reset = reset; // @[RegFile.scala 78:19:@53984.4]
  assign regs_303_io_enable = 1'h1; // @[RegFile.scala 74:20:@53978.4]
  assign regs_304_clock = clock; // @[:@53987.4]
  assign regs_304_reset = io_reset; // @[:@53988.4 RegFile.scala 76:16:@53995.4]
  assign regs_304_io_in = 64'h0; // @[RegFile.scala 75:16:@53994.4]
  assign regs_304_io_reset = reset; // @[RegFile.scala 78:19:@53998.4]
  assign regs_304_io_enable = 1'h1; // @[RegFile.scala 74:20:@53992.4]
  assign regs_305_clock = clock; // @[:@54001.4]
  assign regs_305_reset = io_reset; // @[:@54002.4 RegFile.scala 76:16:@54009.4]
  assign regs_305_io_in = 64'h0; // @[RegFile.scala 75:16:@54008.4]
  assign regs_305_io_reset = reset; // @[RegFile.scala 78:19:@54012.4]
  assign regs_305_io_enable = 1'h1; // @[RegFile.scala 74:20:@54006.4]
  assign regs_306_clock = clock; // @[:@54015.4]
  assign regs_306_reset = io_reset; // @[:@54016.4 RegFile.scala 76:16:@54023.4]
  assign regs_306_io_in = 64'h0; // @[RegFile.scala 75:16:@54022.4]
  assign regs_306_io_reset = reset; // @[RegFile.scala 78:19:@54026.4]
  assign regs_306_io_enable = 1'h1; // @[RegFile.scala 74:20:@54020.4]
  assign regs_307_clock = clock; // @[:@54029.4]
  assign regs_307_reset = io_reset; // @[:@54030.4 RegFile.scala 76:16:@54037.4]
  assign regs_307_io_in = 64'h0; // @[RegFile.scala 75:16:@54036.4]
  assign regs_307_io_reset = reset; // @[RegFile.scala 78:19:@54040.4]
  assign regs_307_io_enable = 1'h1; // @[RegFile.scala 74:20:@54034.4]
  assign regs_308_clock = clock; // @[:@54043.4]
  assign regs_308_reset = io_reset; // @[:@54044.4 RegFile.scala 76:16:@54051.4]
  assign regs_308_io_in = 64'h0; // @[RegFile.scala 75:16:@54050.4]
  assign regs_308_io_reset = reset; // @[RegFile.scala 78:19:@54054.4]
  assign regs_308_io_enable = 1'h1; // @[RegFile.scala 74:20:@54048.4]
  assign regs_309_clock = clock; // @[:@54057.4]
  assign regs_309_reset = io_reset; // @[:@54058.4 RegFile.scala 76:16:@54065.4]
  assign regs_309_io_in = 64'h0; // @[RegFile.scala 75:16:@54064.4]
  assign regs_309_io_reset = reset; // @[RegFile.scala 78:19:@54068.4]
  assign regs_309_io_enable = 1'h1; // @[RegFile.scala 74:20:@54062.4]
  assign regs_310_clock = clock; // @[:@54071.4]
  assign regs_310_reset = io_reset; // @[:@54072.4 RegFile.scala 76:16:@54079.4]
  assign regs_310_io_in = 64'h0; // @[RegFile.scala 75:16:@54078.4]
  assign regs_310_io_reset = reset; // @[RegFile.scala 78:19:@54082.4]
  assign regs_310_io_enable = 1'h1; // @[RegFile.scala 74:20:@54076.4]
  assign regs_311_clock = clock; // @[:@54085.4]
  assign regs_311_reset = io_reset; // @[:@54086.4 RegFile.scala 76:16:@54093.4]
  assign regs_311_io_in = 64'h0; // @[RegFile.scala 75:16:@54092.4]
  assign regs_311_io_reset = reset; // @[RegFile.scala 78:19:@54096.4]
  assign regs_311_io_enable = 1'h1; // @[RegFile.scala 74:20:@54090.4]
  assign regs_312_clock = clock; // @[:@54099.4]
  assign regs_312_reset = io_reset; // @[:@54100.4 RegFile.scala 76:16:@54107.4]
  assign regs_312_io_in = 64'h0; // @[RegFile.scala 75:16:@54106.4]
  assign regs_312_io_reset = reset; // @[RegFile.scala 78:19:@54110.4]
  assign regs_312_io_enable = 1'h1; // @[RegFile.scala 74:20:@54104.4]
  assign regs_313_clock = clock; // @[:@54113.4]
  assign regs_313_reset = io_reset; // @[:@54114.4 RegFile.scala 76:16:@54121.4]
  assign regs_313_io_in = 64'h0; // @[RegFile.scala 75:16:@54120.4]
  assign regs_313_io_reset = reset; // @[RegFile.scala 78:19:@54124.4]
  assign regs_313_io_enable = 1'h1; // @[RegFile.scala 74:20:@54118.4]
  assign regs_314_clock = clock; // @[:@54127.4]
  assign regs_314_reset = io_reset; // @[:@54128.4 RegFile.scala 76:16:@54135.4]
  assign regs_314_io_in = 64'h0; // @[RegFile.scala 75:16:@54134.4]
  assign regs_314_io_reset = reset; // @[RegFile.scala 78:19:@54138.4]
  assign regs_314_io_enable = 1'h1; // @[RegFile.scala 74:20:@54132.4]
  assign regs_315_clock = clock; // @[:@54141.4]
  assign regs_315_reset = io_reset; // @[:@54142.4 RegFile.scala 76:16:@54149.4]
  assign regs_315_io_in = 64'h0; // @[RegFile.scala 75:16:@54148.4]
  assign regs_315_io_reset = reset; // @[RegFile.scala 78:19:@54152.4]
  assign regs_315_io_enable = 1'h1; // @[RegFile.scala 74:20:@54146.4]
  assign regs_316_clock = clock; // @[:@54155.4]
  assign regs_316_reset = io_reset; // @[:@54156.4 RegFile.scala 76:16:@54163.4]
  assign regs_316_io_in = 64'h0; // @[RegFile.scala 75:16:@54162.4]
  assign regs_316_io_reset = reset; // @[RegFile.scala 78:19:@54166.4]
  assign regs_316_io_enable = 1'h1; // @[RegFile.scala 74:20:@54160.4]
  assign regs_317_clock = clock; // @[:@54169.4]
  assign regs_317_reset = io_reset; // @[:@54170.4 RegFile.scala 76:16:@54177.4]
  assign regs_317_io_in = 64'h0; // @[RegFile.scala 75:16:@54176.4]
  assign regs_317_io_reset = reset; // @[RegFile.scala 78:19:@54180.4]
  assign regs_317_io_enable = 1'h1; // @[RegFile.scala 74:20:@54174.4]
  assign regs_318_clock = clock; // @[:@54183.4]
  assign regs_318_reset = io_reset; // @[:@54184.4 RegFile.scala 76:16:@54191.4]
  assign regs_318_io_in = 64'h0; // @[RegFile.scala 75:16:@54190.4]
  assign regs_318_io_reset = reset; // @[RegFile.scala 78:19:@54194.4]
  assign regs_318_io_enable = 1'h1; // @[RegFile.scala 74:20:@54188.4]
  assign regs_319_clock = clock; // @[:@54197.4]
  assign regs_319_reset = io_reset; // @[:@54198.4 RegFile.scala 76:16:@54205.4]
  assign regs_319_io_in = 64'h0; // @[RegFile.scala 75:16:@54204.4]
  assign regs_319_io_reset = reset; // @[RegFile.scala 78:19:@54208.4]
  assign regs_319_io_enable = 1'h1; // @[RegFile.scala 74:20:@54202.4]
  assign regs_320_clock = clock; // @[:@54211.4]
  assign regs_320_reset = io_reset; // @[:@54212.4 RegFile.scala 76:16:@54219.4]
  assign regs_320_io_in = 64'h0; // @[RegFile.scala 75:16:@54218.4]
  assign regs_320_io_reset = reset; // @[RegFile.scala 78:19:@54222.4]
  assign regs_320_io_enable = 1'h1; // @[RegFile.scala 74:20:@54216.4]
  assign regs_321_clock = clock; // @[:@54225.4]
  assign regs_321_reset = io_reset; // @[:@54226.4 RegFile.scala 76:16:@54233.4]
  assign regs_321_io_in = 64'h0; // @[RegFile.scala 75:16:@54232.4]
  assign regs_321_io_reset = reset; // @[RegFile.scala 78:19:@54236.4]
  assign regs_321_io_enable = 1'h1; // @[RegFile.scala 74:20:@54230.4]
  assign regs_322_clock = clock; // @[:@54239.4]
  assign regs_322_reset = io_reset; // @[:@54240.4 RegFile.scala 76:16:@54247.4]
  assign regs_322_io_in = 64'h0; // @[RegFile.scala 75:16:@54246.4]
  assign regs_322_io_reset = reset; // @[RegFile.scala 78:19:@54250.4]
  assign regs_322_io_enable = 1'h1; // @[RegFile.scala 74:20:@54244.4]
  assign regs_323_clock = clock; // @[:@54253.4]
  assign regs_323_reset = io_reset; // @[:@54254.4 RegFile.scala 76:16:@54261.4]
  assign regs_323_io_in = 64'h0; // @[RegFile.scala 75:16:@54260.4]
  assign regs_323_io_reset = reset; // @[RegFile.scala 78:19:@54264.4]
  assign regs_323_io_enable = 1'h1; // @[RegFile.scala 74:20:@54258.4]
  assign regs_324_clock = clock; // @[:@54267.4]
  assign regs_324_reset = io_reset; // @[:@54268.4 RegFile.scala 76:16:@54275.4]
  assign regs_324_io_in = 64'h0; // @[RegFile.scala 75:16:@54274.4]
  assign regs_324_io_reset = reset; // @[RegFile.scala 78:19:@54278.4]
  assign regs_324_io_enable = 1'h1; // @[RegFile.scala 74:20:@54272.4]
  assign regs_325_clock = clock; // @[:@54281.4]
  assign regs_325_reset = io_reset; // @[:@54282.4 RegFile.scala 76:16:@54289.4]
  assign regs_325_io_in = 64'h0; // @[RegFile.scala 75:16:@54288.4]
  assign regs_325_io_reset = reset; // @[RegFile.scala 78:19:@54292.4]
  assign regs_325_io_enable = 1'h1; // @[RegFile.scala 74:20:@54286.4]
  assign regs_326_clock = clock; // @[:@54295.4]
  assign regs_326_reset = io_reset; // @[:@54296.4 RegFile.scala 76:16:@54303.4]
  assign regs_326_io_in = 64'h0; // @[RegFile.scala 75:16:@54302.4]
  assign regs_326_io_reset = reset; // @[RegFile.scala 78:19:@54306.4]
  assign regs_326_io_enable = 1'h1; // @[RegFile.scala 74:20:@54300.4]
  assign regs_327_clock = clock; // @[:@54309.4]
  assign regs_327_reset = io_reset; // @[:@54310.4 RegFile.scala 76:16:@54317.4]
  assign regs_327_io_in = 64'h0; // @[RegFile.scala 75:16:@54316.4]
  assign regs_327_io_reset = reset; // @[RegFile.scala 78:19:@54320.4]
  assign regs_327_io_enable = 1'h1; // @[RegFile.scala 74:20:@54314.4]
  assign regs_328_clock = clock; // @[:@54323.4]
  assign regs_328_reset = io_reset; // @[:@54324.4 RegFile.scala 76:16:@54331.4]
  assign regs_328_io_in = 64'h0; // @[RegFile.scala 75:16:@54330.4]
  assign regs_328_io_reset = reset; // @[RegFile.scala 78:19:@54334.4]
  assign regs_328_io_enable = 1'h1; // @[RegFile.scala 74:20:@54328.4]
  assign regs_329_clock = clock; // @[:@54337.4]
  assign regs_329_reset = io_reset; // @[:@54338.4 RegFile.scala 76:16:@54345.4]
  assign regs_329_io_in = 64'h0; // @[RegFile.scala 75:16:@54344.4]
  assign regs_329_io_reset = reset; // @[RegFile.scala 78:19:@54348.4]
  assign regs_329_io_enable = 1'h1; // @[RegFile.scala 74:20:@54342.4]
  assign regs_330_clock = clock; // @[:@54351.4]
  assign regs_330_reset = io_reset; // @[:@54352.4 RegFile.scala 76:16:@54359.4]
  assign regs_330_io_in = 64'h0; // @[RegFile.scala 75:16:@54358.4]
  assign regs_330_io_reset = reset; // @[RegFile.scala 78:19:@54362.4]
  assign regs_330_io_enable = 1'h1; // @[RegFile.scala 74:20:@54356.4]
  assign regs_331_clock = clock; // @[:@54365.4]
  assign regs_331_reset = io_reset; // @[:@54366.4 RegFile.scala 76:16:@54373.4]
  assign regs_331_io_in = 64'h0; // @[RegFile.scala 75:16:@54372.4]
  assign regs_331_io_reset = reset; // @[RegFile.scala 78:19:@54376.4]
  assign regs_331_io_enable = 1'h1; // @[RegFile.scala 74:20:@54370.4]
  assign regs_332_clock = clock; // @[:@54379.4]
  assign regs_332_reset = io_reset; // @[:@54380.4 RegFile.scala 76:16:@54387.4]
  assign regs_332_io_in = 64'h0; // @[RegFile.scala 75:16:@54386.4]
  assign regs_332_io_reset = reset; // @[RegFile.scala 78:19:@54390.4]
  assign regs_332_io_enable = 1'h1; // @[RegFile.scala 74:20:@54384.4]
  assign regs_333_clock = clock; // @[:@54393.4]
  assign regs_333_reset = io_reset; // @[:@54394.4 RegFile.scala 76:16:@54401.4]
  assign regs_333_io_in = 64'h0; // @[RegFile.scala 75:16:@54400.4]
  assign regs_333_io_reset = reset; // @[RegFile.scala 78:19:@54404.4]
  assign regs_333_io_enable = 1'h1; // @[RegFile.scala 74:20:@54398.4]
  assign regs_334_clock = clock; // @[:@54407.4]
  assign regs_334_reset = io_reset; // @[:@54408.4 RegFile.scala 76:16:@54415.4]
  assign regs_334_io_in = 64'h0; // @[RegFile.scala 75:16:@54414.4]
  assign regs_334_io_reset = reset; // @[RegFile.scala 78:19:@54418.4]
  assign regs_334_io_enable = 1'h1; // @[RegFile.scala 74:20:@54412.4]
  assign regs_335_clock = clock; // @[:@54421.4]
  assign regs_335_reset = io_reset; // @[:@54422.4 RegFile.scala 76:16:@54429.4]
  assign regs_335_io_in = 64'h0; // @[RegFile.scala 75:16:@54428.4]
  assign regs_335_io_reset = reset; // @[RegFile.scala 78:19:@54432.4]
  assign regs_335_io_enable = 1'h1; // @[RegFile.scala 74:20:@54426.4]
  assign regs_336_clock = clock; // @[:@54435.4]
  assign regs_336_reset = io_reset; // @[:@54436.4 RegFile.scala 76:16:@54443.4]
  assign regs_336_io_in = 64'h0; // @[RegFile.scala 75:16:@54442.4]
  assign regs_336_io_reset = reset; // @[RegFile.scala 78:19:@54446.4]
  assign regs_336_io_enable = 1'h1; // @[RegFile.scala 74:20:@54440.4]
  assign regs_337_clock = clock; // @[:@54449.4]
  assign regs_337_reset = io_reset; // @[:@54450.4 RegFile.scala 76:16:@54457.4]
  assign regs_337_io_in = 64'h0; // @[RegFile.scala 75:16:@54456.4]
  assign regs_337_io_reset = reset; // @[RegFile.scala 78:19:@54460.4]
  assign regs_337_io_enable = 1'h1; // @[RegFile.scala 74:20:@54454.4]
  assign regs_338_clock = clock; // @[:@54463.4]
  assign regs_338_reset = io_reset; // @[:@54464.4 RegFile.scala 76:16:@54471.4]
  assign regs_338_io_in = 64'h0; // @[RegFile.scala 75:16:@54470.4]
  assign regs_338_io_reset = reset; // @[RegFile.scala 78:19:@54474.4]
  assign regs_338_io_enable = 1'h1; // @[RegFile.scala 74:20:@54468.4]
  assign regs_339_clock = clock; // @[:@54477.4]
  assign regs_339_reset = io_reset; // @[:@54478.4 RegFile.scala 76:16:@54485.4]
  assign regs_339_io_in = 64'h0; // @[RegFile.scala 75:16:@54484.4]
  assign regs_339_io_reset = reset; // @[RegFile.scala 78:19:@54488.4]
  assign regs_339_io_enable = 1'h1; // @[RegFile.scala 74:20:@54482.4]
  assign regs_340_clock = clock; // @[:@54491.4]
  assign regs_340_reset = io_reset; // @[:@54492.4 RegFile.scala 76:16:@54499.4]
  assign regs_340_io_in = 64'h0; // @[RegFile.scala 75:16:@54498.4]
  assign regs_340_io_reset = reset; // @[RegFile.scala 78:19:@54502.4]
  assign regs_340_io_enable = 1'h1; // @[RegFile.scala 74:20:@54496.4]
  assign regs_341_clock = clock; // @[:@54505.4]
  assign regs_341_reset = io_reset; // @[:@54506.4 RegFile.scala 76:16:@54513.4]
  assign regs_341_io_in = 64'h0; // @[RegFile.scala 75:16:@54512.4]
  assign regs_341_io_reset = reset; // @[RegFile.scala 78:19:@54516.4]
  assign regs_341_io_enable = 1'h1; // @[RegFile.scala 74:20:@54510.4]
  assign regs_342_clock = clock; // @[:@54519.4]
  assign regs_342_reset = io_reset; // @[:@54520.4 RegFile.scala 76:16:@54527.4]
  assign regs_342_io_in = 64'h0; // @[RegFile.scala 75:16:@54526.4]
  assign regs_342_io_reset = reset; // @[RegFile.scala 78:19:@54530.4]
  assign regs_342_io_enable = 1'h1; // @[RegFile.scala 74:20:@54524.4]
  assign regs_343_clock = clock; // @[:@54533.4]
  assign regs_343_reset = io_reset; // @[:@54534.4 RegFile.scala 76:16:@54541.4]
  assign regs_343_io_in = 64'h0; // @[RegFile.scala 75:16:@54540.4]
  assign regs_343_io_reset = reset; // @[RegFile.scala 78:19:@54544.4]
  assign regs_343_io_enable = 1'h1; // @[RegFile.scala 74:20:@54538.4]
  assign regs_344_clock = clock; // @[:@54547.4]
  assign regs_344_reset = io_reset; // @[:@54548.4 RegFile.scala 76:16:@54555.4]
  assign regs_344_io_in = 64'h0; // @[RegFile.scala 75:16:@54554.4]
  assign regs_344_io_reset = reset; // @[RegFile.scala 78:19:@54558.4]
  assign regs_344_io_enable = 1'h1; // @[RegFile.scala 74:20:@54552.4]
  assign regs_345_clock = clock; // @[:@54561.4]
  assign regs_345_reset = io_reset; // @[:@54562.4 RegFile.scala 76:16:@54569.4]
  assign regs_345_io_in = 64'h0; // @[RegFile.scala 75:16:@54568.4]
  assign regs_345_io_reset = reset; // @[RegFile.scala 78:19:@54572.4]
  assign regs_345_io_enable = 1'h1; // @[RegFile.scala 74:20:@54566.4]
  assign regs_346_clock = clock; // @[:@54575.4]
  assign regs_346_reset = io_reset; // @[:@54576.4 RegFile.scala 76:16:@54583.4]
  assign regs_346_io_in = 64'h0; // @[RegFile.scala 75:16:@54582.4]
  assign regs_346_io_reset = reset; // @[RegFile.scala 78:19:@54586.4]
  assign regs_346_io_enable = 1'h1; // @[RegFile.scala 74:20:@54580.4]
  assign regs_347_clock = clock; // @[:@54589.4]
  assign regs_347_reset = io_reset; // @[:@54590.4 RegFile.scala 76:16:@54597.4]
  assign regs_347_io_in = 64'h0; // @[RegFile.scala 75:16:@54596.4]
  assign regs_347_io_reset = reset; // @[RegFile.scala 78:19:@54600.4]
  assign regs_347_io_enable = 1'h1; // @[RegFile.scala 74:20:@54594.4]
  assign regs_348_clock = clock; // @[:@54603.4]
  assign regs_348_reset = io_reset; // @[:@54604.4 RegFile.scala 76:16:@54611.4]
  assign regs_348_io_in = 64'h0; // @[RegFile.scala 75:16:@54610.4]
  assign regs_348_io_reset = reset; // @[RegFile.scala 78:19:@54614.4]
  assign regs_348_io_enable = 1'h1; // @[RegFile.scala 74:20:@54608.4]
  assign regs_349_clock = clock; // @[:@54617.4]
  assign regs_349_reset = io_reset; // @[:@54618.4 RegFile.scala 76:16:@54625.4]
  assign regs_349_io_in = 64'h0; // @[RegFile.scala 75:16:@54624.4]
  assign regs_349_io_reset = reset; // @[RegFile.scala 78:19:@54628.4]
  assign regs_349_io_enable = 1'h1; // @[RegFile.scala 74:20:@54622.4]
  assign regs_350_clock = clock; // @[:@54631.4]
  assign regs_350_reset = io_reset; // @[:@54632.4 RegFile.scala 76:16:@54639.4]
  assign regs_350_io_in = 64'h0; // @[RegFile.scala 75:16:@54638.4]
  assign regs_350_io_reset = reset; // @[RegFile.scala 78:19:@54642.4]
  assign regs_350_io_enable = 1'h1; // @[RegFile.scala 74:20:@54636.4]
  assign regs_351_clock = clock; // @[:@54645.4]
  assign regs_351_reset = io_reset; // @[:@54646.4 RegFile.scala 76:16:@54653.4]
  assign regs_351_io_in = 64'h0; // @[RegFile.scala 75:16:@54652.4]
  assign regs_351_io_reset = reset; // @[RegFile.scala 78:19:@54656.4]
  assign regs_351_io_enable = 1'h1; // @[RegFile.scala 74:20:@54650.4]
  assign regs_352_clock = clock; // @[:@54659.4]
  assign regs_352_reset = io_reset; // @[:@54660.4 RegFile.scala 76:16:@54667.4]
  assign regs_352_io_in = 64'h0; // @[RegFile.scala 75:16:@54666.4]
  assign regs_352_io_reset = reset; // @[RegFile.scala 78:19:@54670.4]
  assign regs_352_io_enable = 1'h1; // @[RegFile.scala 74:20:@54664.4]
  assign regs_353_clock = clock; // @[:@54673.4]
  assign regs_353_reset = io_reset; // @[:@54674.4 RegFile.scala 76:16:@54681.4]
  assign regs_353_io_in = 64'h0; // @[RegFile.scala 75:16:@54680.4]
  assign regs_353_io_reset = reset; // @[RegFile.scala 78:19:@54684.4]
  assign regs_353_io_enable = 1'h1; // @[RegFile.scala 74:20:@54678.4]
  assign regs_354_clock = clock; // @[:@54687.4]
  assign regs_354_reset = io_reset; // @[:@54688.4 RegFile.scala 76:16:@54695.4]
  assign regs_354_io_in = 64'h0; // @[RegFile.scala 75:16:@54694.4]
  assign regs_354_io_reset = reset; // @[RegFile.scala 78:19:@54698.4]
  assign regs_354_io_enable = 1'h1; // @[RegFile.scala 74:20:@54692.4]
  assign regs_355_clock = clock; // @[:@54701.4]
  assign regs_355_reset = io_reset; // @[:@54702.4 RegFile.scala 76:16:@54709.4]
  assign regs_355_io_in = 64'h0; // @[RegFile.scala 75:16:@54708.4]
  assign regs_355_io_reset = reset; // @[RegFile.scala 78:19:@54712.4]
  assign regs_355_io_enable = 1'h1; // @[RegFile.scala 74:20:@54706.4]
  assign regs_356_clock = clock; // @[:@54715.4]
  assign regs_356_reset = io_reset; // @[:@54716.4 RegFile.scala 76:16:@54723.4]
  assign regs_356_io_in = 64'h0; // @[RegFile.scala 75:16:@54722.4]
  assign regs_356_io_reset = reset; // @[RegFile.scala 78:19:@54726.4]
  assign regs_356_io_enable = 1'h1; // @[RegFile.scala 74:20:@54720.4]
  assign regs_357_clock = clock; // @[:@54729.4]
  assign regs_357_reset = io_reset; // @[:@54730.4 RegFile.scala 76:16:@54737.4]
  assign regs_357_io_in = 64'h0; // @[RegFile.scala 75:16:@54736.4]
  assign regs_357_io_reset = reset; // @[RegFile.scala 78:19:@54740.4]
  assign regs_357_io_enable = 1'h1; // @[RegFile.scala 74:20:@54734.4]
  assign regs_358_clock = clock; // @[:@54743.4]
  assign regs_358_reset = io_reset; // @[:@54744.4 RegFile.scala 76:16:@54751.4]
  assign regs_358_io_in = 64'h0; // @[RegFile.scala 75:16:@54750.4]
  assign regs_358_io_reset = reset; // @[RegFile.scala 78:19:@54754.4]
  assign regs_358_io_enable = 1'h1; // @[RegFile.scala 74:20:@54748.4]
  assign regs_359_clock = clock; // @[:@54757.4]
  assign regs_359_reset = io_reset; // @[:@54758.4 RegFile.scala 76:16:@54765.4]
  assign regs_359_io_in = 64'h0; // @[RegFile.scala 75:16:@54764.4]
  assign regs_359_io_reset = reset; // @[RegFile.scala 78:19:@54768.4]
  assign regs_359_io_enable = 1'h1; // @[RegFile.scala 74:20:@54762.4]
  assign regs_360_clock = clock; // @[:@54771.4]
  assign regs_360_reset = io_reset; // @[:@54772.4 RegFile.scala 76:16:@54779.4]
  assign regs_360_io_in = 64'h0; // @[RegFile.scala 75:16:@54778.4]
  assign regs_360_io_reset = reset; // @[RegFile.scala 78:19:@54782.4]
  assign regs_360_io_enable = 1'h1; // @[RegFile.scala 74:20:@54776.4]
  assign regs_361_clock = clock; // @[:@54785.4]
  assign regs_361_reset = io_reset; // @[:@54786.4 RegFile.scala 76:16:@54793.4]
  assign regs_361_io_in = 64'h0; // @[RegFile.scala 75:16:@54792.4]
  assign regs_361_io_reset = reset; // @[RegFile.scala 78:19:@54796.4]
  assign regs_361_io_enable = 1'h1; // @[RegFile.scala 74:20:@54790.4]
  assign regs_362_clock = clock; // @[:@54799.4]
  assign regs_362_reset = io_reset; // @[:@54800.4 RegFile.scala 76:16:@54807.4]
  assign regs_362_io_in = 64'h0; // @[RegFile.scala 75:16:@54806.4]
  assign regs_362_io_reset = reset; // @[RegFile.scala 78:19:@54810.4]
  assign regs_362_io_enable = 1'h1; // @[RegFile.scala 74:20:@54804.4]
  assign regs_363_clock = clock; // @[:@54813.4]
  assign regs_363_reset = io_reset; // @[:@54814.4 RegFile.scala 76:16:@54821.4]
  assign regs_363_io_in = 64'h0; // @[RegFile.scala 75:16:@54820.4]
  assign regs_363_io_reset = reset; // @[RegFile.scala 78:19:@54824.4]
  assign regs_363_io_enable = 1'h1; // @[RegFile.scala 74:20:@54818.4]
  assign regs_364_clock = clock; // @[:@54827.4]
  assign regs_364_reset = io_reset; // @[:@54828.4 RegFile.scala 76:16:@54835.4]
  assign regs_364_io_in = 64'h0; // @[RegFile.scala 75:16:@54834.4]
  assign regs_364_io_reset = reset; // @[RegFile.scala 78:19:@54838.4]
  assign regs_364_io_enable = 1'h1; // @[RegFile.scala 74:20:@54832.4]
  assign regs_365_clock = clock; // @[:@54841.4]
  assign regs_365_reset = io_reset; // @[:@54842.4 RegFile.scala 76:16:@54849.4]
  assign regs_365_io_in = 64'h0; // @[RegFile.scala 75:16:@54848.4]
  assign regs_365_io_reset = reset; // @[RegFile.scala 78:19:@54852.4]
  assign regs_365_io_enable = 1'h1; // @[RegFile.scala 74:20:@54846.4]
  assign regs_366_clock = clock; // @[:@54855.4]
  assign regs_366_reset = io_reset; // @[:@54856.4 RegFile.scala 76:16:@54863.4]
  assign regs_366_io_in = 64'h0; // @[RegFile.scala 75:16:@54862.4]
  assign regs_366_io_reset = reset; // @[RegFile.scala 78:19:@54866.4]
  assign regs_366_io_enable = 1'h1; // @[RegFile.scala 74:20:@54860.4]
  assign regs_367_clock = clock; // @[:@54869.4]
  assign regs_367_reset = io_reset; // @[:@54870.4 RegFile.scala 76:16:@54877.4]
  assign regs_367_io_in = 64'h0; // @[RegFile.scala 75:16:@54876.4]
  assign regs_367_io_reset = reset; // @[RegFile.scala 78:19:@54880.4]
  assign regs_367_io_enable = 1'h1; // @[RegFile.scala 74:20:@54874.4]
  assign regs_368_clock = clock; // @[:@54883.4]
  assign regs_368_reset = io_reset; // @[:@54884.4 RegFile.scala 76:16:@54891.4]
  assign regs_368_io_in = 64'h0; // @[RegFile.scala 75:16:@54890.4]
  assign regs_368_io_reset = reset; // @[RegFile.scala 78:19:@54894.4]
  assign regs_368_io_enable = 1'h1; // @[RegFile.scala 74:20:@54888.4]
  assign regs_369_clock = clock; // @[:@54897.4]
  assign regs_369_reset = io_reset; // @[:@54898.4 RegFile.scala 76:16:@54905.4]
  assign regs_369_io_in = 64'h0; // @[RegFile.scala 75:16:@54904.4]
  assign regs_369_io_reset = reset; // @[RegFile.scala 78:19:@54908.4]
  assign regs_369_io_enable = 1'h1; // @[RegFile.scala 74:20:@54902.4]
  assign regs_370_clock = clock; // @[:@54911.4]
  assign regs_370_reset = io_reset; // @[:@54912.4 RegFile.scala 76:16:@54919.4]
  assign regs_370_io_in = 64'h0; // @[RegFile.scala 75:16:@54918.4]
  assign regs_370_io_reset = reset; // @[RegFile.scala 78:19:@54922.4]
  assign regs_370_io_enable = 1'h1; // @[RegFile.scala 74:20:@54916.4]
  assign regs_371_clock = clock; // @[:@54925.4]
  assign regs_371_reset = io_reset; // @[:@54926.4 RegFile.scala 76:16:@54933.4]
  assign regs_371_io_in = 64'h0; // @[RegFile.scala 75:16:@54932.4]
  assign regs_371_io_reset = reset; // @[RegFile.scala 78:19:@54936.4]
  assign regs_371_io_enable = 1'h1; // @[RegFile.scala 74:20:@54930.4]
  assign regs_372_clock = clock; // @[:@54939.4]
  assign regs_372_reset = io_reset; // @[:@54940.4 RegFile.scala 76:16:@54947.4]
  assign regs_372_io_in = 64'h0; // @[RegFile.scala 75:16:@54946.4]
  assign regs_372_io_reset = reset; // @[RegFile.scala 78:19:@54950.4]
  assign regs_372_io_enable = 1'h1; // @[RegFile.scala 74:20:@54944.4]
  assign regs_373_clock = clock; // @[:@54953.4]
  assign regs_373_reset = io_reset; // @[:@54954.4 RegFile.scala 76:16:@54961.4]
  assign regs_373_io_in = 64'h0; // @[RegFile.scala 75:16:@54960.4]
  assign regs_373_io_reset = reset; // @[RegFile.scala 78:19:@54964.4]
  assign regs_373_io_enable = 1'h1; // @[RegFile.scala 74:20:@54958.4]
  assign regs_374_clock = clock; // @[:@54967.4]
  assign regs_374_reset = io_reset; // @[:@54968.4 RegFile.scala 76:16:@54975.4]
  assign regs_374_io_in = 64'h0; // @[RegFile.scala 75:16:@54974.4]
  assign regs_374_io_reset = reset; // @[RegFile.scala 78:19:@54978.4]
  assign regs_374_io_enable = 1'h1; // @[RegFile.scala 74:20:@54972.4]
  assign regs_375_clock = clock; // @[:@54981.4]
  assign regs_375_reset = io_reset; // @[:@54982.4 RegFile.scala 76:16:@54989.4]
  assign regs_375_io_in = 64'h0; // @[RegFile.scala 75:16:@54988.4]
  assign regs_375_io_reset = reset; // @[RegFile.scala 78:19:@54992.4]
  assign regs_375_io_enable = 1'h1; // @[RegFile.scala 74:20:@54986.4]
  assign regs_376_clock = clock; // @[:@54995.4]
  assign regs_376_reset = io_reset; // @[:@54996.4 RegFile.scala 76:16:@55003.4]
  assign regs_376_io_in = 64'h0; // @[RegFile.scala 75:16:@55002.4]
  assign regs_376_io_reset = reset; // @[RegFile.scala 78:19:@55006.4]
  assign regs_376_io_enable = 1'h1; // @[RegFile.scala 74:20:@55000.4]
  assign regs_377_clock = clock; // @[:@55009.4]
  assign regs_377_reset = io_reset; // @[:@55010.4 RegFile.scala 76:16:@55017.4]
  assign regs_377_io_in = 64'h0; // @[RegFile.scala 75:16:@55016.4]
  assign regs_377_io_reset = reset; // @[RegFile.scala 78:19:@55020.4]
  assign regs_377_io_enable = 1'h1; // @[RegFile.scala 74:20:@55014.4]
  assign regs_378_clock = clock; // @[:@55023.4]
  assign regs_378_reset = io_reset; // @[:@55024.4 RegFile.scala 76:16:@55031.4]
  assign regs_378_io_in = 64'h0; // @[RegFile.scala 75:16:@55030.4]
  assign regs_378_io_reset = reset; // @[RegFile.scala 78:19:@55034.4]
  assign regs_378_io_enable = 1'h1; // @[RegFile.scala 74:20:@55028.4]
  assign regs_379_clock = clock; // @[:@55037.4]
  assign regs_379_reset = io_reset; // @[:@55038.4 RegFile.scala 76:16:@55045.4]
  assign regs_379_io_in = 64'h0; // @[RegFile.scala 75:16:@55044.4]
  assign regs_379_io_reset = reset; // @[RegFile.scala 78:19:@55048.4]
  assign regs_379_io_enable = 1'h1; // @[RegFile.scala 74:20:@55042.4]
  assign regs_380_clock = clock; // @[:@55051.4]
  assign regs_380_reset = io_reset; // @[:@55052.4 RegFile.scala 76:16:@55059.4]
  assign regs_380_io_in = 64'h0; // @[RegFile.scala 75:16:@55058.4]
  assign regs_380_io_reset = reset; // @[RegFile.scala 78:19:@55062.4]
  assign regs_380_io_enable = 1'h1; // @[RegFile.scala 74:20:@55056.4]
  assign regs_381_clock = clock; // @[:@55065.4]
  assign regs_381_reset = io_reset; // @[:@55066.4 RegFile.scala 76:16:@55073.4]
  assign regs_381_io_in = 64'h0; // @[RegFile.scala 75:16:@55072.4]
  assign regs_381_io_reset = reset; // @[RegFile.scala 78:19:@55076.4]
  assign regs_381_io_enable = 1'h1; // @[RegFile.scala 74:20:@55070.4]
  assign regs_382_clock = clock; // @[:@55079.4]
  assign regs_382_reset = io_reset; // @[:@55080.4 RegFile.scala 76:16:@55087.4]
  assign regs_382_io_in = 64'h0; // @[RegFile.scala 75:16:@55086.4]
  assign regs_382_io_reset = reset; // @[RegFile.scala 78:19:@55090.4]
  assign regs_382_io_enable = 1'h1; // @[RegFile.scala 74:20:@55084.4]
  assign regs_383_clock = clock; // @[:@55093.4]
  assign regs_383_reset = io_reset; // @[:@55094.4 RegFile.scala 76:16:@55101.4]
  assign regs_383_io_in = 64'h0; // @[RegFile.scala 75:16:@55100.4]
  assign regs_383_io_reset = reset; // @[RegFile.scala 78:19:@55104.4]
  assign regs_383_io_enable = 1'h1; // @[RegFile.scala 74:20:@55098.4]
  assign regs_384_clock = clock; // @[:@55107.4]
  assign regs_384_reset = io_reset; // @[:@55108.4 RegFile.scala 76:16:@55115.4]
  assign regs_384_io_in = 64'h0; // @[RegFile.scala 75:16:@55114.4]
  assign regs_384_io_reset = reset; // @[RegFile.scala 78:19:@55118.4]
  assign regs_384_io_enable = 1'h1; // @[RegFile.scala 74:20:@55112.4]
  assign regs_385_clock = clock; // @[:@55121.4]
  assign regs_385_reset = io_reset; // @[:@55122.4 RegFile.scala 76:16:@55129.4]
  assign regs_385_io_in = 64'h0; // @[RegFile.scala 75:16:@55128.4]
  assign regs_385_io_reset = reset; // @[RegFile.scala 78:19:@55132.4]
  assign regs_385_io_enable = 1'h1; // @[RegFile.scala 74:20:@55126.4]
  assign regs_386_clock = clock; // @[:@55135.4]
  assign regs_386_reset = io_reset; // @[:@55136.4 RegFile.scala 76:16:@55143.4]
  assign regs_386_io_in = 64'h0; // @[RegFile.scala 75:16:@55142.4]
  assign regs_386_io_reset = reset; // @[RegFile.scala 78:19:@55146.4]
  assign regs_386_io_enable = 1'h1; // @[RegFile.scala 74:20:@55140.4]
  assign regs_387_clock = clock; // @[:@55149.4]
  assign regs_387_reset = io_reset; // @[:@55150.4 RegFile.scala 76:16:@55157.4]
  assign regs_387_io_in = 64'h0; // @[RegFile.scala 75:16:@55156.4]
  assign regs_387_io_reset = reset; // @[RegFile.scala 78:19:@55160.4]
  assign regs_387_io_enable = 1'h1; // @[RegFile.scala 74:20:@55154.4]
  assign regs_388_clock = clock; // @[:@55163.4]
  assign regs_388_reset = io_reset; // @[:@55164.4 RegFile.scala 76:16:@55171.4]
  assign regs_388_io_in = 64'h0; // @[RegFile.scala 75:16:@55170.4]
  assign regs_388_io_reset = reset; // @[RegFile.scala 78:19:@55174.4]
  assign regs_388_io_enable = 1'h1; // @[RegFile.scala 74:20:@55168.4]
  assign regs_389_clock = clock; // @[:@55177.4]
  assign regs_389_reset = io_reset; // @[:@55178.4 RegFile.scala 76:16:@55185.4]
  assign regs_389_io_in = 64'h0; // @[RegFile.scala 75:16:@55184.4]
  assign regs_389_io_reset = reset; // @[RegFile.scala 78:19:@55188.4]
  assign regs_389_io_enable = 1'h1; // @[RegFile.scala 74:20:@55182.4]
  assign regs_390_clock = clock; // @[:@55191.4]
  assign regs_390_reset = io_reset; // @[:@55192.4 RegFile.scala 76:16:@55199.4]
  assign regs_390_io_in = 64'h0; // @[RegFile.scala 75:16:@55198.4]
  assign regs_390_io_reset = reset; // @[RegFile.scala 78:19:@55202.4]
  assign regs_390_io_enable = 1'h1; // @[RegFile.scala 74:20:@55196.4]
  assign regs_391_clock = clock; // @[:@55205.4]
  assign regs_391_reset = io_reset; // @[:@55206.4 RegFile.scala 76:16:@55213.4]
  assign regs_391_io_in = 64'h0; // @[RegFile.scala 75:16:@55212.4]
  assign regs_391_io_reset = reset; // @[RegFile.scala 78:19:@55216.4]
  assign regs_391_io_enable = 1'h1; // @[RegFile.scala 74:20:@55210.4]
  assign regs_392_clock = clock; // @[:@55219.4]
  assign regs_392_reset = io_reset; // @[:@55220.4 RegFile.scala 76:16:@55227.4]
  assign regs_392_io_in = 64'h0; // @[RegFile.scala 75:16:@55226.4]
  assign regs_392_io_reset = reset; // @[RegFile.scala 78:19:@55230.4]
  assign regs_392_io_enable = 1'h1; // @[RegFile.scala 74:20:@55224.4]
  assign regs_393_clock = clock; // @[:@55233.4]
  assign regs_393_reset = io_reset; // @[:@55234.4 RegFile.scala 76:16:@55241.4]
  assign regs_393_io_in = 64'h0; // @[RegFile.scala 75:16:@55240.4]
  assign regs_393_io_reset = reset; // @[RegFile.scala 78:19:@55244.4]
  assign regs_393_io_enable = 1'h1; // @[RegFile.scala 74:20:@55238.4]
  assign regs_394_clock = clock; // @[:@55247.4]
  assign regs_394_reset = io_reset; // @[:@55248.4 RegFile.scala 76:16:@55255.4]
  assign regs_394_io_in = 64'h0; // @[RegFile.scala 75:16:@55254.4]
  assign regs_394_io_reset = reset; // @[RegFile.scala 78:19:@55258.4]
  assign regs_394_io_enable = 1'h1; // @[RegFile.scala 74:20:@55252.4]
  assign regs_395_clock = clock; // @[:@55261.4]
  assign regs_395_reset = io_reset; // @[:@55262.4 RegFile.scala 76:16:@55269.4]
  assign regs_395_io_in = 64'h0; // @[RegFile.scala 75:16:@55268.4]
  assign regs_395_io_reset = reset; // @[RegFile.scala 78:19:@55272.4]
  assign regs_395_io_enable = 1'h1; // @[RegFile.scala 74:20:@55266.4]
  assign regs_396_clock = clock; // @[:@55275.4]
  assign regs_396_reset = io_reset; // @[:@55276.4 RegFile.scala 76:16:@55283.4]
  assign regs_396_io_in = 64'h0; // @[RegFile.scala 75:16:@55282.4]
  assign regs_396_io_reset = reset; // @[RegFile.scala 78:19:@55286.4]
  assign regs_396_io_enable = 1'h1; // @[RegFile.scala 74:20:@55280.4]
  assign regs_397_clock = clock; // @[:@55289.4]
  assign regs_397_reset = io_reset; // @[:@55290.4 RegFile.scala 76:16:@55297.4]
  assign regs_397_io_in = 64'h0; // @[RegFile.scala 75:16:@55296.4]
  assign regs_397_io_reset = reset; // @[RegFile.scala 78:19:@55300.4]
  assign regs_397_io_enable = 1'h1; // @[RegFile.scala 74:20:@55294.4]
  assign regs_398_clock = clock; // @[:@55303.4]
  assign regs_398_reset = io_reset; // @[:@55304.4 RegFile.scala 76:16:@55311.4]
  assign regs_398_io_in = 64'h0; // @[RegFile.scala 75:16:@55310.4]
  assign regs_398_io_reset = reset; // @[RegFile.scala 78:19:@55314.4]
  assign regs_398_io_enable = 1'h1; // @[RegFile.scala 74:20:@55308.4]
  assign regs_399_clock = clock; // @[:@55317.4]
  assign regs_399_reset = io_reset; // @[:@55318.4 RegFile.scala 76:16:@55325.4]
  assign regs_399_io_in = 64'h0; // @[RegFile.scala 75:16:@55324.4]
  assign regs_399_io_reset = reset; // @[RegFile.scala 78:19:@55328.4]
  assign regs_399_io_enable = 1'h1; // @[RegFile.scala 74:20:@55322.4]
  assign regs_400_clock = clock; // @[:@55331.4]
  assign regs_400_reset = io_reset; // @[:@55332.4 RegFile.scala 76:16:@55339.4]
  assign regs_400_io_in = 64'h0; // @[RegFile.scala 75:16:@55338.4]
  assign regs_400_io_reset = reset; // @[RegFile.scala 78:19:@55342.4]
  assign regs_400_io_enable = 1'h1; // @[RegFile.scala 74:20:@55336.4]
  assign regs_401_clock = clock; // @[:@55345.4]
  assign regs_401_reset = io_reset; // @[:@55346.4 RegFile.scala 76:16:@55353.4]
  assign regs_401_io_in = 64'h0; // @[RegFile.scala 75:16:@55352.4]
  assign regs_401_io_reset = reset; // @[RegFile.scala 78:19:@55356.4]
  assign regs_401_io_enable = 1'h1; // @[RegFile.scala 74:20:@55350.4]
  assign regs_402_clock = clock; // @[:@55359.4]
  assign regs_402_reset = io_reset; // @[:@55360.4 RegFile.scala 76:16:@55367.4]
  assign regs_402_io_in = 64'h0; // @[RegFile.scala 75:16:@55366.4]
  assign regs_402_io_reset = reset; // @[RegFile.scala 78:19:@55370.4]
  assign regs_402_io_enable = 1'h1; // @[RegFile.scala 74:20:@55364.4]
  assign regs_403_clock = clock; // @[:@55373.4]
  assign regs_403_reset = io_reset; // @[:@55374.4 RegFile.scala 76:16:@55381.4]
  assign regs_403_io_in = 64'h0; // @[RegFile.scala 75:16:@55380.4]
  assign regs_403_io_reset = reset; // @[RegFile.scala 78:19:@55384.4]
  assign regs_403_io_enable = 1'h1; // @[RegFile.scala 74:20:@55378.4]
  assign regs_404_clock = clock; // @[:@55387.4]
  assign regs_404_reset = io_reset; // @[:@55388.4 RegFile.scala 76:16:@55395.4]
  assign regs_404_io_in = 64'h0; // @[RegFile.scala 75:16:@55394.4]
  assign regs_404_io_reset = reset; // @[RegFile.scala 78:19:@55398.4]
  assign regs_404_io_enable = 1'h1; // @[RegFile.scala 74:20:@55392.4]
  assign regs_405_clock = clock; // @[:@55401.4]
  assign regs_405_reset = io_reset; // @[:@55402.4 RegFile.scala 76:16:@55409.4]
  assign regs_405_io_in = 64'h0; // @[RegFile.scala 75:16:@55408.4]
  assign regs_405_io_reset = reset; // @[RegFile.scala 78:19:@55412.4]
  assign regs_405_io_enable = 1'h1; // @[RegFile.scala 74:20:@55406.4]
  assign regs_406_clock = clock; // @[:@55415.4]
  assign regs_406_reset = io_reset; // @[:@55416.4 RegFile.scala 76:16:@55423.4]
  assign regs_406_io_in = 64'h0; // @[RegFile.scala 75:16:@55422.4]
  assign regs_406_io_reset = reset; // @[RegFile.scala 78:19:@55426.4]
  assign regs_406_io_enable = 1'h1; // @[RegFile.scala 74:20:@55420.4]
  assign regs_407_clock = clock; // @[:@55429.4]
  assign regs_407_reset = io_reset; // @[:@55430.4 RegFile.scala 76:16:@55437.4]
  assign regs_407_io_in = 64'h0; // @[RegFile.scala 75:16:@55436.4]
  assign regs_407_io_reset = reset; // @[RegFile.scala 78:19:@55440.4]
  assign regs_407_io_enable = 1'h1; // @[RegFile.scala 74:20:@55434.4]
  assign regs_408_clock = clock; // @[:@55443.4]
  assign regs_408_reset = io_reset; // @[:@55444.4 RegFile.scala 76:16:@55451.4]
  assign regs_408_io_in = 64'h0; // @[RegFile.scala 75:16:@55450.4]
  assign regs_408_io_reset = reset; // @[RegFile.scala 78:19:@55454.4]
  assign regs_408_io_enable = 1'h1; // @[RegFile.scala 74:20:@55448.4]
  assign regs_409_clock = clock; // @[:@55457.4]
  assign regs_409_reset = io_reset; // @[:@55458.4 RegFile.scala 76:16:@55465.4]
  assign regs_409_io_in = 64'h0; // @[RegFile.scala 75:16:@55464.4]
  assign regs_409_io_reset = reset; // @[RegFile.scala 78:19:@55468.4]
  assign regs_409_io_enable = 1'h1; // @[RegFile.scala 74:20:@55462.4]
  assign regs_410_clock = clock; // @[:@55471.4]
  assign regs_410_reset = io_reset; // @[:@55472.4 RegFile.scala 76:16:@55479.4]
  assign regs_410_io_in = 64'h0; // @[RegFile.scala 75:16:@55478.4]
  assign regs_410_io_reset = reset; // @[RegFile.scala 78:19:@55482.4]
  assign regs_410_io_enable = 1'h1; // @[RegFile.scala 74:20:@55476.4]
  assign regs_411_clock = clock; // @[:@55485.4]
  assign regs_411_reset = io_reset; // @[:@55486.4 RegFile.scala 76:16:@55493.4]
  assign regs_411_io_in = 64'h0; // @[RegFile.scala 75:16:@55492.4]
  assign regs_411_io_reset = reset; // @[RegFile.scala 78:19:@55496.4]
  assign regs_411_io_enable = 1'h1; // @[RegFile.scala 74:20:@55490.4]
  assign regs_412_clock = clock; // @[:@55499.4]
  assign regs_412_reset = io_reset; // @[:@55500.4 RegFile.scala 76:16:@55507.4]
  assign regs_412_io_in = 64'h0; // @[RegFile.scala 75:16:@55506.4]
  assign regs_412_io_reset = reset; // @[RegFile.scala 78:19:@55510.4]
  assign regs_412_io_enable = 1'h1; // @[RegFile.scala 74:20:@55504.4]
  assign regs_413_clock = clock; // @[:@55513.4]
  assign regs_413_reset = io_reset; // @[:@55514.4 RegFile.scala 76:16:@55521.4]
  assign regs_413_io_in = 64'h0; // @[RegFile.scala 75:16:@55520.4]
  assign regs_413_io_reset = reset; // @[RegFile.scala 78:19:@55524.4]
  assign regs_413_io_enable = 1'h1; // @[RegFile.scala 74:20:@55518.4]
  assign regs_414_clock = clock; // @[:@55527.4]
  assign regs_414_reset = io_reset; // @[:@55528.4 RegFile.scala 76:16:@55535.4]
  assign regs_414_io_in = 64'h0; // @[RegFile.scala 75:16:@55534.4]
  assign regs_414_io_reset = reset; // @[RegFile.scala 78:19:@55538.4]
  assign regs_414_io_enable = 1'h1; // @[RegFile.scala 74:20:@55532.4]
  assign regs_415_clock = clock; // @[:@55541.4]
  assign regs_415_reset = io_reset; // @[:@55542.4 RegFile.scala 76:16:@55549.4]
  assign regs_415_io_in = 64'h0; // @[RegFile.scala 75:16:@55548.4]
  assign regs_415_io_reset = reset; // @[RegFile.scala 78:19:@55552.4]
  assign regs_415_io_enable = 1'h1; // @[RegFile.scala 74:20:@55546.4]
  assign regs_416_clock = clock; // @[:@55555.4]
  assign regs_416_reset = io_reset; // @[:@55556.4 RegFile.scala 76:16:@55563.4]
  assign regs_416_io_in = 64'h0; // @[RegFile.scala 75:16:@55562.4]
  assign regs_416_io_reset = reset; // @[RegFile.scala 78:19:@55566.4]
  assign regs_416_io_enable = 1'h1; // @[RegFile.scala 74:20:@55560.4]
  assign regs_417_clock = clock; // @[:@55569.4]
  assign regs_417_reset = io_reset; // @[:@55570.4 RegFile.scala 76:16:@55577.4]
  assign regs_417_io_in = 64'h0; // @[RegFile.scala 75:16:@55576.4]
  assign regs_417_io_reset = reset; // @[RegFile.scala 78:19:@55580.4]
  assign regs_417_io_enable = 1'h1; // @[RegFile.scala 74:20:@55574.4]
  assign regs_418_clock = clock; // @[:@55583.4]
  assign regs_418_reset = io_reset; // @[:@55584.4 RegFile.scala 76:16:@55591.4]
  assign regs_418_io_in = 64'h0; // @[RegFile.scala 75:16:@55590.4]
  assign regs_418_io_reset = reset; // @[RegFile.scala 78:19:@55594.4]
  assign regs_418_io_enable = 1'h1; // @[RegFile.scala 74:20:@55588.4]
  assign regs_419_clock = clock; // @[:@55597.4]
  assign regs_419_reset = io_reset; // @[:@55598.4 RegFile.scala 76:16:@55605.4]
  assign regs_419_io_in = 64'h0; // @[RegFile.scala 75:16:@55604.4]
  assign regs_419_io_reset = reset; // @[RegFile.scala 78:19:@55608.4]
  assign regs_419_io_enable = 1'h1; // @[RegFile.scala 74:20:@55602.4]
  assign regs_420_clock = clock; // @[:@55611.4]
  assign regs_420_reset = io_reset; // @[:@55612.4 RegFile.scala 76:16:@55619.4]
  assign regs_420_io_in = 64'h0; // @[RegFile.scala 75:16:@55618.4]
  assign regs_420_io_reset = reset; // @[RegFile.scala 78:19:@55622.4]
  assign regs_420_io_enable = 1'h1; // @[RegFile.scala 74:20:@55616.4]
  assign regs_421_clock = clock; // @[:@55625.4]
  assign regs_421_reset = io_reset; // @[:@55626.4 RegFile.scala 76:16:@55633.4]
  assign regs_421_io_in = 64'h0; // @[RegFile.scala 75:16:@55632.4]
  assign regs_421_io_reset = reset; // @[RegFile.scala 78:19:@55636.4]
  assign regs_421_io_enable = 1'h1; // @[RegFile.scala 74:20:@55630.4]
  assign regs_422_clock = clock; // @[:@55639.4]
  assign regs_422_reset = io_reset; // @[:@55640.4 RegFile.scala 76:16:@55647.4]
  assign regs_422_io_in = 64'h0; // @[RegFile.scala 75:16:@55646.4]
  assign regs_422_io_reset = reset; // @[RegFile.scala 78:19:@55650.4]
  assign regs_422_io_enable = 1'h1; // @[RegFile.scala 74:20:@55644.4]
  assign regs_423_clock = clock; // @[:@55653.4]
  assign regs_423_reset = io_reset; // @[:@55654.4 RegFile.scala 76:16:@55661.4]
  assign regs_423_io_in = 64'h0; // @[RegFile.scala 75:16:@55660.4]
  assign regs_423_io_reset = reset; // @[RegFile.scala 78:19:@55664.4]
  assign regs_423_io_enable = 1'h1; // @[RegFile.scala 74:20:@55658.4]
  assign regs_424_clock = clock; // @[:@55667.4]
  assign regs_424_reset = io_reset; // @[:@55668.4 RegFile.scala 76:16:@55675.4]
  assign regs_424_io_in = 64'h0; // @[RegFile.scala 75:16:@55674.4]
  assign regs_424_io_reset = reset; // @[RegFile.scala 78:19:@55678.4]
  assign regs_424_io_enable = 1'h1; // @[RegFile.scala 74:20:@55672.4]
  assign regs_425_clock = clock; // @[:@55681.4]
  assign regs_425_reset = io_reset; // @[:@55682.4 RegFile.scala 76:16:@55689.4]
  assign regs_425_io_in = 64'h0; // @[RegFile.scala 75:16:@55688.4]
  assign regs_425_io_reset = reset; // @[RegFile.scala 78:19:@55692.4]
  assign regs_425_io_enable = 1'h1; // @[RegFile.scala 74:20:@55686.4]
  assign regs_426_clock = clock; // @[:@55695.4]
  assign regs_426_reset = io_reset; // @[:@55696.4 RegFile.scala 76:16:@55703.4]
  assign regs_426_io_in = 64'h0; // @[RegFile.scala 75:16:@55702.4]
  assign regs_426_io_reset = reset; // @[RegFile.scala 78:19:@55706.4]
  assign regs_426_io_enable = 1'h1; // @[RegFile.scala 74:20:@55700.4]
  assign regs_427_clock = clock; // @[:@55709.4]
  assign regs_427_reset = io_reset; // @[:@55710.4 RegFile.scala 76:16:@55717.4]
  assign regs_427_io_in = 64'h0; // @[RegFile.scala 75:16:@55716.4]
  assign regs_427_io_reset = reset; // @[RegFile.scala 78:19:@55720.4]
  assign regs_427_io_enable = 1'h1; // @[RegFile.scala 74:20:@55714.4]
  assign regs_428_clock = clock; // @[:@55723.4]
  assign regs_428_reset = io_reset; // @[:@55724.4 RegFile.scala 76:16:@55731.4]
  assign regs_428_io_in = 64'h0; // @[RegFile.scala 75:16:@55730.4]
  assign regs_428_io_reset = reset; // @[RegFile.scala 78:19:@55734.4]
  assign regs_428_io_enable = 1'h1; // @[RegFile.scala 74:20:@55728.4]
  assign regs_429_clock = clock; // @[:@55737.4]
  assign regs_429_reset = io_reset; // @[:@55738.4 RegFile.scala 76:16:@55745.4]
  assign regs_429_io_in = 64'h0; // @[RegFile.scala 75:16:@55744.4]
  assign regs_429_io_reset = reset; // @[RegFile.scala 78:19:@55748.4]
  assign regs_429_io_enable = 1'h1; // @[RegFile.scala 74:20:@55742.4]
  assign regs_430_clock = clock; // @[:@55751.4]
  assign regs_430_reset = io_reset; // @[:@55752.4 RegFile.scala 76:16:@55759.4]
  assign regs_430_io_in = 64'h0; // @[RegFile.scala 75:16:@55758.4]
  assign regs_430_io_reset = reset; // @[RegFile.scala 78:19:@55762.4]
  assign regs_430_io_enable = 1'h1; // @[RegFile.scala 74:20:@55756.4]
  assign regs_431_clock = clock; // @[:@55765.4]
  assign regs_431_reset = io_reset; // @[:@55766.4 RegFile.scala 76:16:@55773.4]
  assign regs_431_io_in = 64'h0; // @[RegFile.scala 75:16:@55772.4]
  assign regs_431_io_reset = reset; // @[RegFile.scala 78:19:@55776.4]
  assign regs_431_io_enable = 1'h1; // @[RegFile.scala 74:20:@55770.4]
  assign regs_432_clock = clock; // @[:@55779.4]
  assign regs_432_reset = io_reset; // @[:@55780.4 RegFile.scala 76:16:@55787.4]
  assign regs_432_io_in = 64'h0; // @[RegFile.scala 75:16:@55786.4]
  assign regs_432_io_reset = reset; // @[RegFile.scala 78:19:@55790.4]
  assign regs_432_io_enable = 1'h1; // @[RegFile.scala 74:20:@55784.4]
  assign regs_433_clock = clock; // @[:@55793.4]
  assign regs_433_reset = io_reset; // @[:@55794.4 RegFile.scala 76:16:@55801.4]
  assign regs_433_io_in = 64'h0; // @[RegFile.scala 75:16:@55800.4]
  assign regs_433_io_reset = reset; // @[RegFile.scala 78:19:@55804.4]
  assign regs_433_io_enable = 1'h1; // @[RegFile.scala 74:20:@55798.4]
  assign regs_434_clock = clock; // @[:@55807.4]
  assign regs_434_reset = io_reset; // @[:@55808.4 RegFile.scala 76:16:@55815.4]
  assign regs_434_io_in = 64'h0; // @[RegFile.scala 75:16:@55814.4]
  assign regs_434_io_reset = reset; // @[RegFile.scala 78:19:@55818.4]
  assign regs_434_io_enable = 1'h1; // @[RegFile.scala 74:20:@55812.4]
  assign regs_435_clock = clock; // @[:@55821.4]
  assign regs_435_reset = io_reset; // @[:@55822.4 RegFile.scala 76:16:@55829.4]
  assign regs_435_io_in = 64'h0; // @[RegFile.scala 75:16:@55828.4]
  assign regs_435_io_reset = reset; // @[RegFile.scala 78:19:@55832.4]
  assign regs_435_io_enable = 1'h1; // @[RegFile.scala 74:20:@55826.4]
  assign regs_436_clock = clock; // @[:@55835.4]
  assign regs_436_reset = io_reset; // @[:@55836.4 RegFile.scala 76:16:@55843.4]
  assign regs_436_io_in = 64'h0; // @[RegFile.scala 75:16:@55842.4]
  assign regs_436_io_reset = reset; // @[RegFile.scala 78:19:@55846.4]
  assign regs_436_io_enable = 1'h1; // @[RegFile.scala 74:20:@55840.4]
  assign regs_437_clock = clock; // @[:@55849.4]
  assign regs_437_reset = io_reset; // @[:@55850.4 RegFile.scala 76:16:@55857.4]
  assign regs_437_io_in = 64'h0; // @[RegFile.scala 75:16:@55856.4]
  assign regs_437_io_reset = reset; // @[RegFile.scala 78:19:@55860.4]
  assign regs_437_io_enable = 1'h1; // @[RegFile.scala 74:20:@55854.4]
  assign regs_438_clock = clock; // @[:@55863.4]
  assign regs_438_reset = io_reset; // @[:@55864.4 RegFile.scala 76:16:@55871.4]
  assign regs_438_io_in = 64'h0; // @[RegFile.scala 75:16:@55870.4]
  assign regs_438_io_reset = reset; // @[RegFile.scala 78:19:@55874.4]
  assign regs_438_io_enable = 1'h1; // @[RegFile.scala 74:20:@55868.4]
  assign regs_439_clock = clock; // @[:@55877.4]
  assign regs_439_reset = io_reset; // @[:@55878.4 RegFile.scala 76:16:@55885.4]
  assign regs_439_io_in = 64'h0; // @[RegFile.scala 75:16:@55884.4]
  assign regs_439_io_reset = reset; // @[RegFile.scala 78:19:@55888.4]
  assign regs_439_io_enable = 1'h1; // @[RegFile.scala 74:20:@55882.4]
  assign regs_440_clock = clock; // @[:@55891.4]
  assign regs_440_reset = io_reset; // @[:@55892.4 RegFile.scala 76:16:@55899.4]
  assign regs_440_io_in = 64'h0; // @[RegFile.scala 75:16:@55898.4]
  assign regs_440_io_reset = reset; // @[RegFile.scala 78:19:@55902.4]
  assign regs_440_io_enable = 1'h1; // @[RegFile.scala 74:20:@55896.4]
  assign regs_441_clock = clock; // @[:@55905.4]
  assign regs_441_reset = io_reset; // @[:@55906.4 RegFile.scala 76:16:@55913.4]
  assign regs_441_io_in = 64'h0; // @[RegFile.scala 75:16:@55912.4]
  assign regs_441_io_reset = reset; // @[RegFile.scala 78:19:@55916.4]
  assign regs_441_io_enable = 1'h1; // @[RegFile.scala 74:20:@55910.4]
  assign regs_442_clock = clock; // @[:@55919.4]
  assign regs_442_reset = io_reset; // @[:@55920.4 RegFile.scala 76:16:@55927.4]
  assign regs_442_io_in = 64'h0; // @[RegFile.scala 75:16:@55926.4]
  assign regs_442_io_reset = reset; // @[RegFile.scala 78:19:@55930.4]
  assign regs_442_io_enable = 1'h1; // @[RegFile.scala 74:20:@55924.4]
  assign regs_443_clock = clock; // @[:@55933.4]
  assign regs_443_reset = io_reset; // @[:@55934.4 RegFile.scala 76:16:@55941.4]
  assign regs_443_io_in = 64'h0; // @[RegFile.scala 75:16:@55940.4]
  assign regs_443_io_reset = reset; // @[RegFile.scala 78:19:@55944.4]
  assign regs_443_io_enable = 1'h1; // @[RegFile.scala 74:20:@55938.4]
  assign regs_444_clock = clock; // @[:@55947.4]
  assign regs_444_reset = io_reset; // @[:@55948.4 RegFile.scala 76:16:@55955.4]
  assign regs_444_io_in = 64'h0; // @[RegFile.scala 75:16:@55954.4]
  assign regs_444_io_reset = reset; // @[RegFile.scala 78:19:@55958.4]
  assign regs_444_io_enable = 1'h1; // @[RegFile.scala 74:20:@55952.4]
  assign regs_445_clock = clock; // @[:@55961.4]
  assign regs_445_reset = io_reset; // @[:@55962.4 RegFile.scala 76:16:@55969.4]
  assign regs_445_io_in = 64'h0; // @[RegFile.scala 75:16:@55968.4]
  assign regs_445_io_reset = reset; // @[RegFile.scala 78:19:@55972.4]
  assign regs_445_io_enable = 1'h1; // @[RegFile.scala 74:20:@55966.4]
  assign regs_446_clock = clock; // @[:@55975.4]
  assign regs_446_reset = io_reset; // @[:@55976.4 RegFile.scala 76:16:@55983.4]
  assign regs_446_io_in = 64'h0; // @[RegFile.scala 75:16:@55982.4]
  assign regs_446_io_reset = reset; // @[RegFile.scala 78:19:@55986.4]
  assign regs_446_io_enable = 1'h1; // @[RegFile.scala 74:20:@55980.4]
  assign regs_447_clock = clock; // @[:@55989.4]
  assign regs_447_reset = io_reset; // @[:@55990.4 RegFile.scala 76:16:@55997.4]
  assign regs_447_io_in = 64'h0; // @[RegFile.scala 75:16:@55996.4]
  assign regs_447_io_reset = reset; // @[RegFile.scala 78:19:@56000.4]
  assign regs_447_io_enable = 1'h1; // @[RegFile.scala 74:20:@55994.4]
  assign regs_448_clock = clock; // @[:@56003.4]
  assign regs_448_reset = io_reset; // @[:@56004.4 RegFile.scala 76:16:@56011.4]
  assign regs_448_io_in = 64'h0; // @[RegFile.scala 75:16:@56010.4]
  assign regs_448_io_reset = reset; // @[RegFile.scala 78:19:@56014.4]
  assign regs_448_io_enable = 1'h1; // @[RegFile.scala 74:20:@56008.4]
  assign regs_449_clock = clock; // @[:@56017.4]
  assign regs_449_reset = io_reset; // @[:@56018.4 RegFile.scala 76:16:@56025.4]
  assign regs_449_io_in = 64'h0; // @[RegFile.scala 75:16:@56024.4]
  assign regs_449_io_reset = reset; // @[RegFile.scala 78:19:@56028.4]
  assign regs_449_io_enable = 1'h1; // @[RegFile.scala 74:20:@56022.4]
  assign regs_450_clock = clock; // @[:@56031.4]
  assign regs_450_reset = io_reset; // @[:@56032.4 RegFile.scala 76:16:@56039.4]
  assign regs_450_io_in = 64'h0; // @[RegFile.scala 75:16:@56038.4]
  assign regs_450_io_reset = reset; // @[RegFile.scala 78:19:@56042.4]
  assign regs_450_io_enable = 1'h1; // @[RegFile.scala 74:20:@56036.4]
  assign regs_451_clock = clock; // @[:@56045.4]
  assign regs_451_reset = io_reset; // @[:@56046.4 RegFile.scala 76:16:@56053.4]
  assign regs_451_io_in = 64'h0; // @[RegFile.scala 75:16:@56052.4]
  assign regs_451_io_reset = reset; // @[RegFile.scala 78:19:@56056.4]
  assign regs_451_io_enable = 1'h1; // @[RegFile.scala 74:20:@56050.4]
  assign regs_452_clock = clock; // @[:@56059.4]
  assign regs_452_reset = io_reset; // @[:@56060.4 RegFile.scala 76:16:@56067.4]
  assign regs_452_io_in = 64'h0; // @[RegFile.scala 75:16:@56066.4]
  assign regs_452_io_reset = reset; // @[RegFile.scala 78:19:@56070.4]
  assign regs_452_io_enable = 1'h1; // @[RegFile.scala 74:20:@56064.4]
  assign regs_453_clock = clock; // @[:@56073.4]
  assign regs_453_reset = io_reset; // @[:@56074.4 RegFile.scala 76:16:@56081.4]
  assign regs_453_io_in = 64'h0; // @[RegFile.scala 75:16:@56080.4]
  assign regs_453_io_reset = reset; // @[RegFile.scala 78:19:@56084.4]
  assign regs_453_io_enable = 1'h1; // @[RegFile.scala 74:20:@56078.4]
  assign regs_454_clock = clock; // @[:@56087.4]
  assign regs_454_reset = io_reset; // @[:@56088.4 RegFile.scala 76:16:@56095.4]
  assign regs_454_io_in = 64'h0; // @[RegFile.scala 75:16:@56094.4]
  assign regs_454_io_reset = reset; // @[RegFile.scala 78:19:@56098.4]
  assign regs_454_io_enable = 1'h1; // @[RegFile.scala 74:20:@56092.4]
  assign regs_455_clock = clock; // @[:@56101.4]
  assign regs_455_reset = io_reset; // @[:@56102.4 RegFile.scala 76:16:@56109.4]
  assign regs_455_io_in = 64'h0; // @[RegFile.scala 75:16:@56108.4]
  assign regs_455_io_reset = reset; // @[RegFile.scala 78:19:@56112.4]
  assign regs_455_io_enable = 1'h1; // @[RegFile.scala 74:20:@56106.4]
  assign regs_456_clock = clock; // @[:@56115.4]
  assign regs_456_reset = io_reset; // @[:@56116.4 RegFile.scala 76:16:@56123.4]
  assign regs_456_io_in = 64'h0; // @[RegFile.scala 75:16:@56122.4]
  assign regs_456_io_reset = reset; // @[RegFile.scala 78:19:@56126.4]
  assign regs_456_io_enable = 1'h1; // @[RegFile.scala 74:20:@56120.4]
  assign regs_457_clock = clock; // @[:@56129.4]
  assign regs_457_reset = io_reset; // @[:@56130.4 RegFile.scala 76:16:@56137.4]
  assign regs_457_io_in = 64'h0; // @[RegFile.scala 75:16:@56136.4]
  assign regs_457_io_reset = reset; // @[RegFile.scala 78:19:@56140.4]
  assign regs_457_io_enable = 1'h1; // @[RegFile.scala 74:20:@56134.4]
  assign regs_458_clock = clock; // @[:@56143.4]
  assign regs_458_reset = io_reset; // @[:@56144.4 RegFile.scala 76:16:@56151.4]
  assign regs_458_io_in = 64'h0; // @[RegFile.scala 75:16:@56150.4]
  assign regs_458_io_reset = reset; // @[RegFile.scala 78:19:@56154.4]
  assign regs_458_io_enable = 1'h1; // @[RegFile.scala 74:20:@56148.4]
  assign regs_459_clock = clock; // @[:@56157.4]
  assign regs_459_reset = io_reset; // @[:@56158.4 RegFile.scala 76:16:@56165.4]
  assign regs_459_io_in = 64'h0; // @[RegFile.scala 75:16:@56164.4]
  assign regs_459_io_reset = reset; // @[RegFile.scala 78:19:@56168.4]
  assign regs_459_io_enable = 1'h1; // @[RegFile.scala 74:20:@56162.4]
  assign regs_460_clock = clock; // @[:@56171.4]
  assign regs_460_reset = io_reset; // @[:@56172.4 RegFile.scala 76:16:@56179.4]
  assign regs_460_io_in = 64'h0; // @[RegFile.scala 75:16:@56178.4]
  assign regs_460_io_reset = reset; // @[RegFile.scala 78:19:@56182.4]
  assign regs_460_io_enable = 1'h1; // @[RegFile.scala 74:20:@56176.4]
  assign regs_461_clock = clock; // @[:@56185.4]
  assign regs_461_reset = io_reset; // @[:@56186.4 RegFile.scala 76:16:@56193.4]
  assign regs_461_io_in = 64'h0; // @[RegFile.scala 75:16:@56192.4]
  assign regs_461_io_reset = reset; // @[RegFile.scala 78:19:@56196.4]
  assign regs_461_io_enable = 1'h1; // @[RegFile.scala 74:20:@56190.4]
  assign regs_462_clock = clock; // @[:@56199.4]
  assign regs_462_reset = io_reset; // @[:@56200.4 RegFile.scala 76:16:@56207.4]
  assign regs_462_io_in = 64'h0; // @[RegFile.scala 75:16:@56206.4]
  assign regs_462_io_reset = reset; // @[RegFile.scala 78:19:@56210.4]
  assign regs_462_io_enable = 1'h1; // @[RegFile.scala 74:20:@56204.4]
  assign regs_463_clock = clock; // @[:@56213.4]
  assign regs_463_reset = io_reset; // @[:@56214.4 RegFile.scala 76:16:@56221.4]
  assign regs_463_io_in = 64'h0; // @[RegFile.scala 75:16:@56220.4]
  assign regs_463_io_reset = reset; // @[RegFile.scala 78:19:@56224.4]
  assign regs_463_io_enable = 1'h1; // @[RegFile.scala 74:20:@56218.4]
  assign regs_464_clock = clock; // @[:@56227.4]
  assign regs_464_reset = io_reset; // @[:@56228.4 RegFile.scala 76:16:@56235.4]
  assign regs_464_io_in = 64'h0; // @[RegFile.scala 75:16:@56234.4]
  assign regs_464_io_reset = reset; // @[RegFile.scala 78:19:@56238.4]
  assign regs_464_io_enable = 1'h1; // @[RegFile.scala 74:20:@56232.4]
  assign regs_465_clock = clock; // @[:@56241.4]
  assign regs_465_reset = io_reset; // @[:@56242.4 RegFile.scala 76:16:@56249.4]
  assign regs_465_io_in = 64'h0; // @[RegFile.scala 75:16:@56248.4]
  assign regs_465_io_reset = reset; // @[RegFile.scala 78:19:@56252.4]
  assign regs_465_io_enable = 1'h1; // @[RegFile.scala 74:20:@56246.4]
  assign regs_466_clock = clock; // @[:@56255.4]
  assign regs_466_reset = io_reset; // @[:@56256.4 RegFile.scala 76:16:@56263.4]
  assign regs_466_io_in = 64'h0; // @[RegFile.scala 75:16:@56262.4]
  assign regs_466_io_reset = reset; // @[RegFile.scala 78:19:@56266.4]
  assign regs_466_io_enable = 1'h1; // @[RegFile.scala 74:20:@56260.4]
  assign regs_467_clock = clock; // @[:@56269.4]
  assign regs_467_reset = io_reset; // @[:@56270.4 RegFile.scala 76:16:@56277.4]
  assign regs_467_io_in = 64'h0; // @[RegFile.scala 75:16:@56276.4]
  assign regs_467_io_reset = reset; // @[RegFile.scala 78:19:@56280.4]
  assign regs_467_io_enable = 1'h1; // @[RegFile.scala 74:20:@56274.4]
  assign regs_468_clock = clock; // @[:@56283.4]
  assign regs_468_reset = io_reset; // @[:@56284.4 RegFile.scala 76:16:@56291.4]
  assign regs_468_io_in = 64'h0; // @[RegFile.scala 75:16:@56290.4]
  assign regs_468_io_reset = reset; // @[RegFile.scala 78:19:@56294.4]
  assign regs_468_io_enable = 1'h1; // @[RegFile.scala 74:20:@56288.4]
  assign regs_469_clock = clock; // @[:@56297.4]
  assign regs_469_reset = io_reset; // @[:@56298.4 RegFile.scala 76:16:@56305.4]
  assign regs_469_io_in = 64'h0; // @[RegFile.scala 75:16:@56304.4]
  assign regs_469_io_reset = reset; // @[RegFile.scala 78:19:@56308.4]
  assign regs_469_io_enable = 1'h1; // @[RegFile.scala 74:20:@56302.4]
  assign regs_470_clock = clock; // @[:@56311.4]
  assign regs_470_reset = io_reset; // @[:@56312.4 RegFile.scala 76:16:@56319.4]
  assign regs_470_io_in = 64'h0; // @[RegFile.scala 75:16:@56318.4]
  assign regs_470_io_reset = reset; // @[RegFile.scala 78:19:@56322.4]
  assign regs_470_io_enable = 1'h1; // @[RegFile.scala 74:20:@56316.4]
  assign regs_471_clock = clock; // @[:@56325.4]
  assign regs_471_reset = io_reset; // @[:@56326.4 RegFile.scala 76:16:@56333.4]
  assign regs_471_io_in = 64'h0; // @[RegFile.scala 75:16:@56332.4]
  assign regs_471_io_reset = reset; // @[RegFile.scala 78:19:@56336.4]
  assign regs_471_io_enable = 1'h1; // @[RegFile.scala 74:20:@56330.4]
  assign regs_472_clock = clock; // @[:@56339.4]
  assign regs_472_reset = io_reset; // @[:@56340.4 RegFile.scala 76:16:@56347.4]
  assign regs_472_io_in = 64'h0; // @[RegFile.scala 75:16:@56346.4]
  assign regs_472_io_reset = reset; // @[RegFile.scala 78:19:@56350.4]
  assign regs_472_io_enable = 1'h1; // @[RegFile.scala 74:20:@56344.4]
  assign regs_473_clock = clock; // @[:@56353.4]
  assign regs_473_reset = io_reset; // @[:@56354.4 RegFile.scala 76:16:@56361.4]
  assign regs_473_io_in = 64'h0; // @[RegFile.scala 75:16:@56360.4]
  assign regs_473_io_reset = reset; // @[RegFile.scala 78:19:@56364.4]
  assign regs_473_io_enable = 1'h1; // @[RegFile.scala 74:20:@56358.4]
  assign regs_474_clock = clock; // @[:@56367.4]
  assign regs_474_reset = io_reset; // @[:@56368.4 RegFile.scala 76:16:@56375.4]
  assign regs_474_io_in = 64'h0; // @[RegFile.scala 75:16:@56374.4]
  assign regs_474_io_reset = reset; // @[RegFile.scala 78:19:@56378.4]
  assign regs_474_io_enable = 1'h1; // @[RegFile.scala 74:20:@56372.4]
  assign regs_475_clock = clock; // @[:@56381.4]
  assign regs_475_reset = io_reset; // @[:@56382.4 RegFile.scala 76:16:@56389.4]
  assign regs_475_io_in = 64'h0; // @[RegFile.scala 75:16:@56388.4]
  assign regs_475_io_reset = reset; // @[RegFile.scala 78:19:@56392.4]
  assign regs_475_io_enable = 1'h1; // @[RegFile.scala 74:20:@56386.4]
  assign regs_476_clock = clock; // @[:@56395.4]
  assign regs_476_reset = io_reset; // @[:@56396.4 RegFile.scala 76:16:@56403.4]
  assign regs_476_io_in = 64'h0; // @[RegFile.scala 75:16:@56402.4]
  assign regs_476_io_reset = reset; // @[RegFile.scala 78:19:@56406.4]
  assign regs_476_io_enable = 1'h1; // @[RegFile.scala 74:20:@56400.4]
  assign regs_477_clock = clock; // @[:@56409.4]
  assign regs_477_reset = io_reset; // @[:@56410.4 RegFile.scala 76:16:@56417.4]
  assign regs_477_io_in = 64'h0; // @[RegFile.scala 75:16:@56416.4]
  assign regs_477_io_reset = reset; // @[RegFile.scala 78:19:@56420.4]
  assign regs_477_io_enable = 1'h1; // @[RegFile.scala 74:20:@56414.4]
  assign regs_478_clock = clock; // @[:@56423.4]
  assign regs_478_reset = io_reset; // @[:@56424.4 RegFile.scala 76:16:@56431.4]
  assign regs_478_io_in = 64'h0; // @[RegFile.scala 75:16:@56430.4]
  assign regs_478_io_reset = reset; // @[RegFile.scala 78:19:@56434.4]
  assign regs_478_io_enable = 1'h1; // @[RegFile.scala 74:20:@56428.4]
  assign regs_479_clock = clock; // @[:@56437.4]
  assign regs_479_reset = io_reset; // @[:@56438.4 RegFile.scala 76:16:@56445.4]
  assign regs_479_io_in = 64'h0; // @[RegFile.scala 75:16:@56444.4]
  assign regs_479_io_reset = reset; // @[RegFile.scala 78:19:@56448.4]
  assign regs_479_io_enable = 1'h1; // @[RegFile.scala 74:20:@56442.4]
  assign regs_480_clock = clock; // @[:@56451.4]
  assign regs_480_reset = io_reset; // @[:@56452.4 RegFile.scala 76:16:@56459.4]
  assign regs_480_io_in = 64'h0; // @[RegFile.scala 75:16:@56458.4]
  assign regs_480_io_reset = reset; // @[RegFile.scala 78:19:@56462.4]
  assign regs_480_io_enable = 1'h1; // @[RegFile.scala 74:20:@56456.4]
  assign regs_481_clock = clock; // @[:@56465.4]
  assign regs_481_reset = io_reset; // @[:@56466.4 RegFile.scala 76:16:@56473.4]
  assign regs_481_io_in = 64'h0; // @[RegFile.scala 75:16:@56472.4]
  assign regs_481_io_reset = reset; // @[RegFile.scala 78:19:@56476.4]
  assign regs_481_io_enable = 1'h1; // @[RegFile.scala 74:20:@56470.4]
  assign regs_482_clock = clock; // @[:@56479.4]
  assign regs_482_reset = io_reset; // @[:@56480.4 RegFile.scala 76:16:@56487.4]
  assign regs_482_io_in = 64'h0; // @[RegFile.scala 75:16:@56486.4]
  assign regs_482_io_reset = reset; // @[RegFile.scala 78:19:@56490.4]
  assign regs_482_io_enable = 1'h1; // @[RegFile.scala 74:20:@56484.4]
  assign regs_483_clock = clock; // @[:@56493.4]
  assign regs_483_reset = io_reset; // @[:@56494.4 RegFile.scala 76:16:@56501.4]
  assign regs_483_io_in = 64'h0; // @[RegFile.scala 75:16:@56500.4]
  assign regs_483_io_reset = reset; // @[RegFile.scala 78:19:@56504.4]
  assign regs_483_io_enable = 1'h1; // @[RegFile.scala 74:20:@56498.4]
  assign regs_484_clock = clock; // @[:@56507.4]
  assign regs_484_reset = io_reset; // @[:@56508.4 RegFile.scala 76:16:@56515.4]
  assign regs_484_io_in = 64'h0; // @[RegFile.scala 75:16:@56514.4]
  assign regs_484_io_reset = reset; // @[RegFile.scala 78:19:@56518.4]
  assign regs_484_io_enable = 1'h1; // @[RegFile.scala 74:20:@56512.4]
  assign regs_485_clock = clock; // @[:@56521.4]
  assign regs_485_reset = io_reset; // @[:@56522.4 RegFile.scala 76:16:@56529.4]
  assign regs_485_io_in = 64'h0; // @[RegFile.scala 75:16:@56528.4]
  assign regs_485_io_reset = reset; // @[RegFile.scala 78:19:@56532.4]
  assign regs_485_io_enable = 1'h1; // @[RegFile.scala 74:20:@56526.4]
  assign regs_486_clock = clock; // @[:@56535.4]
  assign regs_486_reset = io_reset; // @[:@56536.4 RegFile.scala 76:16:@56543.4]
  assign regs_486_io_in = 64'h0; // @[RegFile.scala 75:16:@56542.4]
  assign regs_486_io_reset = reset; // @[RegFile.scala 78:19:@56546.4]
  assign regs_486_io_enable = 1'h1; // @[RegFile.scala 74:20:@56540.4]
  assign regs_487_clock = clock; // @[:@56549.4]
  assign regs_487_reset = io_reset; // @[:@56550.4 RegFile.scala 76:16:@56557.4]
  assign regs_487_io_in = 64'h0; // @[RegFile.scala 75:16:@56556.4]
  assign regs_487_io_reset = reset; // @[RegFile.scala 78:19:@56560.4]
  assign regs_487_io_enable = 1'h1; // @[RegFile.scala 74:20:@56554.4]
  assign regs_488_clock = clock; // @[:@56563.4]
  assign regs_488_reset = io_reset; // @[:@56564.4 RegFile.scala 76:16:@56571.4]
  assign regs_488_io_in = 64'h0; // @[RegFile.scala 75:16:@56570.4]
  assign regs_488_io_reset = reset; // @[RegFile.scala 78:19:@56574.4]
  assign regs_488_io_enable = 1'h1; // @[RegFile.scala 74:20:@56568.4]
  assign regs_489_clock = clock; // @[:@56577.4]
  assign regs_489_reset = io_reset; // @[:@56578.4 RegFile.scala 76:16:@56585.4]
  assign regs_489_io_in = 64'h0; // @[RegFile.scala 75:16:@56584.4]
  assign regs_489_io_reset = reset; // @[RegFile.scala 78:19:@56588.4]
  assign regs_489_io_enable = 1'h1; // @[RegFile.scala 74:20:@56582.4]
  assign regs_490_clock = clock; // @[:@56591.4]
  assign regs_490_reset = io_reset; // @[:@56592.4 RegFile.scala 76:16:@56599.4]
  assign regs_490_io_in = 64'h0; // @[RegFile.scala 75:16:@56598.4]
  assign regs_490_io_reset = reset; // @[RegFile.scala 78:19:@56602.4]
  assign regs_490_io_enable = 1'h1; // @[RegFile.scala 74:20:@56596.4]
  assign regs_491_clock = clock; // @[:@56605.4]
  assign regs_491_reset = io_reset; // @[:@56606.4 RegFile.scala 76:16:@56613.4]
  assign regs_491_io_in = 64'h0; // @[RegFile.scala 75:16:@56612.4]
  assign regs_491_io_reset = reset; // @[RegFile.scala 78:19:@56616.4]
  assign regs_491_io_enable = 1'h1; // @[RegFile.scala 74:20:@56610.4]
  assign regs_492_clock = clock; // @[:@56619.4]
  assign regs_492_reset = io_reset; // @[:@56620.4 RegFile.scala 76:16:@56627.4]
  assign regs_492_io_in = 64'h0; // @[RegFile.scala 75:16:@56626.4]
  assign regs_492_io_reset = reset; // @[RegFile.scala 78:19:@56630.4]
  assign regs_492_io_enable = 1'h1; // @[RegFile.scala 74:20:@56624.4]
  assign regs_493_clock = clock; // @[:@56633.4]
  assign regs_493_reset = io_reset; // @[:@56634.4 RegFile.scala 76:16:@56641.4]
  assign regs_493_io_in = 64'h0; // @[RegFile.scala 75:16:@56640.4]
  assign regs_493_io_reset = reset; // @[RegFile.scala 78:19:@56644.4]
  assign regs_493_io_enable = 1'h1; // @[RegFile.scala 74:20:@56638.4]
  assign regs_494_clock = clock; // @[:@56647.4]
  assign regs_494_reset = io_reset; // @[:@56648.4 RegFile.scala 76:16:@56655.4]
  assign regs_494_io_in = 64'h0; // @[RegFile.scala 75:16:@56654.4]
  assign regs_494_io_reset = reset; // @[RegFile.scala 78:19:@56658.4]
  assign regs_494_io_enable = 1'h1; // @[RegFile.scala 74:20:@56652.4]
  assign regs_495_clock = clock; // @[:@56661.4]
  assign regs_495_reset = io_reset; // @[:@56662.4 RegFile.scala 76:16:@56669.4]
  assign regs_495_io_in = 64'h0; // @[RegFile.scala 75:16:@56668.4]
  assign regs_495_io_reset = reset; // @[RegFile.scala 78:19:@56672.4]
  assign regs_495_io_enable = 1'h1; // @[RegFile.scala 74:20:@56666.4]
  assign regs_496_clock = clock; // @[:@56675.4]
  assign regs_496_reset = io_reset; // @[:@56676.4 RegFile.scala 76:16:@56683.4]
  assign regs_496_io_in = 64'h0; // @[RegFile.scala 75:16:@56682.4]
  assign regs_496_io_reset = reset; // @[RegFile.scala 78:19:@56686.4]
  assign regs_496_io_enable = 1'h1; // @[RegFile.scala 74:20:@56680.4]
  assign regs_497_clock = clock; // @[:@56689.4]
  assign regs_497_reset = io_reset; // @[:@56690.4 RegFile.scala 76:16:@56697.4]
  assign regs_497_io_in = 64'h0; // @[RegFile.scala 75:16:@56696.4]
  assign regs_497_io_reset = reset; // @[RegFile.scala 78:19:@56700.4]
  assign regs_497_io_enable = 1'h1; // @[RegFile.scala 74:20:@56694.4]
  assign regs_498_clock = clock; // @[:@56703.4]
  assign regs_498_reset = io_reset; // @[:@56704.4 RegFile.scala 76:16:@56711.4]
  assign regs_498_io_in = 64'h0; // @[RegFile.scala 75:16:@56710.4]
  assign regs_498_io_reset = reset; // @[RegFile.scala 78:19:@56714.4]
  assign regs_498_io_enable = 1'h1; // @[RegFile.scala 74:20:@56708.4]
  assign regs_499_clock = clock; // @[:@56717.4]
  assign regs_499_reset = io_reset; // @[:@56718.4 RegFile.scala 76:16:@56725.4]
  assign regs_499_io_in = 64'h0; // @[RegFile.scala 75:16:@56724.4]
  assign regs_499_io_reset = reset; // @[RegFile.scala 78:19:@56728.4]
  assign regs_499_io_enable = 1'h1; // @[RegFile.scala 74:20:@56722.4]
  assign regs_500_clock = clock; // @[:@56731.4]
  assign regs_500_reset = io_reset; // @[:@56732.4 RegFile.scala 76:16:@56739.4]
  assign regs_500_io_in = 64'h0; // @[RegFile.scala 75:16:@56738.4]
  assign regs_500_io_reset = reset; // @[RegFile.scala 78:19:@56742.4]
  assign regs_500_io_enable = 1'h1; // @[RegFile.scala 74:20:@56736.4]
  assign regs_501_clock = clock; // @[:@56745.4]
  assign regs_501_reset = io_reset; // @[:@56746.4 RegFile.scala 76:16:@56753.4]
  assign regs_501_io_in = 64'h0; // @[RegFile.scala 75:16:@56752.4]
  assign regs_501_io_reset = reset; // @[RegFile.scala 78:19:@56756.4]
  assign regs_501_io_enable = 1'h1; // @[RegFile.scala 74:20:@56750.4]
  assign regs_502_clock = clock; // @[:@56759.4]
  assign regs_502_reset = io_reset; // @[:@56760.4 RegFile.scala 76:16:@56767.4]
  assign regs_502_io_in = 64'h0; // @[RegFile.scala 75:16:@56766.4]
  assign regs_502_io_reset = reset; // @[RegFile.scala 78:19:@56770.4]
  assign regs_502_io_enable = 1'h1; // @[RegFile.scala 74:20:@56764.4]
  assign regs_503_clock = clock; // @[:@56773.4]
  assign regs_503_reset = io_reset; // @[:@56774.4 RegFile.scala 76:16:@56781.4]
  assign regs_503_io_in = 64'h0; // @[RegFile.scala 75:16:@56780.4]
  assign regs_503_io_reset = reset; // @[RegFile.scala 78:19:@56784.4]
  assign regs_503_io_enable = 1'h1; // @[RegFile.scala 74:20:@56778.4]
  assign regs_504_clock = clock; // @[:@56787.4]
  assign regs_504_reset = io_reset; // @[:@56788.4 RegFile.scala 76:16:@56795.4]
  assign regs_504_io_in = 64'h0; // @[RegFile.scala 75:16:@56794.4]
  assign regs_504_io_reset = reset; // @[RegFile.scala 78:19:@56798.4]
  assign regs_504_io_enable = 1'h1; // @[RegFile.scala 74:20:@56792.4]
  assign regs_505_clock = clock; // @[:@56801.4]
  assign regs_505_reset = io_reset; // @[:@56802.4 RegFile.scala 76:16:@56809.4]
  assign regs_505_io_in = 64'h0; // @[RegFile.scala 75:16:@56808.4]
  assign regs_505_io_reset = reset; // @[RegFile.scala 78:19:@56812.4]
  assign regs_505_io_enable = 1'h1; // @[RegFile.scala 74:20:@56806.4]
  assign regs_506_clock = clock; // @[:@56815.4]
  assign regs_506_reset = io_reset; // @[:@56816.4 RegFile.scala 76:16:@56823.4]
  assign regs_506_io_in = 64'h0; // @[RegFile.scala 75:16:@56822.4]
  assign regs_506_io_reset = reset; // @[RegFile.scala 78:19:@56826.4]
  assign regs_506_io_enable = 1'h1; // @[RegFile.scala 74:20:@56820.4]
  assign regs_507_clock = clock; // @[:@56829.4]
  assign regs_507_reset = io_reset; // @[:@56830.4 RegFile.scala 76:16:@56837.4]
  assign regs_507_io_in = 64'h0; // @[RegFile.scala 75:16:@56836.4]
  assign regs_507_io_reset = reset; // @[RegFile.scala 78:19:@56840.4]
  assign regs_507_io_enable = 1'h1; // @[RegFile.scala 74:20:@56834.4]
  assign regs_508_clock = clock; // @[:@56843.4]
  assign regs_508_reset = io_reset; // @[:@56844.4 RegFile.scala 76:16:@56851.4]
  assign regs_508_io_in = 64'h0; // @[RegFile.scala 75:16:@56850.4]
  assign regs_508_io_reset = reset; // @[RegFile.scala 78:19:@56854.4]
  assign regs_508_io_enable = 1'h1; // @[RegFile.scala 74:20:@56848.4]
  assign regs_509_clock = clock; // @[:@56857.4]
  assign regs_509_reset = io_reset; // @[:@56858.4 RegFile.scala 76:16:@56865.4]
  assign regs_509_io_in = 64'h0; // @[RegFile.scala 75:16:@56864.4]
  assign regs_509_io_reset = reset; // @[RegFile.scala 78:19:@56868.4]
  assign regs_509_io_enable = 1'h1; // @[RegFile.scala 74:20:@56862.4]
  assign regs_510_clock = clock; // @[:@56871.4]
  assign regs_510_reset = io_reset; // @[:@56872.4 RegFile.scala 76:16:@56879.4]
  assign regs_510_io_in = 64'h0; // @[RegFile.scala 75:16:@56878.4]
  assign regs_510_io_reset = reset; // @[RegFile.scala 78:19:@56882.4]
  assign regs_510_io_enable = 1'h1; // @[RegFile.scala 74:20:@56876.4]
  assign regs_511_clock = clock; // @[:@56885.4]
  assign regs_511_reset = io_reset; // @[:@56886.4 RegFile.scala 76:16:@56893.4]
  assign regs_511_io_in = 64'h0; // @[RegFile.scala 75:16:@56892.4]
  assign regs_511_io_reset = reset; // @[RegFile.scala 78:19:@56896.4]
  assign regs_511_io_enable = 1'h1; // @[RegFile.scala 74:20:@56890.4]
  assign regs_512_clock = clock; // @[:@56899.4]
  assign regs_512_reset = io_reset; // @[:@56900.4 RegFile.scala 76:16:@56907.4]
  assign regs_512_io_in = 64'h0; // @[RegFile.scala 75:16:@56906.4]
  assign regs_512_io_reset = reset; // @[RegFile.scala 78:19:@56910.4]
  assign regs_512_io_enable = 1'h1; // @[RegFile.scala 74:20:@56904.4]
  assign regs_513_clock = clock; // @[:@56913.4]
  assign regs_513_reset = io_reset; // @[:@56914.4 RegFile.scala 76:16:@56921.4]
  assign regs_513_io_in = 64'h0; // @[RegFile.scala 75:16:@56920.4]
  assign regs_513_io_reset = reset; // @[RegFile.scala 78:19:@56924.4]
  assign regs_513_io_enable = 1'h1; // @[RegFile.scala 74:20:@56918.4]
  assign regs_514_clock = clock; // @[:@56927.4]
  assign regs_514_reset = io_reset; // @[:@56928.4 RegFile.scala 76:16:@56935.4]
  assign regs_514_io_in = 64'h0; // @[RegFile.scala 75:16:@56934.4]
  assign regs_514_io_reset = reset; // @[RegFile.scala 78:19:@56938.4]
  assign regs_514_io_enable = 1'h1; // @[RegFile.scala 74:20:@56932.4]
  assign regs_515_clock = clock; // @[:@56941.4]
  assign regs_515_reset = io_reset; // @[:@56942.4 RegFile.scala 76:16:@56949.4]
  assign regs_515_io_in = 64'h0; // @[RegFile.scala 75:16:@56948.4]
  assign regs_515_io_reset = reset; // @[RegFile.scala 78:19:@56952.4]
  assign regs_515_io_enable = 1'h1; // @[RegFile.scala 74:20:@56946.4]
  assign regs_516_clock = clock; // @[:@56955.4]
  assign regs_516_reset = io_reset; // @[:@56956.4 RegFile.scala 76:16:@56963.4]
  assign regs_516_io_in = 64'h0; // @[RegFile.scala 75:16:@56962.4]
  assign regs_516_io_reset = reset; // @[RegFile.scala 78:19:@56966.4]
  assign regs_516_io_enable = 1'h1; // @[RegFile.scala 74:20:@56960.4]
  assign regs_517_clock = clock; // @[:@56969.4]
  assign regs_517_reset = io_reset; // @[:@56970.4 RegFile.scala 76:16:@56977.4]
  assign regs_517_io_in = 64'h0; // @[RegFile.scala 75:16:@56976.4]
  assign regs_517_io_reset = reset; // @[RegFile.scala 78:19:@56980.4]
  assign regs_517_io_enable = 1'h1; // @[RegFile.scala 74:20:@56974.4]
  assign rport_io_ins_0 = regs_0_io_out; // @[RegFile.scala 97:16:@57504.4]
  assign rport_io_ins_1 = regs_1_io_out; // @[RegFile.scala 97:16:@57505.4]
  assign rport_io_ins_2 = regs_2_io_out; // @[RegFile.scala 97:16:@57506.4]
  assign rport_io_ins_3 = regs_3_io_out; // @[RegFile.scala 97:16:@57507.4]
  assign rport_io_ins_4 = regs_4_io_out; // @[RegFile.scala 97:16:@57508.4]
  assign rport_io_ins_5 = regs_5_io_out; // @[RegFile.scala 97:16:@57509.4]
  assign rport_io_ins_6 = regs_6_io_out; // @[RegFile.scala 97:16:@57510.4]
  assign rport_io_ins_7 = regs_7_io_out; // @[RegFile.scala 97:16:@57511.4]
  assign rport_io_ins_8 = regs_8_io_out; // @[RegFile.scala 97:16:@57512.4]
  assign rport_io_ins_9 = regs_9_io_out; // @[RegFile.scala 97:16:@57513.4]
  assign rport_io_ins_10 = regs_10_io_out; // @[RegFile.scala 97:16:@57514.4]
  assign rport_io_ins_11 = regs_11_io_out; // @[RegFile.scala 97:16:@57515.4]
  assign rport_io_ins_12 = regs_12_io_out; // @[RegFile.scala 97:16:@57516.4]
  assign rport_io_ins_13 = regs_13_io_out; // @[RegFile.scala 97:16:@57517.4]
  assign rport_io_ins_14 = regs_14_io_out; // @[RegFile.scala 97:16:@57518.4]
  assign rport_io_ins_15 = regs_15_io_out; // @[RegFile.scala 97:16:@57519.4]
  assign rport_io_ins_16 = regs_16_io_out; // @[RegFile.scala 97:16:@57520.4]
  assign rport_io_ins_17 = regs_17_io_out; // @[RegFile.scala 97:16:@57521.4]
  assign rport_io_ins_18 = regs_18_io_out; // @[RegFile.scala 97:16:@57522.4]
  assign rport_io_ins_19 = regs_19_io_out; // @[RegFile.scala 97:16:@57523.4]
  assign rport_io_ins_20 = regs_20_io_out; // @[RegFile.scala 97:16:@57524.4]
  assign rport_io_ins_21 = regs_21_io_out; // @[RegFile.scala 97:16:@57525.4]
  assign rport_io_ins_22 = regs_22_io_out; // @[RegFile.scala 97:16:@57526.4]
  assign rport_io_ins_23 = regs_23_io_out; // @[RegFile.scala 97:16:@57527.4]
  assign rport_io_ins_24 = regs_24_io_out; // @[RegFile.scala 97:16:@57528.4]
  assign rport_io_ins_25 = regs_25_io_out; // @[RegFile.scala 97:16:@57529.4]
  assign rport_io_ins_26 = regs_26_io_out; // @[RegFile.scala 97:16:@57530.4]
  assign rport_io_ins_27 = regs_27_io_out; // @[RegFile.scala 97:16:@57531.4]
  assign rport_io_ins_28 = regs_28_io_out; // @[RegFile.scala 97:16:@57532.4]
  assign rport_io_ins_29 = regs_29_io_out; // @[RegFile.scala 97:16:@57533.4]
  assign rport_io_ins_30 = regs_30_io_out; // @[RegFile.scala 97:16:@57534.4]
  assign rport_io_ins_31 = regs_31_io_out; // @[RegFile.scala 97:16:@57535.4]
  assign rport_io_ins_32 = regs_32_io_out; // @[RegFile.scala 97:16:@57536.4]
  assign rport_io_ins_33 = regs_33_io_out; // @[RegFile.scala 97:16:@57537.4]
  assign rport_io_ins_34 = regs_34_io_out; // @[RegFile.scala 97:16:@57538.4]
  assign rport_io_ins_35 = regs_35_io_out; // @[RegFile.scala 97:16:@57539.4]
  assign rport_io_ins_36 = regs_36_io_out; // @[RegFile.scala 97:16:@57540.4]
  assign rport_io_ins_37 = regs_37_io_out; // @[RegFile.scala 97:16:@57541.4]
  assign rport_io_ins_38 = regs_38_io_out; // @[RegFile.scala 97:16:@57542.4]
  assign rport_io_ins_39 = regs_39_io_out; // @[RegFile.scala 97:16:@57543.4]
  assign rport_io_ins_40 = regs_40_io_out; // @[RegFile.scala 97:16:@57544.4]
  assign rport_io_ins_41 = regs_41_io_out; // @[RegFile.scala 97:16:@57545.4]
  assign rport_io_ins_42 = regs_42_io_out; // @[RegFile.scala 97:16:@57546.4]
  assign rport_io_ins_43 = regs_43_io_out; // @[RegFile.scala 97:16:@57547.4]
  assign rport_io_ins_44 = regs_44_io_out; // @[RegFile.scala 97:16:@57548.4]
  assign rport_io_ins_45 = regs_45_io_out; // @[RegFile.scala 97:16:@57549.4]
  assign rport_io_ins_46 = regs_46_io_out; // @[RegFile.scala 97:16:@57550.4]
  assign rport_io_ins_47 = regs_47_io_out; // @[RegFile.scala 97:16:@57551.4]
  assign rport_io_ins_48 = regs_48_io_out; // @[RegFile.scala 97:16:@57552.4]
  assign rport_io_ins_49 = regs_49_io_out; // @[RegFile.scala 97:16:@57553.4]
  assign rport_io_ins_50 = regs_50_io_out; // @[RegFile.scala 97:16:@57554.4]
  assign rport_io_ins_51 = regs_51_io_out; // @[RegFile.scala 97:16:@57555.4]
  assign rport_io_ins_52 = regs_52_io_out; // @[RegFile.scala 97:16:@57556.4]
  assign rport_io_ins_53 = regs_53_io_out; // @[RegFile.scala 97:16:@57557.4]
  assign rport_io_ins_54 = regs_54_io_out; // @[RegFile.scala 97:16:@57558.4]
  assign rport_io_ins_55 = regs_55_io_out; // @[RegFile.scala 97:16:@57559.4]
  assign rport_io_ins_56 = regs_56_io_out; // @[RegFile.scala 97:16:@57560.4]
  assign rport_io_ins_57 = regs_57_io_out; // @[RegFile.scala 97:16:@57561.4]
  assign rport_io_ins_58 = regs_58_io_out; // @[RegFile.scala 97:16:@57562.4]
  assign rport_io_ins_59 = regs_59_io_out; // @[RegFile.scala 97:16:@57563.4]
  assign rport_io_ins_60 = regs_60_io_out; // @[RegFile.scala 97:16:@57564.4]
  assign rport_io_ins_61 = regs_61_io_out; // @[RegFile.scala 97:16:@57565.4]
  assign rport_io_ins_62 = regs_62_io_out; // @[RegFile.scala 97:16:@57566.4]
  assign rport_io_ins_63 = regs_63_io_out; // @[RegFile.scala 97:16:@57567.4]
  assign rport_io_ins_64 = regs_64_io_out; // @[RegFile.scala 97:16:@57568.4]
  assign rport_io_ins_65 = regs_65_io_out; // @[RegFile.scala 97:16:@57569.4]
  assign rport_io_ins_66 = regs_66_io_out; // @[RegFile.scala 97:16:@57570.4]
  assign rport_io_ins_67 = regs_67_io_out; // @[RegFile.scala 97:16:@57571.4]
  assign rport_io_ins_68 = regs_68_io_out; // @[RegFile.scala 97:16:@57572.4]
  assign rport_io_ins_69 = regs_69_io_out; // @[RegFile.scala 97:16:@57573.4]
  assign rport_io_ins_70 = regs_70_io_out; // @[RegFile.scala 97:16:@57574.4]
  assign rport_io_ins_71 = regs_71_io_out; // @[RegFile.scala 97:16:@57575.4]
  assign rport_io_ins_72 = regs_72_io_out; // @[RegFile.scala 97:16:@57576.4]
  assign rport_io_ins_73 = regs_73_io_out; // @[RegFile.scala 97:16:@57577.4]
  assign rport_io_ins_74 = regs_74_io_out; // @[RegFile.scala 97:16:@57578.4]
  assign rport_io_ins_75 = regs_75_io_out; // @[RegFile.scala 97:16:@57579.4]
  assign rport_io_ins_76 = regs_76_io_out; // @[RegFile.scala 97:16:@57580.4]
  assign rport_io_ins_77 = regs_77_io_out; // @[RegFile.scala 97:16:@57581.4]
  assign rport_io_ins_78 = regs_78_io_out; // @[RegFile.scala 97:16:@57582.4]
  assign rport_io_ins_79 = regs_79_io_out; // @[RegFile.scala 97:16:@57583.4]
  assign rport_io_ins_80 = regs_80_io_out; // @[RegFile.scala 97:16:@57584.4]
  assign rport_io_ins_81 = regs_81_io_out; // @[RegFile.scala 97:16:@57585.4]
  assign rport_io_ins_82 = regs_82_io_out; // @[RegFile.scala 97:16:@57586.4]
  assign rport_io_ins_83 = regs_83_io_out; // @[RegFile.scala 97:16:@57587.4]
  assign rport_io_ins_84 = regs_84_io_out; // @[RegFile.scala 97:16:@57588.4]
  assign rport_io_ins_85 = regs_85_io_out; // @[RegFile.scala 97:16:@57589.4]
  assign rport_io_ins_86 = regs_86_io_out; // @[RegFile.scala 97:16:@57590.4]
  assign rport_io_ins_87 = regs_87_io_out; // @[RegFile.scala 97:16:@57591.4]
  assign rport_io_ins_88 = regs_88_io_out; // @[RegFile.scala 97:16:@57592.4]
  assign rport_io_ins_89 = regs_89_io_out; // @[RegFile.scala 97:16:@57593.4]
  assign rport_io_ins_90 = regs_90_io_out; // @[RegFile.scala 97:16:@57594.4]
  assign rport_io_ins_91 = regs_91_io_out; // @[RegFile.scala 97:16:@57595.4]
  assign rport_io_ins_92 = regs_92_io_out; // @[RegFile.scala 97:16:@57596.4]
  assign rport_io_ins_93 = regs_93_io_out; // @[RegFile.scala 97:16:@57597.4]
  assign rport_io_ins_94 = regs_94_io_out; // @[RegFile.scala 97:16:@57598.4]
  assign rport_io_ins_95 = regs_95_io_out; // @[RegFile.scala 97:16:@57599.4]
  assign rport_io_ins_96 = regs_96_io_out; // @[RegFile.scala 97:16:@57600.4]
  assign rport_io_ins_97 = regs_97_io_out; // @[RegFile.scala 97:16:@57601.4]
  assign rport_io_ins_98 = regs_98_io_out; // @[RegFile.scala 97:16:@57602.4]
  assign rport_io_ins_99 = regs_99_io_out; // @[RegFile.scala 97:16:@57603.4]
  assign rport_io_ins_100 = regs_100_io_out; // @[RegFile.scala 97:16:@57604.4]
  assign rport_io_ins_101 = regs_101_io_out; // @[RegFile.scala 97:16:@57605.4]
  assign rport_io_ins_102 = regs_102_io_out; // @[RegFile.scala 97:16:@57606.4]
  assign rport_io_ins_103 = regs_103_io_out; // @[RegFile.scala 97:16:@57607.4]
  assign rport_io_ins_104 = regs_104_io_out; // @[RegFile.scala 97:16:@57608.4]
  assign rport_io_ins_105 = regs_105_io_out; // @[RegFile.scala 97:16:@57609.4]
  assign rport_io_ins_106 = regs_106_io_out; // @[RegFile.scala 97:16:@57610.4]
  assign rport_io_ins_107 = regs_107_io_out; // @[RegFile.scala 97:16:@57611.4]
  assign rport_io_ins_108 = regs_108_io_out; // @[RegFile.scala 97:16:@57612.4]
  assign rport_io_ins_109 = regs_109_io_out; // @[RegFile.scala 97:16:@57613.4]
  assign rport_io_ins_110 = regs_110_io_out; // @[RegFile.scala 97:16:@57614.4]
  assign rport_io_ins_111 = regs_111_io_out; // @[RegFile.scala 97:16:@57615.4]
  assign rport_io_ins_112 = regs_112_io_out; // @[RegFile.scala 97:16:@57616.4]
  assign rport_io_ins_113 = regs_113_io_out; // @[RegFile.scala 97:16:@57617.4]
  assign rport_io_ins_114 = regs_114_io_out; // @[RegFile.scala 97:16:@57618.4]
  assign rport_io_ins_115 = regs_115_io_out; // @[RegFile.scala 97:16:@57619.4]
  assign rport_io_ins_116 = regs_116_io_out; // @[RegFile.scala 97:16:@57620.4]
  assign rport_io_ins_117 = regs_117_io_out; // @[RegFile.scala 97:16:@57621.4]
  assign rport_io_ins_118 = regs_118_io_out; // @[RegFile.scala 97:16:@57622.4]
  assign rport_io_ins_119 = regs_119_io_out; // @[RegFile.scala 97:16:@57623.4]
  assign rport_io_ins_120 = regs_120_io_out; // @[RegFile.scala 97:16:@57624.4]
  assign rport_io_ins_121 = regs_121_io_out; // @[RegFile.scala 97:16:@57625.4]
  assign rport_io_ins_122 = regs_122_io_out; // @[RegFile.scala 97:16:@57626.4]
  assign rport_io_ins_123 = regs_123_io_out; // @[RegFile.scala 97:16:@57627.4]
  assign rport_io_ins_124 = regs_124_io_out; // @[RegFile.scala 97:16:@57628.4]
  assign rport_io_ins_125 = regs_125_io_out; // @[RegFile.scala 97:16:@57629.4]
  assign rport_io_ins_126 = regs_126_io_out; // @[RegFile.scala 97:16:@57630.4]
  assign rport_io_ins_127 = regs_127_io_out; // @[RegFile.scala 97:16:@57631.4]
  assign rport_io_ins_128 = regs_128_io_out; // @[RegFile.scala 97:16:@57632.4]
  assign rport_io_ins_129 = regs_129_io_out; // @[RegFile.scala 97:16:@57633.4]
  assign rport_io_ins_130 = regs_130_io_out; // @[RegFile.scala 97:16:@57634.4]
  assign rport_io_ins_131 = regs_131_io_out; // @[RegFile.scala 97:16:@57635.4]
  assign rport_io_ins_132 = regs_132_io_out; // @[RegFile.scala 97:16:@57636.4]
  assign rport_io_ins_133 = regs_133_io_out; // @[RegFile.scala 97:16:@57637.4]
  assign rport_io_ins_134 = regs_134_io_out; // @[RegFile.scala 97:16:@57638.4]
  assign rport_io_ins_135 = regs_135_io_out; // @[RegFile.scala 97:16:@57639.4]
  assign rport_io_ins_136 = regs_136_io_out; // @[RegFile.scala 97:16:@57640.4]
  assign rport_io_ins_137 = regs_137_io_out; // @[RegFile.scala 97:16:@57641.4]
  assign rport_io_ins_138 = regs_138_io_out; // @[RegFile.scala 97:16:@57642.4]
  assign rport_io_ins_139 = regs_139_io_out; // @[RegFile.scala 97:16:@57643.4]
  assign rport_io_ins_140 = regs_140_io_out; // @[RegFile.scala 97:16:@57644.4]
  assign rport_io_ins_141 = regs_141_io_out; // @[RegFile.scala 97:16:@57645.4]
  assign rport_io_ins_142 = regs_142_io_out; // @[RegFile.scala 97:16:@57646.4]
  assign rport_io_ins_143 = regs_143_io_out; // @[RegFile.scala 97:16:@57647.4]
  assign rport_io_ins_144 = regs_144_io_out; // @[RegFile.scala 97:16:@57648.4]
  assign rport_io_ins_145 = regs_145_io_out; // @[RegFile.scala 97:16:@57649.4]
  assign rport_io_ins_146 = regs_146_io_out; // @[RegFile.scala 97:16:@57650.4]
  assign rport_io_ins_147 = regs_147_io_out; // @[RegFile.scala 97:16:@57651.4]
  assign rport_io_ins_148 = regs_148_io_out; // @[RegFile.scala 97:16:@57652.4]
  assign rport_io_ins_149 = regs_149_io_out; // @[RegFile.scala 97:16:@57653.4]
  assign rport_io_ins_150 = regs_150_io_out; // @[RegFile.scala 97:16:@57654.4]
  assign rport_io_ins_151 = regs_151_io_out; // @[RegFile.scala 97:16:@57655.4]
  assign rport_io_ins_152 = regs_152_io_out; // @[RegFile.scala 97:16:@57656.4]
  assign rport_io_ins_153 = regs_153_io_out; // @[RegFile.scala 97:16:@57657.4]
  assign rport_io_ins_154 = regs_154_io_out; // @[RegFile.scala 97:16:@57658.4]
  assign rport_io_ins_155 = regs_155_io_out; // @[RegFile.scala 97:16:@57659.4]
  assign rport_io_ins_156 = regs_156_io_out; // @[RegFile.scala 97:16:@57660.4]
  assign rport_io_ins_157 = regs_157_io_out; // @[RegFile.scala 97:16:@57661.4]
  assign rport_io_ins_158 = regs_158_io_out; // @[RegFile.scala 97:16:@57662.4]
  assign rport_io_ins_159 = regs_159_io_out; // @[RegFile.scala 97:16:@57663.4]
  assign rport_io_ins_160 = regs_160_io_out; // @[RegFile.scala 97:16:@57664.4]
  assign rport_io_ins_161 = regs_161_io_out; // @[RegFile.scala 97:16:@57665.4]
  assign rport_io_ins_162 = regs_162_io_out; // @[RegFile.scala 97:16:@57666.4]
  assign rport_io_ins_163 = regs_163_io_out; // @[RegFile.scala 97:16:@57667.4]
  assign rport_io_ins_164 = regs_164_io_out; // @[RegFile.scala 97:16:@57668.4]
  assign rport_io_ins_165 = regs_165_io_out; // @[RegFile.scala 97:16:@57669.4]
  assign rport_io_ins_166 = regs_166_io_out; // @[RegFile.scala 97:16:@57670.4]
  assign rport_io_ins_167 = regs_167_io_out; // @[RegFile.scala 97:16:@57671.4]
  assign rport_io_ins_168 = regs_168_io_out; // @[RegFile.scala 97:16:@57672.4]
  assign rport_io_ins_169 = regs_169_io_out; // @[RegFile.scala 97:16:@57673.4]
  assign rport_io_ins_170 = regs_170_io_out; // @[RegFile.scala 97:16:@57674.4]
  assign rport_io_ins_171 = regs_171_io_out; // @[RegFile.scala 97:16:@57675.4]
  assign rport_io_ins_172 = regs_172_io_out; // @[RegFile.scala 97:16:@57676.4]
  assign rport_io_ins_173 = regs_173_io_out; // @[RegFile.scala 97:16:@57677.4]
  assign rport_io_ins_174 = regs_174_io_out; // @[RegFile.scala 97:16:@57678.4]
  assign rport_io_ins_175 = regs_175_io_out; // @[RegFile.scala 97:16:@57679.4]
  assign rport_io_ins_176 = regs_176_io_out; // @[RegFile.scala 97:16:@57680.4]
  assign rport_io_ins_177 = regs_177_io_out; // @[RegFile.scala 97:16:@57681.4]
  assign rport_io_ins_178 = regs_178_io_out; // @[RegFile.scala 97:16:@57682.4]
  assign rport_io_ins_179 = regs_179_io_out; // @[RegFile.scala 97:16:@57683.4]
  assign rport_io_ins_180 = regs_180_io_out; // @[RegFile.scala 97:16:@57684.4]
  assign rport_io_ins_181 = regs_181_io_out; // @[RegFile.scala 97:16:@57685.4]
  assign rport_io_ins_182 = regs_182_io_out; // @[RegFile.scala 97:16:@57686.4]
  assign rport_io_ins_183 = regs_183_io_out; // @[RegFile.scala 97:16:@57687.4]
  assign rport_io_ins_184 = regs_184_io_out; // @[RegFile.scala 97:16:@57688.4]
  assign rport_io_ins_185 = regs_185_io_out; // @[RegFile.scala 97:16:@57689.4]
  assign rport_io_ins_186 = regs_186_io_out; // @[RegFile.scala 97:16:@57690.4]
  assign rport_io_ins_187 = regs_187_io_out; // @[RegFile.scala 97:16:@57691.4]
  assign rport_io_ins_188 = regs_188_io_out; // @[RegFile.scala 97:16:@57692.4]
  assign rport_io_ins_189 = regs_189_io_out; // @[RegFile.scala 97:16:@57693.4]
  assign rport_io_ins_190 = regs_190_io_out; // @[RegFile.scala 97:16:@57694.4]
  assign rport_io_ins_191 = regs_191_io_out; // @[RegFile.scala 97:16:@57695.4]
  assign rport_io_ins_192 = regs_192_io_out; // @[RegFile.scala 97:16:@57696.4]
  assign rport_io_ins_193 = regs_193_io_out; // @[RegFile.scala 97:16:@57697.4]
  assign rport_io_ins_194 = regs_194_io_out; // @[RegFile.scala 97:16:@57698.4]
  assign rport_io_ins_195 = regs_195_io_out; // @[RegFile.scala 97:16:@57699.4]
  assign rport_io_ins_196 = regs_196_io_out; // @[RegFile.scala 97:16:@57700.4]
  assign rport_io_ins_197 = regs_197_io_out; // @[RegFile.scala 97:16:@57701.4]
  assign rport_io_ins_198 = regs_198_io_out; // @[RegFile.scala 97:16:@57702.4]
  assign rport_io_ins_199 = regs_199_io_out; // @[RegFile.scala 97:16:@57703.4]
  assign rport_io_ins_200 = regs_200_io_out; // @[RegFile.scala 97:16:@57704.4]
  assign rport_io_ins_201 = regs_201_io_out; // @[RegFile.scala 97:16:@57705.4]
  assign rport_io_ins_202 = regs_202_io_out; // @[RegFile.scala 97:16:@57706.4]
  assign rport_io_ins_203 = regs_203_io_out; // @[RegFile.scala 97:16:@57707.4]
  assign rport_io_ins_204 = regs_204_io_out; // @[RegFile.scala 97:16:@57708.4]
  assign rport_io_ins_205 = regs_205_io_out; // @[RegFile.scala 97:16:@57709.4]
  assign rport_io_ins_206 = regs_206_io_out; // @[RegFile.scala 97:16:@57710.4]
  assign rport_io_ins_207 = regs_207_io_out; // @[RegFile.scala 97:16:@57711.4]
  assign rport_io_ins_208 = regs_208_io_out; // @[RegFile.scala 97:16:@57712.4]
  assign rport_io_ins_209 = regs_209_io_out; // @[RegFile.scala 97:16:@57713.4]
  assign rport_io_ins_210 = regs_210_io_out; // @[RegFile.scala 97:16:@57714.4]
  assign rport_io_ins_211 = regs_211_io_out; // @[RegFile.scala 97:16:@57715.4]
  assign rport_io_ins_212 = regs_212_io_out; // @[RegFile.scala 97:16:@57716.4]
  assign rport_io_ins_213 = regs_213_io_out; // @[RegFile.scala 97:16:@57717.4]
  assign rport_io_ins_214 = regs_214_io_out; // @[RegFile.scala 97:16:@57718.4]
  assign rport_io_ins_215 = regs_215_io_out; // @[RegFile.scala 97:16:@57719.4]
  assign rport_io_ins_216 = regs_216_io_out; // @[RegFile.scala 97:16:@57720.4]
  assign rport_io_ins_217 = regs_217_io_out; // @[RegFile.scala 97:16:@57721.4]
  assign rport_io_ins_218 = regs_218_io_out; // @[RegFile.scala 97:16:@57722.4]
  assign rport_io_ins_219 = regs_219_io_out; // @[RegFile.scala 97:16:@57723.4]
  assign rport_io_ins_220 = regs_220_io_out; // @[RegFile.scala 97:16:@57724.4]
  assign rport_io_ins_221 = regs_221_io_out; // @[RegFile.scala 97:16:@57725.4]
  assign rport_io_ins_222 = regs_222_io_out; // @[RegFile.scala 97:16:@57726.4]
  assign rport_io_ins_223 = regs_223_io_out; // @[RegFile.scala 97:16:@57727.4]
  assign rport_io_ins_224 = regs_224_io_out; // @[RegFile.scala 97:16:@57728.4]
  assign rport_io_ins_225 = regs_225_io_out; // @[RegFile.scala 97:16:@57729.4]
  assign rport_io_ins_226 = regs_226_io_out; // @[RegFile.scala 97:16:@57730.4]
  assign rport_io_ins_227 = regs_227_io_out; // @[RegFile.scala 97:16:@57731.4]
  assign rport_io_ins_228 = regs_228_io_out; // @[RegFile.scala 97:16:@57732.4]
  assign rport_io_ins_229 = regs_229_io_out; // @[RegFile.scala 97:16:@57733.4]
  assign rport_io_ins_230 = regs_230_io_out; // @[RegFile.scala 97:16:@57734.4]
  assign rport_io_ins_231 = regs_231_io_out; // @[RegFile.scala 97:16:@57735.4]
  assign rport_io_ins_232 = regs_232_io_out; // @[RegFile.scala 97:16:@57736.4]
  assign rport_io_ins_233 = regs_233_io_out; // @[RegFile.scala 97:16:@57737.4]
  assign rport_io_ins_234 = regs_234_io_out; // @[RegFile.scala 97:16:@57738.4]
  assign rport_io_ins_235 = regs_235_io_out; // @[RegFile.scala 97:16:@57739.4]
  assign rport_io_ins_236 = regs_236_io_out; // @[RegFile.scala 97:16:@57740.4]
  assign rport_io_ins_237 = regs_237_io_out; // @[RegFile.scala 97:16:@57741.4]
  assign rport_io_ins_238 = regs_238_io_out; // @[RegFile.scala 97:16:@57742.4]
  assign rport_io_ins_239 = regs_239_io_out; // @[RegFile.scala 97:16:@57743.4]
  assign rport_io_ins_240 = regs_240_io_out; // @[RegFile.scala 97:16:@57744.4]
  assign rport_io_ins_241 = regs_241_io_out; // @[RegFile.scala 97:16:@57745.4]
  assign rport_io_ins_242 = regs_242_io_out; // @[RegFile.scala 97:16:@57746.4]
  assign rport_io_ins_243 = regs_243_io_out; // @[RegFile.scala 97:16:@57747.4]
  assign rport_io_ins_244 = regs_244_io_out; // @[RegFile.scala 97:16:@57748.4]
  assign rport_io_ins_245 = regs_245_io_out; // @[RegFile.scala 97:16:@57749.4]
  assign rport_io_ins_246 = regs_246_io_out; // @[RegFile.scala 97:16:@57750.4]
  assign rport_io_ins_247 = regs_247_io_out; // @[RegFile.scala 97:16:@57751.4]
  assign rport_io_ins_248 = regs_248_io_out; // @[RegFile.scala 97:16:@57752.4]
  assign rport_io_ins_249 = regs_249_io_out; // @[RegFile.scala 97:16:@57753.4]
  assign rport_io_ins_250 = regs_250_io_out; // @[RegFile.scala 97:16:@57754.4]
  assign rport_io_ins_251 = regs_251_io_out; // @[RegFile.scala 97:16:@57755.4]
  assign rport_io_ins_252 = regs_252_io_out; // @[RegFile.scala 97:16:@57756.4]
  assign rport_io_ins_253 = regs_253_io_out; // @[RegFile.scala 97:16:@57757.4]
  assign rport_io_ins_254 = regs_254_io_out; // @[RegFile.scala 97:16:@57758.4]
  assign rport_io_ins_255 = regs_255_io_out; // @[RegFile.scala 97:16:@57759.4]
  assign rport_io_ins_256 = regs_256_io_out; // @[RegFile.scala 97:16:@57760.4]
  assign rport_io_ins_257 = regs_257_io_out; // @[RegFile.scala 97:16:@57761.4]
  assign rport_io_ins_258 = regs_258_io_out; // @[RegFile.scala 97:16:@57762.4]
  assign rport_io_ins_259 = regs_259_io_out; // @[RegFile.scala 97:16:@57763.4]
  assign rport_io_ins_260 = regs_260_io_out; // @[RegFile.scala 97:16:@57764.4]
  assign rport_io_ins_261 = regs_261_io_out; // @[RegFile.scala 97:16:@57765.4]
  assign rport_io_ins_262 = regs_262_io_out; // @[RegFile.scala 97:16:@57766.4]
  assign rport_io_ins_263 = regs_263_io_out; // @[RegFile.scala 97:16:@57767.4]
  assign rport_io_ins_264 = regs_264_io_out; // @[RegFile.scala 97:16:@57768.4]
  assign rport_io_ins_265 = regs_265_io_out; // @[RegFile.scala 97:16:@57769.4]
  assign rport_io_ins_266 = regs_266_io_out; // @[RegFile.scala 97:16:@57770.4]
  assign rport_io_ins_267 = regs_267_io_out; // @[RegFile.scala 97:16:@57771.4]
  assign rport_io_ins_268 = regs_268_io_out; // @[RegFile.scala 97:16:@57772.4]
  assign rport_io_ins_269 = regs_269_io_out; // @[RegFile.scala 97:16:@57773.4]
  assign rport_io_ins_270 = regs_270_io_out; // @[RegFile.scala 97:16:@57774.4]
  assign rport_io_ins_271 = regs_271_io_out; // @[RegFile.scala 97:16:@57775.4]
  assign rport_io_ins_272 = regs_272_io_out; // @[RegFile.scala 97:16:@57776.4]
  assign rport_io_ins_273 = regs_273_io_out; // @[RegFile.scala 97:16:@57777.4]
  assign rport_io_ins_274 = regs_274_io_out; // @[RegFile.scala 97:16:@57778.4]
  assign rport_io_ins_275 = regs_275_io_out; // @[RegFile.scala 97:16:@57779.4]
  assign rport_io_ins_276 = regs_276_io_out; // @[RegFile.scala 97:16:@57780.4]
  assign rport_io_ins_277 = regs_277_io_out; // @[RegFile.scala 97:16:@57781.4]
  assign rport_io_ins_278 = regs_278_io_out; // @[RegFile.scala 97:16:@57782.4]
  assign rport_io_ins_279 = regs_279_io_out; // @[RegFile.scala 97:16:@57783.4]
  assign rport_io_ins_280 = regs_280_io_out; // @[RegFile.scala 97:16:@57784.4]
  assign rport_io_ins_281 = regs_281_io_out; // @[RegFile.scala 97:16:@57785.4]
  assign rport_io_ins_282 = regs_282_io_out; // @[RegFile.scala 97:16:@57786.4]
  assign rport_io_ins_283 = regs_283_io_out; // @[RegFile.scala 97:16:@57787.4]
  assign rport_io_ins_284 = regs_284_io_out; // @[RegFile.scala 97:16:@57788.4]
  assign rport_io_ins_285 = regs_285_io_out; // @[RegFile.scala 97:16:@57789.4]
  assign rport_io_ins_286 = regs_286_io_out; // @[RegFile.scala 97:16:@57790.4]
  assign rport_io_ins_287 = regs_287_io_out; // @[RegFile.scala 97:16:@57791.4]
  assign rport_io_ins_288 = regs_288_io_out; // @[RegFile.scala 97:16:@57792.4]
  assign rport_io_ins_289 = regs_289_io_out; // @[RegFile.scala 97:16:@57793.4]
  assign rport_io_ins_290 = regs_290_io_out; // @[RegFile.scala 97:16:@57794.4]
  assign rport_io_ins_291 = regs_291_io_out; // @[RegFile.scala 97:16:@57795.4]
  assign rport_io_ins_292 = regs_292_io_out; // @[RegFile.scala 97:16:@57796.4]
  assign rport_io_ins_293 = regs_293_io_out; // @[RegFile.scala 97:16:@57797.4]
  assign rport_io_ins_294 = regs_294_io_out; // @[RegFile.scala 97:16:@57798.4]
  assign rport_io_ins_295 = regs_295_io_out; // @[RegFile.scala 97:16:@57799.4]
  assign rport_io_ins_296 = regs_296_io_out; // @[RegFile.scala 97:16:@57800.4]
  assign rport_io_ins_297 = regs_297_io_out; // @[RegFile.scala 97:16:@57801.4]
  assign rport_io_ins_298 = regs_298_io_out; // @[RegFile.scala 97:16:@57802.4]
  assign rport_io_ins_299 = regs_299_io_out; // @[RegFile.scala 97:16:@57803.4]
  assign rport_io_ins_300 = regs_300_io_out; // @[RegFile.scala 97:16:@57804.4]
  assign rport_io_ins_301 = regs_301_io_out; // @[RegFile.scala 97:16:@57805.4]
  assign rport_io_ins_302 = regs_302_io_out; // @[RegFile.scala 97:16:@57806.4]
  assign rport_io_ins_303 = regs_303_io_out; // @[RegFile.scala 97:16:@57807.4]
  assign rport_io_ins_304 = regs_304_io_out; // @[RegFile.scala 97:16:@57808.4]
  assign rport_io_ins_305 = regs_305_io_out; // @[RegFile.scala 97:16:@57809.4]
  assign rport_io_ins_306 = regs_306_io_out; // @[RegFile.scala 97:16:@57810.4]
  assign rport_io_ins_307 = regs_307_io_out; // @[RegFile.scala 97:16:@57811.4]
  assign rport_io_ins_308 = regs_308_io_out; // @[RegFile.scala 97:16:@57812.4]
  assign rport_io_ins_309 = regs_309_io_out; // @[RegFile.scala 97:16:@57813.4]
  assign rport_io_ins_310 = regs_310_io_out; // @[RegFile.scala 97:16:@57814.4]
  assign rport_io_ins_311 = regs_311_io_out; // @[RegFile.scala 97:16:@57815.4]
  assign rport_io_ins_312 = regs_312_io_out; // @[RegFile.scala 97:16:@57816.4]
  assign rport_io_ins_313 = regs_313_io_out; // @[RegFile.scala 97:16:@57817.4]
  assign rport_io_ins_314 = regs_314_io_out; // @[RegFile.scala 97:16:@57818.4]
  assign rport_io_ins_315 = regs_315_io_out; // @[RegFile.scala 97:16:@57819.4]
  assign rport_io_ins_316 = regs_316_io_out; // @[RegFile.scala 97:16:@57820.4]
  assign rport_io_ins_317 = regs_317_io_out; // @[RegFile.scala 97:16:@57821.4]
  assign rport_io_ins_318 = regs_318_io_out; // @[RegFile.scala 97:16:@57822.4]
  assign rport_io_ins_319 = regs_319_io_out; // @[RegFile.scala 97:16:@57823.4]
  assign rport_io_ins_320 = regs_320_io_out; // @[RegFile.scala 97:16:@57824.4]
  assign rport_io_ins_321 = regs_321_io_out; // @[RegFile.scala 97:16:@57825.4]
  assign rport_io_ins_322 = regs_322_io_out; // @[RegFile.scala 97:16:@57826.4]
  assign rport_io_ins_323 = regs_323_io_out; // @[RegFile.scala 97:16:@57827.4]
  assign rport_io_ins_324 = regs_324_io_out; // @[RegFile.scala 97:16:@57828.4]
  assign rport_io_ins_325 = regs_325_io_out; // @[RegFile.scala 97:16:@57829.4]
  assign rport_io_ins_326 = regs_326_io_out; // @[RegFile.scala 97:16:@57830.4]
  assign rport_io_ins_327 = regs_327_io_out; // @[RegFile.scala 97:16:@57831.4]
  assign rport_io_ins_328 = regs_328_io_out; // @[RegFile.scala 97:16:@57832.4]
  assign rport_io_ins_329 = regs_329_io_out; // @[RegFile.scala 97:16:@57833.4]
  assign rport_io_ins_330 = regs_330_io_out; // @[RegFile.scala 97:16:@57834.4]
  assign rport_io_ins_331 = regs_331_io_out; // @[RegFile.scala 97:16:@57835.4]
  assign rport_io_ins_332 = regs_332_io_out; // @[RegFile.scala 97:16:@57836.4]
  assign rport_io_ins_333 = regs_333_io_out; // @[RegFile.scala 97:16:@57837.4]
  assign rport_io_ins_334 = regs_334_io_out; // @[RegFile.scala 97:16:@57838.4]
  assign rport_io_ins_335 = regs_335_io_out; // @[RegFile.scala 97:16:@57839.4]
  assign rport_io_ins_336 = regs_336_io_out; // @[RegFile.scala 97:16:@57840.4]
  assign rport_io_ins_337 = regs_337_io_out; // @[RegFile.scala 97:16:@57841.4]
  assign rport_io_ins_338 = regs_338_io_out; // @[RegFile.scala 97:16:@57842.4]
  assign rport_io_ins_339 = regs_339_io_out; // @[RegFile.scala 97:16:@57843.4]
  assign rport_io_ins_340 = regs_340_io_out; // @[RegFile.scala 97:16:@57844.4]
  assign rport_io_ins_341 = regs_341_io_out; // @[RegFile.scala 97:16:@57845.4]
  assign rport_io_ins_342 = regs_342_io_out; // @[RegFile.scala 97:16:@57846.4]
  assign rport_io_ins_343 = regs_343_io_out; // @[RegFile.scala 97:16:@57847.4]
  assign rport_io_ins_344 = regs_344_io_out; // @[RegFile.scala 97:16:@57848.4]
  assign rport_io_ins_345 = regs_345_io_out; // @[RegFile.scala 97:16:@57849.4]
  assign rport_io_ins_346 = regs_346_io_out; // @[RegFile.scala 97:16:@57850.4]
  assign rport_io_ins_347 = regs_347_io_out; // @[RegFile.scala 97:16:@57851.4]
  assign rport_io_ins_348 = regs_348_io_out; // @[RegFile.scala 97:16:@57852.4]
  assign rport_io_ins_349 = regs_349_io_out; // @[RegFile.scala 97:16:@57853.4]
  assign rport_io_ins_350 = regs_350_io_out; // @[RegFile.scala 97:16:@57854.4]
  assign rport_io_ins_351 = regs_351_io_out; // @[RegFile.scala 97:16:@57855.4]
  assign rport_io_ins_352 = regs_352_io_out; // @[RegFile.scala 97:16:@57856.4]
  assign rport_io_ins_353 = regs_353_io_out; // @[RegFile.scala 97:16:@57857.4]
  assign rport_io_ins_354 = regs_354_io_out; // @[RegFile.scala 97:16:@57858.4]
  assign rport_io_ins_355 = regs_355_io_out; // @[RegFile.scala 97:16:@57859.4]
  assign rport_io_ins_356 = regs_356_io_out; // @[RegFile.scala 97:16:@57860.4]
  assign rport_io_ins_357 = regs_357_io_out; // @[RegFile.scala 97:16:@57861.4]
  assign rport_io_ins_358 = regs_358_io_out; // @[RegFile.scala 97:16:@57862.4]
  assign rport_io_ins_359 = regs_359_io_out; // @[RegFile.scala 97:16:@57863.4]
  assign rport_io_ins_360 = regs_360_io_out; // @[RegFile.scala 97:16:@57864.4]
  assign rport_io_ins_361 = regs_361_io_out; // @[RegFile.scala 97:16:@57865.4]
  assign rport_io_ins_362 = regs_362_io_out; // @[RegFile.scala 97:16:@57866.4]
  assign rport_io_ins_363 = regs_363_io_out; // @[RegFile.scala 97:16:@57867.4]
  assign rport_io_ins_364 = regs_364_io_out; // @[RegFile.scala 97:16:@57868.4]
  assign rport_io_ins_365 = regs_365_io_out; // @[RegFile.scala 97:16:@57869.4]
  assign rport_io_ins_366 = regs_366_io_out; // @[RegFile.scala 97:16:@57870.4]
  assign rport_io_ins_367 = regs_367_io_out; // @[RegFile.scala 97:16:@57871.4]
  assign rport_io_ins_368 = regs_368_io_out; // @[RegFile.scala 97:16:@57872.4]
  assign rport_io_ins_369 = regs_369_io_out; // @[RegFile.scala 97:16:@57873.4]
  assign rport_io_ins_370 = regs_370_io_out; // @[RegFile.scala 97:16:@57874.4]
  assign rport_io_ins_371 = regs_371_io_out; // @[RegFile.scala 97:16:@57875.4]
  assign rport_io_ins_372 = regs_372_io_out; // @[RegFile.scala 97:16:@57876.4]
  assign rport_io_ins_373 = regs_373_io_out; // @[RegFile.scala 97:16:@57877.4]
  assign rport_io_ins_374 = regs_374_io_out; // @[RegFile.scala 97:16:@57878.4]
  assign rport_io_ins_375 = regs_375_io_out; // @[RegFile.scala 97:16:@57879.4]
  assign rport_io_ins_376 = regs_376_io_out; // @[RegFile.scala 97:16:@57880.4]
  assign rport_io_ins_377 = regs_377_io_out; // @[RegFile.scala 97:16:@57881.4]
  assign rport_io_ins_378 = regs_378_io_out; // @[RegFile.scala 97:16:@57882.4]
  assign rport_io_ins_379 = regs_379_io_out; // @[RegFile.scala 97:16:@57883.4]
  assign rport_io_ins_380 = regs_380_io_out; // @[RegFile.scala 97:16:@57884.4]
  assign rport_io_ins_381 = regs_381_io_out; // @[RegFile.scala 97:16:@57885.4]
  assign rport_io_ins_382 = regs_382_io_out; // @[RegFile.scala 97:16:@57886.4]
  assign rport_io_ins_383 = regs_383_io_out; // @[RegFile.scala 97:16:@57887.4]
  assign rport_io_ins_384 = regs_384_io_out; // @[RegFile.scala 97:16:@57888.4]
  assign rport_io_ins_385 = regs_385_io_out; // @[RegFile.scala 97:16:@57889.4]
  assign rport_io_ins_386 = regs_386_io_out; // @[RegFile.scala 97:16:@57890.4]
  assign rport_io_ins_387 = regs_387_io_out; // @[RegFile.scala 97:16:@57891.4]
  assign rport_io_ins_388 = regs_388_io_out; // @[RegFile.scala 97:16:@57892.4]
  assign rport_io_ins_389 = regs_389_io_out; // @[RegFile.scala 97:16:@57893.4]
  assign rport_io_ins_390 = regs_390_io_out; // @[RegFile.scala 97:16:@57894.4]
  assign rport_io_ins_391 = regs_391_io_out; // @[RegFile.scala 97:16:@57895.4]
  assign rport_io_ins_392 = regs_392_io_out; // @[RegFile.scala 97:16:@57896.4]
  assign rport_io_ins_393 = regs_393_io_out; // @[RegFile.scala 97:16:@57897.4]
  assign rport_io_ins_394 = regs_394_io_out; // @[RegFile.scala 97:16:@57898.4]
  assign rport_io_ins_395 = regs_395_io_out; // @[RegFile.scala 97:16:@57899.4]
  assign rport_io_ins_396 = regs_396_io_out; // @[RegFile.scala 97:16:@57900.4]
  assign rport_io_ins_397 = regs_397_io_out; // @[RegFile.scala 97:16:@57901.4]
  assign rport_io_ins_398 = regs_398_io_out; // @[RegFile.scala 97:16:@57902.4]
  assign rport_io_ins_399 = regs_399_io_out; // @[RegFile.scala 97:16:@57903.4]
  assign rport_io_ins_400 = regs_400_io_out; // @[RegFile.scala 97:16:@57904.4]
  assign rport_io_ins_401 = regs_401_io_out; // @[RegFile.scala 97:16:@57905.4]
  assign rport_io_ins_402 = regs_402_io_out; // @[RegFile.scala 97:16:@57906.4]
  assign rport_io_ins_403 = regs_403_io_out; // @[RegFile.scala 97:16:@57907.4]
  assign rport_io_ins_404 = regs_404_io_out; // @[RegFile.scala 97:16:@57908.4]
  assign rport_io_ins_405 = regs_405_io_out; // @[RegFile.scala 97:16:@57909.4]
  assign rport_io_ins_406 = regs_406_io_out; // @[RegFile.scala 97:16:@57910.4]
  assign rport_io_ins_407 = regs_407_io_out; // @[RegFile.scala 97:16:@57911.4]
  assign rport_io_ins_408 = regs_408_io_out; // @[RegFile.scala 97:16:@57912.4]
  assign rport_io_ins_409 = regs_409_io_out; // @[RegFile.scala 97:16:@57913.4]
  assign rport_io_ins_410 = regs_410_io_out; // @[RegFile.scala 97:16:@57914.4]
  assign rport_io_ins_411 = regs_411_io_out; // @[RegFile.scala 97:16:@57915.4]
  assign rport_io_ins_412 = regs_412_io_out; // @[RegFile.scala 97:16:@57916.4]
  assign rport_io_ins_413 = regs_413_io_out; // @[RegFile.scala 97:16:@57917.4]
  assign rport_io_ins_414 = regs_414_io_out; // @[RegFile.scala 97:16:@57918.4]
  assign rport_io_ins_415 = regs_415_io_out; // @[RegFile.scala 97:16:@57919.4]
  assign rport_io_ins_416 = regs_416_io_out; // @[RegFile.scala 97:16:@57920.4]
  assign rport_io_ins_417 = regs_417_io_out; // @[RegFile.scala 97:16:@57921.4]
  assign rport_io_ins_418 = regs_418_io_out; // @[RegFile.scala 97:16:@57922.4]
  assign rport_io_ins_419 = regs_419_io_out; // @[RegFile.scala 97:16:@57923.4]
  assign rport_io_ins_420 = regs_420_io_out; // @[RegFile.scala 97:16:@57924.4]
  assign rport_io_ins_421 = regs_421_io_out; // @[RegFile.scala 97:16:@57925.4]
  assign rport_io_ins_422 = regs_422_io_out; // @[RegFile.scala 97:16:@57926.4]
  assign rport_io_ins_423 = regs_423_io_out; // @[RegFile.scala 97:16:@57927.4]
  assign rport_io_ins_424 = regs_424_io_out; // @[RegFile.scala 97:16:@57928.4]
  assign rport_io_ins_425 = regs_425_io_out; // @[RegFile.scala 97:16:@57929.4]
  assign rport_io_ins_426 = regs_426_io_out; // @[RegFile.scala 97:16:@57930.4]
  assign rport_io_ins_427 = regs_427_io_out; // @[RegFile.scala 97:16:@57931.4]
  assign rport_io_ins_428 = regs_428_io_out; // @[RegFile.scala 97:16:@57932.4]
  assign rport_io_ins_429 = regs_429_io_out; // @[RegFile.scala 97:16:@57933.4]
  assign rport_io_ins_430 = regs_430_io_out; // @[RegFile.scala 97:16:@57934.4]
  assign rport_io_ins_431 = regs_431_io_out; // @[RegFile.scala 97:16:@57935.4]
  assign rport_io_ins_432 = regs_432_io_out; // @[RegFile.scala 97:16:@57936.4]
  assign rport_io_ins_433 = regs_433_io_out; // @[RegFile.scala 97:16:@57937.4]
  assign rport_io_ins_434 = regs_434_io_out; // @[RegFile.scala 97:16:@57938.4]
  assign rport_io_ins_435 = regs_435_io_out; // @[RegFile.scala 97:16:@57939.4]
  assign rport_io_ins_436 = regs_436_io_out; // @[RegFile.scala 97:16:@57940.4]
  assign rport_io_ins_437 = regs_437_io_out; // @[RegFile.scala 97:16:@57941.4]
  assign rport_io_ins_438 = regs_438_io_out; // @[RegFile.scala 97:16:@57942.4]
  assign rport_io_ins_439 = regs_439_io_out; // @[RegFile.scala 97:16:@57943.4]
  assign rport_io_ins_440 = regs_440_io_out; // @[RegFile.scala 97:16:@57944.4]
  assign rport_io_ins_441 = regs_441_io_out; // @[RegFile.scala 97:16:@57945.4]
  assign rport_io_ins_442 = regs_442_io_out; // @[RegFile.scala 97:16:@57946.4]
  assign rport_io_ins_443 = regs_443_io_out; // @[RegFile.scala 97:16:@57947.4]
  assign rport_io_ins_444 = regs_444_io_out; // @[RegFile.scala 97:16:@57948.4]
  assign rport_io_ins_445 = regs_445_io_out; // @[RegFile.scala 97:16:@57949.4]
  assign rport_io_ins_446 = regs_446_io_out; // @[RegFile.scala 97:16:@57950.4]
  assign rport_io_ins_447 = regs_447_io_out; // @[RegFile.scala 97:16:@57951.4]
  assign rport_io_ins_448 = regs_448_io_out; // @[RegFile.scala 97:16:@57952.4]
  assign rport_io_ins_449 = regs_449_io_out; // @[RegFile.scala 97:16:@57953.4]
  assign rport_io_ins_450 = regs_450_io_out; // @[RegFile.scala 97:16:@57954.4]
  assign rport_io_ins_451 = regs_451_io_out; // @[RegFile.scala 97:16:@57955.4]
  assign rport_io_ins_452 = regs_452_io_out; // @[RegFile.scala 97:16:@57956.4]
  assign rport_io_ins_453 = regs_453_io_out; // @[RegFile.scala 97:16:@57957.4]
  assign rport_io_ins_454 = regs_454_io_out; // @[RegFile.scala 97:16:@57958.4]
  assign rport_io_ins_455 = regs_455_io_out; // @[RegFile.scala 97:16:@57959.4]
  assign rport_io_ins_456 = regs_456_io_out; // @[RegFile.scala 97:16:@57960.4]
  assign rport_io_ins_457 = regs_457_io_out; // @[RegFile.scala 97:16:@57961.4]
  assign rport_io_ins_458 = regs_458_io_out; // @[RegFile.scala 97:16:@57962.4]
  assign rport_io_ins_459 = regs_459_io_out; // @[RegFile.scala 97:16:@57963.4]
  assign rport_io_ins_460 = regs_460_io_out; // @[RegFile.scala 97:16:@57964.4]
  assign rport_io_ins_461 = regs_461_io_out; // @[RegFile.scala 97:16:@57965.4]
  assign rport_io_ins_462 = regs_462_io_out; // @[RegFile.scala 97:16:@57966.4]
  assign rport_io_ins_463 = regs_463_io_out; // @[RegFile.scala 97:16:@57967.4]
  assign rport_io_ins_464 = regs_464_io_out; // @[RegFile.scala 97:16:@57968.4]
  assign rport_io_ins_465 = regs_465_io_out; // @[RegFile.scala 97:16:@57969.4]
  assign rport_io_ins_466 = regs_466_io_out; // @[RegFile.scala 97:16:@57970.4]
  assign rport_io_ins_467 = regs_467_io_out; // @[RegFile.scala 97:16:@57971.4]
  assign rport_io_ins_468 = regs_468_io_out; // @[RegFile.scala 97:16:@57972.4]
  assign rport_io_ins_469 = regs_469_io_out; // @[RegFile.scala 97:16:@57973.4]
  assign rport_io_ins_470 = regs_470_io_out; // @[RegFile.scala 97:16:@57974.4]
  assign rport_io_ins_471 = regs_471_io_out; // @[RegFile.scala 97:16:@57975.4]
  assign rport_io_ins_472 = regs_472_io_out; // @[RegFile.scala 97:16:@57976.4]
  assign rport_io_ins_473 = regs_473_io_out; // @[RegFile.scala 97:16:@57977.4]
  assign rport_io_ins_474 = regs_474_io_out; // @[RegFile.scala 97:16:@57978.4]
  assign rport_io_ins_475 = regs_475_io_out; // @[RegFile.scala 97:16:@57979.4]
  assign rport_io_ins_476 = regs_476_io_out; // @[RegFile.scala 97:16:@57980.4]
  assign rport_io_ins_477 = regs_477_io_out; // @[RegFile.scala 97:16:@57981.4]
  assign rport_io_ins_478 = regs_478_io_out; // @[RegFile.scala 97:16:@57982.4]
  assign rport_io_ins_479 = regs_479_io_out; // @[RegFile.scala 97:16:@57983.4]
  assign rport_io_ins_480 = regs_480_io_out; // @[RegFile.scala 97:16:@57984.4]
  assign rport_io_ins_481 = regs_481_io_out; // @[RegFile.scala 97:16:@57985.4]
  assign rport_io_ins_482 = regs_482_io_out; // @[RegFile.scala 97:16:@57986.4]
  assign rport_io_ins_483 = regs_483_io_out; // @[RegFile.scala 97:16:@57987.4]
  assign rport_io_ins_484 = regs_484_io_out; // @[RegFile.scala 97:16:@57988.4]
  assign rport_io_ins_485 = regs_485_io_out; // @[RegFile.scala 97:16:@57989.4]
  assign rport_io_ins_486 = regs_486_io_out; // @[RegFile.scala 97:16:@57990.4]
  assign rport_io_ins_487 = regs_487_io_out; // @[RegFile.scala 97:16:@57991.4]
  assign rport_io_ins_488 = regs_488_io_out; // @[RegFile.scala 97:16:@57992.4]
  assign rport_io_ins_489 = regs_489_io_out; // @[RegFile.scala 97:16:@57993.4]
  assign rport_io_ins_490 = regs_490_io_out; // @[RegFile.scala 97:16:@57994.4]
  assign rport_io_ins_491 = regs_491_io_out; // @[RegFile.scala 97:16:@57995.4]
  assign rport_io_ins_492 = regs_492_io_out; // @[RegFile.scala 97:16:@57996.4]
  assign rport_io_ins_493 = regs_493_io_out; // @[RegFile.scala 97:16:@57997.4]
  assign rport_io_ins_494 = regs_494_io_out; // @[RegFile.scala 97:16:@57998.4]
  assign rport_io_ins_495 = regs_495_io_out; // @[RegFile.scala 97:16:@57999.4]
  assign rport_io_ins_496 = regs_496_io_out; // @[RegFile.scala 97:16:@58000.4]
  assign rport_io_ins_497 = regs_497_io_out; // @[RegFile.scala 97:16:@58001.4]
  assign rport_io_ins_498 = regs_498_io_out; // @[RegFile.scala 97:16:@58002.4]
  assign rport_io_ins_499 = regs_499_io_out; // @[RegFile.scala 97:16:@58003.4]
  assign rport_io_ins_500 = regs_500_io_out; // @[RegFile.scala 97:16:@58004.4]
  assign rport_io_ins_501 = regs_501_io_out; // @[RegFile.scala 97:16:@58005.4]
  assign rport_io_ins_502 = regs_502_io_out; // @[RegFile.scala 97:16:@58006.4]
  assign rport_io_ins_503 = regs_503_io_out; // @[RegFile.scala 97:16:@58007.4]
  assign rport_io_ins_504 = regs_504_io_out; // @[RegFile.scala 97:16:@58008.4]
  assign rport_io_ins_505 = regs_505_io_out; // @[RegFile.scala 97:16:@58009.4]
  assign rport_io_ins_506 = regs_506_io_out; // @[RegFile.scala 97:16:@58010.4]
  assign rport_io_ins_507 = regs_507_io_out; // @[RegFile.scala 97:16:@58011.4]
  assign rport_io_ins_508 = regs_508_io_out; // @[RegFile.scala 97:16:@58012.4]
  assign rport_io_ins_509 = regs_509_io_out; // @[RegFile.scala 97:16:@58013.4]
  assign rport_io_ins_510 = regs_510_io_out; // @[RegFile.scala 97:16:@58014.4]
  assign rport_io_ins_511 = regs_511_io_out; // @[RegFile.scala 97:16:@58015.4]
  assign rport_io_ins_512 = regs_512_io_out; // @[RegFile.scala 97:16:@58016.4]
  assign rport_io_ins_513 = regs_513_io_out; // @[RegFile.scala 97:16:@58017.4]
  assign rport_io_ins_514 = regs_514_io_out; // @[RegFile.scala 97:16:@58018.4]
  assign rport_io_ins_515 = regs_515_io_out; // @[RegFile.scala 97:16:@58019.4]
  assign rport_io_ins_516 = regs_516_io_out; // @[RegFile.scala 97:16:@58020.4]
  assign rport_io_ins_517 = regs_517_io_out; // @[RegFile.scala 97:16:@58021.4]
  assign rport_io_sel = io_raddr[9:0]; // @[RegFile.scala 106:18:@58022.4]
endmodule
module RetimeWrapper_623( // @[:@58044.2]
  input         clock, // @[:@58045.4]
  input         reset, // @[:@58046.4]
  input  [39:0] io_in, // @[:@58047.4]
  output [39:0] io_out // @[:@58047.4]
);
  wire [39:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@58049.4]
  wire [39:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@58049.4]
  wire [39:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@58049.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@58049.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@58049.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@58049.4]
  RetimeShiftRegister #(.WIDTH(40), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@58049.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@58062.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@58061.4]
  assign sr_init = 40'h0; // @[RetimeShiftRegister.scala 19:16:@58060.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@58059.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@58058.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@58056.4]
endmodule
module FringeFF_518( // @[:@58064.2]
  input         clock, // @[:@58065.4]
  input         reset, // @[:@58066.4]
  input  [39:0] io_in, // @[:@58067.4]
  output [39:0] io_out, // @[:@58067.4]
  input         io_enable // @[:@58067.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@58070.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@58070.4]
  wire [39:0] RetimeWrapper_io_in; // @[package.scala 93:22:@58070.4]
  wire [39:0] RetimeWrapper_io_out; // @[package.scala 93:22:@58070.4]
  wire [39:0] _T_18; // @[package.scala 96:25:@58075.4 package.scala 96:25:@58076.4]
  RetimeWrapper_623 RetimeWrapper ( // @[package.scala 93:22:@58070.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@58075.4 package.scala 96:25:@58076.4]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@58087.4]
  assign RetimeWrapper_clock = clock; // @[:@58071.4]
  assign RetimeWrapper_reset = reset; // @[:@58072.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _T_18; // @[package.scala 94:16:@58073.4]
endmodule
module FringeCounter( // @[:@58089.2]
  input   clock, // @[:@58090.4]
  input   reset, // @[:@58091.4]
  input   io_enable, // @[:@58092.4]
  output  io_done // @[:@58092.4]
);
  wire  reg$_clock; // @[FringeCounter.scala 24:19:@58094.4]
  wire  reg$_reset; // @[FringeCounter.scala 24:19:@58094.4]
  wire [39:0] reg$_io_in; // @[FringeCounter.scala 24:19:@58094.4]
  wire [39:0] reg$_io_out; // @[FringeCounter.scala 24:19:@58094.4]
  wire  reg$_io_enable; // @[FringeCounter.scala 24:19:@58094.4]
  wire [40:0] count; // @[Cat.scala 30:58:@58101.4]
  wire [41:0] _T_25; // @[FringeCounter.scala 31:22:@58102.4]
  wire [40:0] newval; // @[FringeCounter.scala 31:22:@58103.4]
  wire  isMax; // @[FringeCounter.scala 32:22:@58104.4]
  wire [40:0] next; // @[FringeCounter.scala 33:17:@58106.4]
  FringeFF_518 reg$ ( // @[FringeCounter.scala 24:19:@58094.4]
    .clock(reg$_clock),
    .reset(reg$_reset),
    .io_in(reg$_io_in),
    .io_out(reg$_io_out),
    .io_enable(reg$_io_enable)
  );
  assign count = {1'h0,reg$_io_out}; // @[Cat.scala 30:58:@58101.4]
  assign _T_25 = count + 41'h1; // @[FringeCounter.scala 31:22:@58102.4]
  assign newval = count + 41'h1; // @[FringeCounter.scala 31:22:@58103.4]
  assign isMax = newval >= 41'h2cb417800; // @[FringeCounter.scala 32:22:@58104.4]
  assign next = isMax ? count : newval; // @[FringeCounter.scala 33:17:@58106.4]
  assign io_done = io_enable & isMax; // @[FringeCounter.scala 43:11:@58117.4]
  assign reg$_clock = clock; // @[:@58095.4]
  assign reg$_reset = reset; // @[:@58096.4]
  assign reg$_io_in = next[39:0]; // @[FringeCounter.scala 35:15:@58108.6 FringeCounter.scala 37:15:@58111.6]
  assign reg$_io_enable = io_enable; // @[FringeCounter.scala 27:17:@58099.4]
endmodule
module FringeFF_519( // @[:@58151.2]
  input   clock, // @[:@58152.4]
  input   reset, // @[:@58153.4]
  input   io_in, // @[:@58154.4]
  input   io_reset, // @[:@58154.4]
  output  io_out, // @[:@58154.4]
  input   io_enable // @[:@58154.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@58157.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@58157.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@58157.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@58157.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@58157.4]
  wire  _T_18; // @[package.scala 96:25:@58162.4 package.scala 96:25:@58163.4]
  wire  _GEN_0; // @[FringeFF.scala 21:27:@58168.6]
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@58157.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@58162.4 package.scala 96:25:@58163.4]
  assign _GEN_0 = io_reset ? 1'h0 : _T_18; // @[FringeFF.scala 21:27:@58168.6]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@58174.4]
  assign RetimeWrapper_clock = clock; // @[:@58158.4]
  assign RetimeWrapper_reset = reset; // @[:@58159.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@58161.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _GEN_0; // @[package.scala 94:16:@58160.4]
endmodule
module Depulser( // @[:@58176.2]
  input   clock, // @[:@58177.4]
  input   reset, // @[:@58178.4]
  input   io_in, // @[:@58179.4]
  input   io_rst, // @[:@58179.4]
  output  io_out // @[:@58179.4]
);
  wire  r_clock; // @[Depulser.scala 14:17:@58181.4]
  wire  r_reset; // @[Depulser.scala 14:17:@58181.4]
  wire  r_io_in; // @[Depulser.scala 14:17:@58181.4]
  wire  r_io_reset; // @[Depulser.scala 14:17:@58181.4]
  wire  r_io_out; // @[Depulser.scala 14:17:@58181.4]
  wire  r_io_enable; // @[Depulser.scala 14:17:@58181.4]
  FringeFF_519 r ( // @[Depulser.scala 14:17:@58181.4]
    .clock(r_clock),
    .reset(r_reset),
    .io_in(r_io_in),
    .io_reset(r_io_reset),
    .io_out(r_io_out),
    .io_enable(r_io_enable)
  );
  assign io_out = r_io_out; // @[Depulser.scala 19:10:@58190.4]
  assign r_clock = clock; // @[:@58182.4]
  assign r_reset = reset; // @[:@58183.4]
  assign r_io_in = io_rst ? 1'h0 : io_in; // @[Depulser.scala 15:11:@58185.4]
  assign r_io_reset = io_rst; // @[Depulser.scala 18:14:@58189.4]
  assign r_io_enable = io_in | io_rst; // @[Depulser.scala 17:15:@58188.4]
endmodule
module Fringe( // @[:@58192.2]
  input         clock, // @[:@58193.4]
  input         reset, // @[:@58194.4]
  input  [31:0] io_raddr, // @[:@58195.4]
  input         io_wen, // @[:@58195.4]
  input  [31:0] io_waddr, // @[:@58195.4]
  input  [63:0] io_wdata, // @[:@58195.4]
  output [63:0] io_rdata, // @[:@58195.4]
  output        io_enable, // @[:@58195.4]
  input         io_done, // @[:@58195.4]
  output        io_reset, // @[:@58195.4]
  output [63:0] io_argIns_0, // @[:@58195.4]
  input         io_argOuts_0_valid, // @[:@58195.4]
  input  [63:0] io_argOuts_0_bits, // @[:@58195.4]
  input         io_argOuts_1_valid, // @[:@58195.4]
  input  [63:0] io_argOuts_1_bits, // @[:@58195.4]
  input         io_argOuts_2_valid, // @[:@58195.4]
  input  [63:0] io_argOuts_2_bits, // @[:@58195.4]
  input         io_argOuts_3_valid, // @[:@58195.4]
  input  [63:0] io_argOuts_3_bits, // @[:@58195.4]
  input         io_argOuts_4_valid, // @[:@58195.4]
  input  [63:0] io_argOuts_4_bits, // @[:@58195.4]
  input         io_argOuts_5_valid, // @[:@58195.4]
  input  [63:0] io_argOuts_5_bits, // @[:@58195.4]
  input         io_argOuts_6_valid, // @[:@58195.4]
  input  [63:0] io_argOuts_6_bits, // @[:@58195.4]
  input         io_argOuts_7_valid, // @[:@58195.4]
  input  [63:0] io_argOuts_7_bits, // @[:@58195.4]
  input         io_argOuts_8_valid, // @[:@58195.4]
  input  [63:0] io_argOuts_8_bits, // @[:@58195.4]
  input         io_argOuts_9_valid, // @[:@58195.4]
  input  [63:0] io_argOuts_9_bits, // @[:@58195.4]
  input         io_argOuts_10_valid, // @[:@58195.4]
  input  [63:0] io_argOuts_10_bits, // @[:@58195.4]
  input         io_argOuts_11_valid, // @[:@58195.4]
  input  [63:0] io_argOuts_11_bits, // @[:@58195.4]
  input         io_argOuts_12_valid, // @[:@58195.4]
  input  [63:0] io_argOuts_12_bits, // @[:@58195.4]
  input         io_argOuts_13_valid, // @[:@58195.4]
  input  [63:0] io_argOuts_13_bits, // @[:@58195.4]
  input         io_argOuts_14_valid, // @[:@58195.4]
  input  [63:0] io_argOuts_14_bits, // @[:@58195.4]
  input         io_argOuts_15_valid, // @[:@58195.4]
  input  [63:0] io_argOuts_15_bits, // @[:@58195.4]
  output        io_memStreams_loads_0_cmd_ready, // @[:@58195.4]
  input         io_memStreams_loads_0_cmd_valid, // @[:@58195.4]
  input  [63:0] io_memStreams_loads_0_cmd_bits_addr, // @[:@58195.4]
  input  [31:0] io_memStreams_loads_0_cmd_bits_size, // @[:@58195.4]
  input         io_memStreams_loads_0_data_ready, // @[:@58195.4]
  output        io_memStreams_loads_0_data_valid, // @[:@58195.4]
  output [31:0] io_memStreams_loads_0_data_bits_rdata_0, // @[:@58195.4]
  input         io_memStreams_stores_0_cmd_valid, // @[:@58195.4]
  input  [63:0] io_memStreams_stores_0_cmd_bits_addr, // @[:@58195.4]
  input  [31:0] io_memStreams_stores_0_cmd_bits_size, // @[:@58195.4]
  input         io_memStreams_stores_0_data_valid, // @[:@58195.4]
  input  [31:0] io_memStreams_stores_0_data_bits_wdata_0, // @[:@58195.4]
  input  [15:0] io_memStreams_stores_0_data_bits_wstrb, // @[:@58195.4]
  input         io_dram_0_cmd_ready, // @[:@58195.4]
  output        io_dram_0_cmd_valid, // @[:@58195.4]
  output [63:0] io_dram_0_cmd_bits_addr, // @[:@58195.4]
  output [31:0] io_dram_0_cmd_bits_size, // @[:@58195.4]
  output [31:0] io_dram_0_cmd_bits_tag, // @[:@58195.4]
  input         io_dram_0_wdata_ready, // @[:@58195.4]
  output        io_dram_0_wdata_bits_wlast, // @[:@58195.4]
  output        io_dram_0_rresp_ready, // @[:@58195.4]
  input         io_dram_0_rresp_valid, // @[:@58195.4]
  input  [31:0] io_dram_0_rresp_bits_rdata_0, // @[:@58195.4]
  input  [31:0] io_dram_0_rresp_bits_rdata_1, // @[:@58195.4]
  input  [31:0] io_dram_0_rresp_bits_rdata_2, // @[:@58195.4]
  input  [31:0] io_dram_0_rresp_bits_rdata_3, // @[:@58195.4]
  input  [31:0] io_dram_0_rresp_bits_rdata_4, // @[:@58195.4]
  input  [31:0] io_dram_0_rresp_bits_rdata_5, // @[:@58195.4]
  input  [31:0] io_dram_0_rresp_bits_rdata_6, // @[:@58195.4]
  input  [31:0] io_dram_0_rresp_bits_rdata_7, // @[:@58195.4]
  input  [31:0] io_dram_0_rresp_bits_rdata_8, // @[:@58195.4]
  input  [31:0] io_dram_0_rresp_bits_rdata_9, // @[:@58195.4]
  input  [31:0] io_dram_0_rresp_bits_rdata_10, // @[:@58195.4]
  input  [31:0] io_dram_0_rresp_bits_rdata_11, // @[:@58195.4]
  input  [31:0] io_dram_0_rresp_bits_rdata_12, // @[:@58195.4]
  input  [31:0] io_dram_0_rresp_bits_rdata_13, // @[:@58195.4]
  input  [31:0] io_dram_0_rresp_bits_rdata_14, // @[:@58195.4]
  input  [31:0] io_dram_0_rresp_bits_rdata_15, // @[:@58195.4]
  input  [31:0] io_dram_0_rresp_bits_tag, // @[:@58195.4]
  output        io_dram_0_wresp_ready, // @[:@58195.4]
  input         io_dram_0_wresp_valid, // @[:@58195.4]
  input  [31:0] io_dram_0_wresp_bits_tag, // @[:@58195.4]
  input         io_heap_0_req_valid, // @[:@58195.4]
  input         io_heap_0_req_bits_allocDealloc, // @[:@58195.4]
  input  [63:0] io_heap_0_req_bits_sizeAddr, // @[:@58195.4]
  output        io_heap_0_resp_valid, // @[:@58195.4]
  output        io_heap_0_resp_bits_allocDealloc, // @[:@58195.4]
  output [63:0] io_heap_0_resp_bits_sizeAddr // @[:@58195.4]
);
  wire  dramArbs_0_clock; // @[Fringe.scala 91:25:@58261.4]
  wire  dramArbs_0_reset; // @[Fringe.scala 91:25:@58261.4]
  wire  dramArbs_0_io_enable; // @[Fringe.scala 91:25:@58261.4]
  wire  dramArbs_0_io_app_loads_0_cmd_ready; // @[Fringe.scala 91:25:@58261.4]
  wire  dramArbs_0_io_app_loads_0_cmd_valid; // @[Fringe.scala 91:25:@58261.4]
  wire [63:0] dramArbs_0_io_app_loads_0_cmd_bits_addr; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_app_loads_0_cmd_bits_size; // @[Fringe.scala 91:25:@58261.4]
  wire  dramArbs_0_io_app_loads_0_data_ready; // @[Fringe.scala 91:25:@58261.4]
  wire  dramArbs_0_io_app_loads_0_data_valid; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_app_loads_0_data_bits_rdata_0; // @[Fringe.scala 91:25:@58261.4]
  wire  dramArbs_0_io_app_stores_0_cmd_ready; // @[Fringe.scala 91:25:@58261.4]
  wire  dramArbs_0_io_app_stores_0_cmd_valid; // @[Fringe.scala 91:25:@58261.4]
  wire [63:0] dramArbs_0_io_app_stores_0_cmd_bits_addr; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_app_stores_0_cmd_bits_size; // @[Fringe.scala 91:25:@58261.4]
  wire  dramArbs_0_io_app_stores_0_data_ready; // @[Fringe.scala 91:25:@58261.4]
  wire  dramArbs_0_io_app_stores_0_data_valid; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_app_stores_0_data_bits_wdata_0; // @[Fringe.scala 91:25:@58261.4]
  wire [15:0] dramArbs_0_io_app_stores_0_data_bits_wstrb; // @[Fringe.scala 91:25:@58261.4]
  wire  dramArbs_0_io_dram_cmd_ready; // @[Fringe.scala 91:25:@58261.4]
  wire  dramArbs_0_io_dram_cmd_valid; // @[Fringe.scala 91:25:@58261.4]
  wire [63:0] dramArbs_0_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@58261.4]
  wire  dramArbs_0_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@58261.4]
  wire  dramArbs_0_io_dram_wdata_ready; // @[Fringe.scala 91:25:@58261.4]
  wire  dramArbs_0_io_dram_wdata_valid; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@58261.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@58261.4]
  wire  dramArbs_0_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@58261.4]
  wire  dramArbs_0_io_dram_rresp_ready; // @[Fringe.scala 91:25:@58261.4]
  wire  dramArbs_0_io_dram_rresp_valid; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_dram_rresp_bits_rdata_0; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_dram_rresp_bits_rdata_1; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_dram_rresp_bits_rdata_2; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_dram_rresp_bits_rdata_3; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_dram_rresp_bits_rdata_4; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_dram_rresp_bits_rdata_5; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_dram_rresp_bits_rdata_6; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_dram_rresp_bits_rdata_7; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_dram_rresp_bits_rdata_8; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_dram_rresp_bits_rdata_9; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_dram_rresp_bits_rdata_10; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_dram_rresp_bits_rdata_11; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_dram_rresp_bits_rdata_12; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_dram_rresp_bits_rdata_13; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_dram_rresp_bits_rdata_14; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_dram_rresp_bits_rdata_15; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_dram_rresp_bits_tag; // @[Fringe.scala 91:25:@58261.4]
  wire  dramArbs_0_io_dram_wresp_ready; // @[Fringe.scala 91:25:@58261.4]
  wire  dramArbs_0_io_dram_wresp_valid; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_debugSignals_0; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_debugSignals_1; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_debugSignals_2; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_debugSignals_3; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_debugSignals_4; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_debugSignals_5; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_debugSignals_6; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_debugSignals_7; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_debugSignals_8; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_debugSignals_9; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_debugSignals_10; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_debugSignals_11; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_debugSignals_12; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_debugSignals_13; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_debugSignals_14; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_debugSignals_15; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_debugSignals_16; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_debugSignals_17; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_debugSignals_18; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_debugSignals_19; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_debugSignals_20; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_debugSignals_21; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_debugSignals_22; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_debugSignals_23; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_debugSignals_24; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_debugSignals_25; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_debugSignals_26; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_debugSignals_27; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_debugSignals_28; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_debugSignals_29; // @[Fringe.scala 91:25:@58261.4]
  wire [31:0] dramArbs_0_io_debugSignals_40; // @[Fringe.scala 91:25:@58261.4]
  wire  heap_io_accel_0_req_valid; // @[Fringe.scala 107:20:@59254.4]
  wire  heap_io_accel_0_req_bits_allocDealloc; // @[Fringe.scala 107:20:@59254.4]
  wire [63:0] heap_io_accel_0_req_bits_sizeAddr; // @[Fringe.scala 107:20:@59254.4]
  wire  heap_io_accel_0_resp_valid; // @[Fringe.scala 107:20:@59254.4]
  wire  heap_io_accel_0_resp_bits_allocDealloc; // @[Fringe.scala 107:20:@59254.4]
  wire [63:0] heap_io_accel_0_resp_bits_sizeAddr; // @[Fringe.scala 107:20:@59254.4]
  wire  heap_io_host_0_req_valid; // @[Fringe.scala 107:20:@59254.4]
  wire  heap_io_host_0_req_bits_allocDealloc; // @[Fringe.scala 107:20:@59254.4]
  wire [63:0] heap_io_host_0_req_bits_sizeAddr; // @[Fringe.scala 107:20:@59254.4]
  wire  heap_io_host_0_resp_valid; // @[Fringe.scala 107:20:@59254.4]
  wire  heap_io_host_0_resp_bits_allocDealloc; // @[Fringe.scala 107:20:@59254.4]
  wire [63:0] heap_io_host_0_resp_bits_sizeAddr; // @[Fringe.scala 107:20:@59254.4]
  wire  regs_clock; // @[Fringe.scala 116:20:@59263.4]
  wire  regs_reset; // @[Fringe.scala 116:20:@59263.4]
  wire [31:0] regs_io_raddr; // @[Fringe.scala 116:20:@59263.4]
  wire  regs_io_wen; // @[Fringe.scala 116:20:@59263.4]
  wire [31:0] regs_io_waddr; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_wdata; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_rdata; // @[Fringe.scala 116:20:@59263.4]
  wire  regs_io_reset; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argIns_0; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argIns_1; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argIns_2; // @[Fringe.scala 116:20:@59263.4]
  wire  regs_io_argOuts_0_valid; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argOuts_0_bits; // @[Fringe.scala 116:20:@59263.4]
  wire  regs_io_argOuts_1_valid; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argOuts_1_bits; // @[Fringe.scala 116:20:@59263.4]
  wire  regs_io_argOuts_2_valid; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argOuts_2_bits; // @[Fringe.scala 116:20:@59263.4]
  wire  regs_io_argOuts_3_valid; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argOuts_3_bits; // @[Fringe.scala 116:20:@59263.4]
  wire  regs_io_argOuts_4_valid; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argOuts_4_bits; // @[Fringe.scala 116:20:@59263.4]
  wire  regs_io_argOuts_5_valid; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argOuts_5_bits; // @[Fringe.scala 116:20:@59263.4]
  wire  regs_io_argOuts_6_valid; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argOuts_6_bits; // @[Fringe.scala 116:20:@59263.4]
  wire  regs_io_argOuts_7_valid; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argOuts_7_bits; // @[Fringe.scala 116:20:@59263.4]
  wire  regs_io_argOuts_8_valid; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argOuts_8_bits; // @[Fringe.scala 116:20:@59263.4]
  wire  regs_io_argOuts_9_valid; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argOuts_9_bits; // @[Fringe.scala 116:20:@59263.4]
  wire  regs_io_argOuts_10_valid; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argOuts_10_bits; // @[Fringe.scala 116:20:@59263.4]
  wire  regs_io_argOuts_11_valid; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argOuts_11_bits; // @[Fringe.scala 116:20:@59263.4]
  wire  regs_io_argOuts_12_valid; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argOuts_12_bits; // @[Fringe.scala 116:20:@59263.4]
  wire  regs_io_argOuts_13_valid; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argOuts_13_bits; // @[Fringe.scala 116:20:@59263.4]
  wire  regs_io_argOuts_14_valid; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argOuts_14_bits; // @[Fringe.scala 116:20:@59263.4]
  wire  regs_io_argOuts_15_valid; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argOuts_15_bits; // @[Fringe.scala 116:20:@59263.4]
  wire  regs_io_argOuts_16_valid; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argOuts_16_bits; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argOuts_17_bits; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argOuts_18_bits; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argOuts_19_bits; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argOuts_20_bits; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argOuts_21_bits; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argOuts_22_bits; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argOuts_23_bits; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argOuts_24_bits; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argOuts_25_bits; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argOuts_26_bits; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argOuts_27_bits; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argOuts_28_bits; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argOuts_29_bits; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argOuts_30_bits; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argOuts_31_bits; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argOuts_32_bits; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argOuts_33_bits; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argOuts_34_bits; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argOuts_35_bits; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argOuts_36_bits; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argOuts_37_bits; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argOuts_38_bits; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argOuts_39_bits; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argOuts_40_bits; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argOuts_41_bits; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argOuts_42_bits; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argOuts_43_bits; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argOuts_44_bits; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argOuts_45_bits; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argOuts_46_bits; // @[Fringe.scala 116:20:@59263.4]
  wire [63:0] regs_io_argOuts_57_bits; // @[Fringe.scala 116:20:@59263.4]
  wire  timeoutCtr_clock; // @[Fringe.scala 143:26:@61372.4]
  wire  timeoutCtr_reset; // @[Fringe.scala 143:26:@61372.4]
  wire  timeoutCtr_io_enable; // @[Fringe.scala 143:26:@61372.4]
  wire  timeoutCtr_io_done; // @[Fringe.scala 143:26:@61372.4]
  wire  depulser_clock; // @[Fringe.scala 153:24:@61390.4]
  wire  depulser_reset; // @[Fringe.scala 153:24:@61390.4]
  wire  depulser_io_in; // @[Fringe.scala 153:24:@61390.4]
  wire  depulser_io_rst; // @[Fringe.scala 153:24:@61390.4]
  wire  depulser_io_out; // @[Fringe.scala 153:24:@61390.4]
  wire [63:0] _T_916; // @[:@61349.4 :@61350.4]
  wire  curStatus_done; // @[Fringe.scala 133:45:@61351.4]
  wire  curStatus_timeout; // @[Fringe.scala 133:45:@61353.4]
  wire [2:0] curStatus_allocDealloc; // @[Fringe.scala 133:45:@61355.4]
  wire [58:0] curStatus_sizeAddr; // @[Fringe.scala 133:45:@61357.4]
  wire  _T_921; // @[Fringe.scala 134:28:@61359.4]
  wire  _T_925; // @[Fringe.scala 134:42:@61361.4]
  wire  _T_926; // @[Fringe.scala 135:27:@61363.4]
  wire [63:0] _T_936; // @[Fringe.scala 156:22:@61398.4]
  reg  _T_943; // @[package.scala 152:20:@61401.4]
  reg [31:0] _RAND_0;
  wire  _T_944; // @[package.scala 153:13:@61403.4]
  wire  _T_945; // @[package.scala 153:8:@61404.4]
  wire  _T_948; // @[Fringe.scala 160:55:@61408.4]
  wire  status_bits_done; // @[Fringe.scala 160:26:@61409.4]
  wire  _T_951; // @[Fringe.scala 161:58:@61412.4]
  wire  status_bits_timeout; // @[Fringe.scala 161:29:@61413.4]
  wire [1:0] _T_955; // @[Fringe.scala 162:57:@61415.4]
  wire [1:0] _T_957; // @[Fringe.scala 162:34:@61416.4]
  wire [63:0] _T_959; // @[Fringe.scala 163:30:@61418.4]
  wire [1:0] _T_960; // @[Fringe.scala 171:37:@61421.4]
  wire [58:0] status_bits_sizeAddr; // @[Fringe.scala 158:20:@61400.4 Fringe.scala 163:24:@61419.4]
  wire [2:0] status_bits_allocDealloc; // @[Fringe.scala 158:20:@61400.4 Fringe.scala 162:28:@61417.4]
  wire [61:0] _T_961; // @[Fringe.scala 171:37:@61422.4]
  wire  alloc; // @[Fringe.scala 202:38:@62752.4]
  wire  dealloc; // @[Fringe.scala 203:40:@62753.4]
  wire  _T_1465; // @[Fringe.scala 204:37:@62754.4]
  reg  _T_1468; // @[package.scala 152:20:@62755.4]
  reg [31:0] _RAND_1;
  wire  _T_1469; // @[package.scala 153:13:@62757.4]
  DRAMArbiter dramArbs_0 ( // @[Fringe.scala 91:25:@58261.4]
    .clock(dramArbs_0_clock),
    .reset(dramArbs_0_reset),
    .io_enable(dramArbs_0_io_enable),
    .io_app_loads_0_cmd_ready(dramArbs_0_io_app_loads_0_cmd_ready),
    .io_app_loads_0_cmd_valid(dramArbs_0_io_app_loads_0_cmd_valid),
    .io_app_loads_0_cmd_bits_addr(dramArbs_0_io_app_loads_0_cmd_bits_addr),
    .io_app_loads_0_cmd_bits_size(dramArbs_0_io_app_loads_0_cmd_bits_size),
    .io_app_loads_0_data_ready(dramArbs_0_io_app_loads_0_data_ready),
    .io_app_loads_0_data_valid(dramArbs_0_io_app_loads_0_data_valid),
    .io_app_loads_0_data_bits_rdata_0(dramArbs_0_io_app_loads_0_data_bits_rdata_0),
    .io_app_stores_0_cmd_ready(dramArbs_0_io_app_stores_0_cmd_ready),
    .io_app_stores_0_cmd_valid(dramArbs_0_io_app_stores_0_cmd_valid),
    .io_app_stores_0_cmd_bits_addr(dramArbs_0_io_app_stores_0_cmd_bits_addr),
    .io_app_stores_0_cmd_bits_size(dramArbs_0_io_app_stores_0_cmd_bits_size),
    .io_app_stores_0_data_ready(dramArbs_0_io_app_stores_0_data_ready),
    .io_app_stores_0_data_valid(dramArbs_0_io_app_stores_0_data_valid),
    .io_app_stores_0_data_bits_wdata_0(dramArbs_0_io_app_stores_0_data_bits_wdata_0),
    .io_app_stores_0_data_bits_wstrb(dramArbs_0_io_app_stores_0_data_bits_wstrb),
    .io_dram_cmd_ready(dramArbs_0_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_0_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_0_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_0_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_0_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_0_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_0_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_0_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_0_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wstrb_0(dramArbs_0_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wlast(dramArbs_0_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_0_io_dram_rresp_ready),
    .io_dram_rresp_valid(dramArbs_0_io_dram_rresp_valid),
    .io_dram_rresp_bits_rdata_0(dramArbs_0_io_dram_rresp_bits_rdata_0),
    .io_dram_rresp_bits_rdata_1(dramArbs_0_io_dram_rresp_bits_rdata_1),
    .io_dram_rresp_bits_rdata_2(dramArbs_0_io_dram_rresp_bits_rdata_2),
    .io_dram_rresp_bits_rdata_3(dramArbs_0_io_dram_rresp_bits_rdata_3),
    .io_dram_rresp_bits_rdata_4(dramArbs_0_io_dram_rresp_bits_rdata_4),
    .io_dram_rresp_bits_rdata_5(dramArbs_0_io_dram_rresp_bits_rdata_5),
    .io_dram_rresp_bits_rdata_6(dramArbs_0_io_dram_rresp_bits_rdata_6),
    .io_dram_rresp_bits_rdata_7(dramArbs_0_io_dram_rresp_bits_rdata_7),
    .io_dram_rresp_bits_rdata_8(dramArbs_0_io_dram_rresp_bits_rdata_8),
    .io_dram_rresp_bits_rdata_9(dramArbs_0_io_dram_rresp_bits_rdata_9),
    .io_dram_rresp_bits_rdata_10(dramArbs_0_io_dram_rresp_bits_rdata_10),
    .io_dram_rresp_bits_rdata_11(dramArbs_0_io_dram_rresp_bits_rdata_11),
    .io_dram_rresp_bits_rdata_12(dramArbs_0_io_dram_rresp_bits_rdata_12),
    .io_dram_rresp_bits_rdata_13(dramArbs_0_io_dram_rresp_bits_rdata_13),
    .io_dram_rresp_bits_rdata_14(dramArbs_0_io_dram_rresp_bits_rdata_14),
    .io_dram_rresp_bits_rdata_15(dramArbs_0_io_dram_rresp_bits_rdata_15),
    .io_dram_rresp_bits_tag(dramArbs_0_io_dram_rresp_bits_tag),
    .io_dram_wresp_ready(dramArbs_0_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_0_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_0_io_dram_wresp_bits_tag),
    .io_debugSignals_0(dramArbs_0_io_debugSignals_0),
    .io_debugSignals_1(dramArbs_0_io_debugSignals_1),
    .io_debugSignals_2(dramArbs_0_io_debugSignals_2),
    .io_debugSignals_3(dramArbs_0_io_debugSignals_3),
    .io_debugSignals_4(dramArbs_0_io_debugSignals_4),
    .io_debugSignals_5(dramArbs_0_io_debugSignals_5),
    .io_debugSignals_6(dramArbs_0_io_debugSignals_6),
    .io_debugSignals_7(dramArbs_0_io_debugSignals_7),
    .io_debugSignals_8(dramArbs_0_io_debugSignals_8),
    .io_debugSignals_9(dramArbs_0_io_debugSignals_9),
    .io_debugSignals_10(dramArbs_0_io_debugSignals_10),
    .io_debugSignals_11(dramArbs_0_io_debugSignals_11),
    .io_debugSignals_12(dramArbs_0_io_debugSignals_12),
    .io_debugSignals_13(dramArbs_0_io_debugSignals_13),
    .io_debugSignals_14(dramArbs_0_io_debugSignals_14),
    .io_debugSignals_15(dramArbs_0_io_debugSignals_15),
    .io_debugSignals_16(dramArbs_0_io_debugSignals_16),
    .io_debugSignals_17(dramArbs_0_io_debugSignals_17),
    .io_debugSignals_18(dramArbs_0_io_debugSignals_18),
    .io_debugSignals_19(dramArbs_0_io_debugSignals_19),
    .io_debugSignals_20(dramArbs_0_io_debugSignals_20),
    .io_debugSignals_21(dramArbs_0_io_debugSignals_21),
    .io_debugSignals_22(dramArbs_0_io_debugSignals_22),
    .io_debugSignals_23(dramArbs_0_io_debugSignals_23),
    .io_debugSignals_24(dramArbs_0_io_debugSignals_24),
    .io_debugSignals_25(dramArbs_0_io_debugSignals_25),
    .io_debugSignals_26(dramArbs_0_io_debugSignals_26),
    .io_debugSignals_27(dramArbs_0_io_debugSignals_27),
    .io_debugSignals_28(dramArbs_0_io_debugSignals_28),
    .io_debugSignals_29(dramArbs_0_io_debugSignals_29),
    .io_debugSignals_40(dramArbs_0_io_debugSignals_40)
  );
  DRAMHeap heap ( // @[Fringe.scala 107:20:@59254.4]
    .io_accel_0_req_valid(heap_io_accel_0_req_valid),
    .io_accel_0_req_bits_allocDealloc(heap_io_accel_0_req_bits_allocDealloc),
    .io_accel_0_req_bits_sizeAddr(heap_io_accel_0_req_bits_sizeAddr),
    .io_accel_0_resp_valid(heap_io_accel_0_resp_valid),
    .io_accel_0_resp_bits_allocDealloc(heap_io_accel_0_resp_bits_allocDealloc),
    .io_accel_0_resp_bits_sizeAddr(heap_io_accel_0_resp_bits_sizeAddr),
    .io_host_0_req_valid(heap_io_host_0_req_valid),
    .io_host_0_req_bits_allocDealloc(heap_io_host_0_req_bits_allocDealloc),
    .io_host_0_req_bits_sizeAddr(heap_io_host_0_req_bits_sizeAddr),
    .io_host_0_resp_valid(heap_io_host_0_resp_valid),
    .io_host_0_resp_bits_allocDealloc(heap_io_host_0_resp_bits_allocDealloc),
    .io_host_0_resp_bits_sizeAddr(heap_io_host_0_resp_bits_sizeAddr)
  );
  RegFile regs ( // @[Fringe.scala 116:20:@59263.4]
    .clock(regs_clock),
    .reset(regs_reset),
    .io_raddr(regs_io_raddr),
    .io_wen(regs_io_wen),
    .io_waddr(regs_io_waddr),
    .io_wdata(regs_io_wdata),
    .io_rdata(regs_io_rdata),
    .io_reset(regs_io_reset),
    .io_argIns_0(regs_io_argIns_0),
    .io_argIns_1(regs_io_argIns_1),
    .io_argIns_2(regs_io_argIns_2),
    .io_argOuts_0_valid(regs_io_argOuts_0_valid),
    .io_argOuts_0_bits(regs_io_argOuts_0_bits),
    .io_argOuts_1_valid(regs_io_argOuts_1_valid),
    .io_argOuts_1_bits(regs_io_argOuts_1_bits),
    .io_argOuts_2_valid(regs_io_argOuts_2_valid),
    .io_argOuts_2_bits(regs_io_argOuts_2_bits),
    .io_argOuts_3_valid(regs_io_argOuts_3_valid),
    .io_argOuts_3_bits(regs_io_argOuts_3_bits),
    .io_argOuts_4_valid(regs_io_argOuts_4_valid),
    .io_argOuts_4_bits(regs_io_argOuts_4_bits),
    .io_argOuts_5_valid(regs_io_argOuts_5_valid),
    .io_argOuts_5_bits(regs_io_argOuts_5_bits),
    .io_argOuts_6_valid(regs_io_argOuts_6_valid),
    .io_argOuts_6_bits(regs_io_argOuts_6_bits),
    .io_argOuts_7_valid(regs_io_argOuts_7_valid),
    .io_argOuts_7_bits(regs_io_argOuts_7_bits),
    .io_argOuts_8_valid(regs_io_argOuts_8_valid),
    .io_argOuts_8_bits(regs_io_argOuts_8_bits),
    .io_argOuts_9_valid(regs_io_argOuts_9_valid),
    .io_argOuts_9_bits(regs_io_argOuts_9_bits),
    .io_argOuts_10_valid(regs_io_argOuts_10_valid),
    .io_argOuts_10_bits(regs_io_argOuts_10_bits),
    .io_argOuts_11_valid(regs_io_argOuts_11_valid),
    .io_argOuts_11_bits(regs_io_argOuts_11_bits),
    .io_argOuts_12_valid(regs_io_argOuts_12_valid),
    .io_argOuts_12_bits(regs_io_argOuts_12_bits),
    .io_argOuts_13_valid(regs_io_argOuts_13_valid),
    .io_argOuts_13_bits(regs_io_argOuts_13_bits),
    .io_argOuts_14_valid(regs_io_argOuts_14_valid),
    .io_argOuts_14_bits(regs_io_argOuts_14_bits),
    .io_argOuts_15_valid(regs_io_argOuts_15_valid),
    .io_argOuts_15_bits(regs_io_argOuts_15_bits),
    .io_argOuts_16_valid(regs_io_argOuts_16_valid),
    .io_argOuts_16_bits(regs_io_argOuts_16_bits),
    .io_argOuts_17_bits(regs_io_argOuts_17_bits),
    .io_argOuts_18_bits(regs_io_argOuts_18_bits),
    .io_argOuts_19_bits(regs_io_argOuts_19_bits),
    .io_argOuts_20_bits(regs_io_argOuts_20_bits),
    .io_argOuts_21_bits(regs_io_argOuts_21_bits),
    .io_argOuts_22_bits(regs_io_argOuts_22_bits),
    .io_argOuts_23_bits(regs_io_argOuts_23_bits),
    .io_argOuts_24_bits(regs_io_argOuts_24_bits),
    .io_argOuts_25_bits(regs_io_argOuts_25_bits),
    .io_argOuts_26_bits(regs_io_argOuts_26_bits),
    .io_argOuts_27_bits(regs_io_argOuts_27_bits),
    .io_argOuts_28_bits(regs_io_argOuts_28_bits),
    .io_argOuts_29_bits(regs_io_argOuts_29_bits),
    .io_argOuts_30_bits(regs_io_argOuts_30_bits),
    .io_argOuts_31_bits(regs_io_argOuts_31_bits),
    .io_argOuts_32_bits(regs_io_argOuts_32_bits),
    .io_argOuts_33_bits(regs_io_argOuts_33_bits),
    .io_argOuts_34_bits(regs_io_argOuts_34_bits),
    .io_argOuts_35_bits(regs_io_argOuts_35_bits),
    .io_argOuts_36_bits(regs_io_argOuts_36_bits),
    .io_argOuts_37_bits(regs_io_argOuts_37_bits),
    .io_argOuts_38_bits(regs_io_argOuts_38_bits),
    .io_argOuts_39_bits(regs_io_argOuts_39_bits),
    .io_argOuts_40_bits(regs_io_argOuts_40_bits),
    .io_argOuts_41_bits(regs_io_argOuts_41_bits),
    .io_argOuts_42_bits(regs_io_argOuts_42_bits),
    .io_argOuts_43_bits(regs_io_argOuts_43_bits),
    .io_argOuts_44_bits(regs_io_argOuts_44_bits),
    .io_argOuts_45_bits(regs_io_argOuts_45_bits),
    .io_argOuts_46_bits(regs_io_argOuts_46_bits),
    .io_argOuts_57_bits(regs_io_argOuts_57_bits)
  );
  FringeCounter timeoutCtr ( // @[Fringe.scala 143:26:@61372.4]
    .clock(timeoutCtr_clock),
    .reset(timeoutCtr_reset),
    .io_enable(timeoutCtr_io_enable),
    .io_done(timeoutCtr_io_done)
  );
  Depulser depulser ( // @[Fringe.scala 153:24:@61390.4]
    .clock(depulser_clock),
    .reset(depulser_reset),
    .io_in(depulser_io_in),
    .io_rst(depulser_io_rst),
    .io_out(depulser_io_out)
  );
  assign _T_916 = regs_io_argIns_1; // @[:@61349.4 :@61350.4]
  assign curStatus_done = _T_916[0]; // @[Fringe.scala 133:45:@61351.4]
  assign curStatus_timeout = _T_916[1]; // @[Fringe.scala 133:45:@61353.4]
  assign curStatus_allocDealloc = _T_916[4:2]; // @[Fringe.scala 133:45:@61355.4]
  assign curStatus_sizeAddr = _T_916[63:5]; // @[Fringe.scala 133:45:@61357.4]
  assign _T_921 = regs_io_argIns_0[0]; // @[Fringe.scala 134:28:@61359.4]
  assign _T_925 = curStatus_done == 1'h0; // @[Fringe.scala 134:42:@61361.4]
  assign _T_926 = regs_io_argIns_0[1]; // @[Fringe.scala 135:27:@61363.4]
  assign _T_936 = ~ regs_io_argIns_0; // @[Fringe.scala 156:22:@61398.4]
  assign _T_944 = _T_943 ^ heap_io_host_0_req_valid; // @[package.scala 153:13:@61403.4]
  assign _T_945 = heap_io_host_0_req_valid & _T_944; // @[package.scala 153:8:@61404.4]
  assign _T_948 = _T_921 & depulser_io_out; // @[Fringe.scala 160:55:@61408.4]
  assign status_bits_done = depulser_io_out ? _T_948 : curStatus_done; // @[Fringe.scala 160:26:@61409.4]
  assign _T_951 = _T_921 & timeoutCtr_io_done; // @[Fringe.scala 161:58:@61412.4]
  assign status_bits_timeout = depulser_io_out ? _T_951 : curStatus_timeout; // @[Fringe.scala 161:29:@61413.4]
  assign _T_955 = heap_io_host_0_req_bits_allocDealloc ? 2'h1 : 2'h2; // @[Fringe.scala 162:57:@61415.4]
  assign _T_957 = heap_io_host_0_req_valid ? _T_955 : 2'h0; // @[Fringe.scala 162:34:@61416.4]
  assign _T_959 = heap_io_host_0_req_valid ? heap_io_host_0_req_bits_sizeAddr : 64'h0; // @[Fringe.scala 163:30:@61418.4]
  assign _T_960 = {status_bits_timeout,status_bits_done}; // @[Fringe.scala 171:37:@61421.4]
  assign status_bits_sizeAddr = _T_959[58:0]; // @[Fringe.scala 158:20:@61400.4 Fringe.scala 163:24:@61419.4]
  assign status_bits_allocDealloc = {{1'd0}, _T_957}; // @[Fringe.scala 158:20:@61400.4 Fringe.scala 162:28:@61417.4]
  assign _T_961 = {status_bits_sizeAddr,status_bits_allocDealloc}; // @[Fringe.scala 171:37:@61422.4]
  assign alloc = curStatus_allocDealloc == 3'h3; // @[Fringe.scala 202:38:@62752.4]
  assign dealloc = curStatus_allocDealloc == 3'h4; // @[Fringe.scala 203:40:@62753.4]
  assign _T_1465 = alloc | dealloc; // @[Fringe.scala 204:37:@62754.4]
  assign _T_1469 = _T_1468 ^ _T_1465; // @[package.scala 153:13:@62757.4]
  assign io_rdata = regs_io_rdata; // @[Fringe.scala 125:14:@61347.4]
  assign io_enable = _T_921 & _T_925; // @[Fringe.scala 136:13:@61367.4]
  assign io_reset = _T_926 | reset; // @[Fringe.scala 137:12:@61368.4]
  assign io_argIns_0 = regs_io_argIns_2; // @[Fringe.scala 151:51:@61389.4]
  assign io_memStreams_loads_0_cmd_ready = dramArbs_0_io_app_loads_0_cmd_ready; // @[Fringe.scala 100:70:@59154.4]
  assign io_memStreams_loads_0_data_valid = dramArbs_0_io_app_loads_0_data_valid; // @[Fringe.scala 100:70:@59149.4]
  assign io_memStreams_loads_0_data_bits_rdata_0 = dramArbs_0_io_app_loads_0_data_bits_rdata_0; // @[Fringe.scala 100:70:@59148.4]
  assign io_dram_0_cmd_valid = dramArbs_0_io_dram_cmd_valid; // @[Fringe.scala 195:72:@62586.4]
  assign io_dram_0_cmd_bits_addr = dramArbs_0_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@62585.4]
  assign io_dram_0_cmd_bits_size = dramArbs_0_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@62584.4]
  assign io_dram_0_cmd_bits_tag = dramArbs_0_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@62581.4]
  assign io_dram_0_wdata_bits_wlast = dramArbs_0_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@62498.4]
  assign io_dram_0_rresp_ready = dramArbs_0_io_dram_rresp_ready; // @[Fringe.scala 195:72:@62497.4]
  assign io_dram_0_wresp_ready = dramArbs_0_io_dram_wresp_ready; // @[Fringe.scala 195:72:@62478.4]
  assign io_heap_0_resp_valid = heap_io_accel_0_resp_valid; // @[Fringe.scala 108:17:@59259.4]
  assign io_heap_0_resp_bits_allocDealloc = heap_io_accel_0_resp_bits_allocDealloc; // @[Fringe.scala 108:17:@59258.4]
  assign io_heap_0_resp_bits_sizeAddr = heap_io_accel_0_resp_bits_sizeAddr; // @[Fringe.scala 108:17:@59257.4]
  assign dramArbs_0_clock = clock; // @[:@58262.4]
  assign dramArbs_0_reset = _T_926 | reset; // @[:@58263.4 Fringe.scala 187:30:@62474.4]
  assign dramArbs_0_io_enable = _T_921 & _T_925; // @[Fringe.scala 192:36:@62475.4]
  assign dramArbs_0_io_app_loads_0_cmd_valid = io_memStreams_loads_0_cmd_valid; // @[Fringe.scala 100:70:@59153.4]
  assign dramArbs_0_io_app_loads_0_cmd_bits_addr = io_memStreams_loads_0_cmd_bits_addr; // @[Fringe.scala 100:70:@59152.4]
  assign dramArbs_0_io_app_loads_0_cmd_bits_size = io_memStreams_loads_0_cmd_bits_size; // @[Fringe.scala 100:70:@59151.4]
  assign dramArbs_0_io_app_loads_0_data_ready = io_memStreams_loads_0_data_ready; // @[Fringe.scala 100:70:@59150.4]
  assign dramArbs_0_io_app_stores_0_cmd_valid = io_memStreams_stores_0_cmd_valid; // @[Fringe.scala 101:72:@59179.4]
  assign dramArbs_0_io_app_stores_0_cmd_bits_addr = io_memStreams_stores_0_cmd_bits_addr; // @[Fringe.scala 101:72:@59178.4]
  assign dramArbs_0_io_app_stores_0_cmd_bits_size = io_memStreams_stores_0_cmd_bits_size; // @[Fringe.scala 101:72:@59177.4]
  assign dramArbs_0_io_app_stores_0_data_valid = io_memStreams_stores_0_data_valid; // @[Fringe.scala 101:72:@59175.4]
  assign dramArbs_0_io_app_stores_0_data_bits_wdata_0 = io_memStreams_stores_0_data_bits_wdata_0; // @[Fringe.scala 101:72:@59159.4]
  assign dramArbs_0_io_app_stores_0_data_bits_wstrb = io_memStreams_stores_0_data_bits_wstrb; // @[Fringe.scala 101:72:@59158.4]
  assign dramArbs_0_io_dram_cmd_ready = io_dram_0_cmd_ready; // @[Fringe.scala 195:72:@62587.4]
  assign dramArbs_0_io_dram_wdata_ready = io_dram_0_wdata_ready; // @[Fringe.scala 195:72:@62580.4]
  assign dramArbs_0_io_dram_rresp_valid = io_dram_0_rresp_valid; // @[Fringe.scala 195:72:@62496.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_0 = io_dram_0_rresp_bits_rdata_0; // @[Fringe.scala 195:72:@62480.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_1 = io_dram_0_rresp_bits_rdata_1; // @[Fringe.scala 195:72:@62481.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_2 = io_dram_0_rresp_bits_rdata_2; // @[Fringe.scala 195:72:@62482.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_3 = io_dram_0_rresp_bits_rdata_3; // @[Fringe.scala 195:72:@62483.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_4 = io_dram_0_rresp_bits_rdata_4; // @[Fringe.scala 195:72:@62484.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_5 = io_dram_0_rresp_bits_rdata_5; // @[Fringe.scala 195:72:@62485.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_6 = io_dram_0_rresp_bits_rdata_6; // @[Fringe.scala 195:72:@62486.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_7 = io_dram_0_rresp_bits_rdata_7; // @[Fringe.scala 195:72:@62487.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_8 = io_dram_0_rresp_bits_rdata_8; // @[Fringe.scala 195:72:@62488.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_9 = io_dram_0_rresp_bits_rdata_9; // @[Fringe.scala 195:72:@62489.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_10 = io_dram_0_rresp_bits_rdata_10; // @[Fringe.scala 195:72:@62490.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_11 = io_dram_0_rresp_bits_rdata_11; // @[Fringe.scala 195:72:@62491.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_12 = io_dram_0_rresp_bits_rdata_12; // @[Fringe.scala 195:72:@62492.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_13 = io_dram_0_rresp_bits_rdata_13; // @[Fringe.scala 195:72:@62493.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_14 = io_dram_0_rresp_bits_rdata_14; // @[Fringe.scala 195:72:@62494.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_15 = io_dram_0_rresp_bits_rdata_15; // @[Fringe.scala 195:72:@62495.4]
  assign dramArbs_0_io_dram_rresp_bits_tag = io_dram_0_rresp_bits_tag; // @[Fringe.scala 195:72:@62479.4]
  assign dramArbs_0_io_dram_wresp_valid = io_dram_0_wresp_valid; // @[Fringe.scala 195:72:@62477.4]
  assign dramArbs_0_io_dram_wresp_bits_tag = io_dram_0_wresp_bits_tag; // @[Fringe.scala 195:72:@62476.4]
  assign heap_io_accel_0_req_valid = io_heap_0_req_valid; // @[Fringe.scala 108:17:@59262.4]
  assign heap_io_accel_0_req_bits_allocDealloc = io_heap_0_req_bits_allocDealloc; // @[Fringe.scala 108:17:@59261.4]
  assign heap_io_accel_0_req_bits_sizeAddr = io_heap_0_req_bits_sizeAddr; // @[Fringe.scala 108:17:@59260.4]
  assign heap_io_host_0_resp_valid = _T_1465 & _T_1469; // @[Fringe.scala 204:22:@62759.4]
  assign heap_io_host_0_resp_bits_allocDealloc = curStatus_allocDealloc == 3'h3; // @[Fringe.scala 205:34:@62760.4]
  assign heap_io_host_0_resp_bits_sizeAddr = {{5'd0}, curStatus_sizeAddr}; // @[Fringe.scala 206:30:@62761.4]
  assign regs_clock = clock; // @[:@59264.4]
  assign regs_reset = reset; // @[:@59265.4 Fringe.scala 139:14:@61371.4]
  assign regs_io_raddr = io_raddr; // @[Fringe.scala 118:17:@61343.4]
  assign regs_io_wen = io_wen; // @[Fringe.scala 120:15:@61345.4]
  assign regs_io_waddr = io_waddr; // @[Fringe.scala 119:17:@61344.4]
  assign regs_io_wdata = io_wdata; // @[Fringe.scala 121:17:@61346.4]
  assign regs_io_reset = _T_926 | reset; // @[Fringe.scala 138:17:@61369.4]
  assign regs_io_argOuts_0_valid = depulser_io_out | _T_945; // @[Fringe.scala 170:23:@61420.4]
  assign regs_io_argOuts_0_bits = {_T_961,_T_960}; // @[Fringe.scala 171:22:@61424.4]
  assign regs_io_argOuts_1_valid = io_argOuts_0_valid; // @[Fringe.scala 176:23:@61427.4]
  assign regs_io_argOuts_1_bits = io_argOuts_0_bits; // @[Fringe.scala 175:22:@61426.4]
  assign regs_io_argOuts_2_valid = io_argOuts_1_valid; // @[Fringe.scala 176:23:@61430.4]
  assign regs_io_argOuts_2_bits = io_argOuts_1_bits; // @[Fringe.scala 175:22:@61429.4]
  assign regs_io_argOuts_3_valid = io_argOuts_2_valid; // @[Fringe.scala 176:23:@61433.4]
  assign regs_io_argOuts_3_bits = io_argOuts_2_bits; // @[Fringe.scala 175:22:@61432.4]
  assign regs_io_argOuts_4_valid = io_argOuts_3_valid; // @[Fringe.scala 176:23:@61436.4]
  assign regs_io_argOuts_4_bits = io_argOuts_3_bits; // @[Fringe.scala 175:22:@61435.4]
  assign regs_io_argOuts_5_valid = io_argOuts_4_valid; // @[Fringe.scala 176:23:@61439.4]
  assign regs_io_argOuts_5_bits = io_argOuts_4_bits; // @[Fringe.scala 175:22:@61438.4]
  assign regs_io_argOuts_6_valid = io_argOuts_5_valid; // @[Fringe.scala 176:23:@61442.4]
  assign regs_io_argOuts_6_bits = io_argOuts_5_bits; // @[Fringe.scala 175:22:@61441.4]
  assign regs_io_argOuts_7_valid = io_argOuts_6_valid; // @[Fringe.scala 176:23:@61445.4]
  assign regs_io_argOuts_7_bits = io_argOuts_6_bits; // @[Fringe.scala 175:22:@61444.4]
  assign regs_io_argOuts_8_valid = io_argOuts_7_valid; // @[Fringe.scala 176:23:@61448.4]
  assign regs_io_argOuts_8_bits = io_argOuts_7_bits; // @[Fringe.scala 175:22:@61447.4]
  assign regs_io_argOuts_9_valid = io_argOuts_8_valid; // @[Fringe.scala 176:23:@61451.4]
  assign regs_io_argOuts_9_bits = io_argOuts_8_bits; // @[Fringe.scala 175:22:@61450.4]
  assign regs_io_argOuts_10_valid = io_argOuts_9_valid; // @[Fringe.scala 176:23:@61454.4]
  assign regs_io_argOuts_10_bits = io_argOuts_9_bits; // @[Fringe.scala 175:22:@61453.4]
  assign regs_io_argOuts_11_valid = io_argOuts_10_valid; // @[Fringe.scala 176:23:@61457.4]
  assign regs_io_argOuts_11_bits = io_argOuts_10_bits; // @[Fringe.scala 175:22:@61456.4]
  assign regs_io_argOuts_12_valid = io_argOuts_11_valid; // @[Fringe.scala 176:23:@61460.4]
  assign regs_io_argOuts_12_bits = io_argOuts_11_bits; // @[Fringe.scala 175:22:@61459.4]
  assign regs_io_argOuts_13_valid = io_argOuts_12_valid; // @[Fringe.scala 176:23:@61463.4]
  assign regs_io_argOuts_13_bits = io_argOuts_12_bits; // @[Fringe.scala 175:22:@61462.4]
  assign regs_io_argOuts_14_valid = io_argOuts_13_valid; // @[Fringe.scala 176:23:@61466.4]
  assign regs_io_argOuts_14_bits = io_argOuts_13_bits; // @[Fringe.scala 175:22:@61465.4]
  assign regs_io_argOuts_15_valid = io_argOuts_14_valid; // @[Fringe.scala 176:23:@61469.4]
  assign regs_io_argOuts_15_bits = io_argOuts_14_bits; // @[Fringe.scala 175:22:@61468.4]
  assign regs_io_argOuts_16_valid = io_argOuts_15_valid; // @[Fringe.scala 176:23:@61472.4]
  assign regs_io_argOuts_16_bits = io_argOuts_15_bits; // @[Fringe.scala 175:22:@61471.4]
  assign regs_io_argOuts_17_bits = {{32'd0}, dramArbs_0_io_debugSignals_0}; // @[Fringe.scala 179:22:@61473.4]
  assign regs_io_argOuts_18_bits = {{32'd0}, dramArbs_0_io_debugSignals_1}; // @[Fringe.scala 179:22:@61475.4]
  assign regs_io_argOuts_19_bits = {{32'd0}, dramArbs_0_io_debugSignals_2}; // @[Fringe.scala 179:22:@61477.4]
  assign regs_io_argOuts_20_bits = {{32'd0}, dramArbs_0_io_debugSignals_3}; // @[Fringe.scala 179:22:@61479.4]
  assign regs_io_argOuts_21_bits = {{32'd0}, dramArbs_0_io_debugSignals_4}; // @[Fringe.scala 179:22:@61481.4]
  assign regs_io_argOuts_22_bits = {{32'd0}, dramArbs_0_io_debugSignals_5}; // @[Fringe.scala 179:22:@61483.4]
  assign regs_io_argOuts_23_bits = {{32'd0}, dramArbs_0_io_debugSignals_6}; // @[Fringe.scala 179:22:@61485.4]
  assign regs_io_argOuts_24_bits = {{32'd0}, dramArbs_0_io_debugSignals_7}; // @[Fringe.scala 179:22:@61487.4]
  assign regs_io_argOuts_25_bits = {{32'd0}, dramArbs_0_io_debugSignals_8}; // @[Fringe.scala 179:22:@61489.4]
  assign regs_io_argOuts_26_bits = {{32'd0}, dramArbs_0_io_debugSignals_9}; // @[Fringe.scala 179:22:@61491.4]
  assign regs_io_argOuts_27_bits = {{32'd0}, dramArbs_0_io_debugSignals_10}; // @[Fringe.scala 179:22:@61493.4]
  assign regs_io_argOuts_28_bits = {{32'd0}, dramArbs_0_io_debugSignals_11}; // @[Fringe.scala 179:22:@61495.4]
  assign regs_io_argOuts_29_bits = {{32'd0}, dramArbs_0_io_debugSignals_12}; // @[Fringe.scala 179:22:@61497.4]
  assign regs_io_argOuts_30_bits = {{32'd0}, dramArbs_0_io_debugSignals_13}; // @[Fringe.scala 179:22:@61499.4]
  assign regs_io_argOuts_31_bits = {{32'd0}, dramArbs_0_io_debugSignals_14}; // @[Fringe.scala 179:22:@61501.4]
  assign regs_io_argOuts_32_bits = {{32'd0}, dramArbs_0_io_debugSignals_15}; // @[Fringe.scala 179:22:@61503.4]
  assign regs_io_argOuts_33_bits = {{32'd0}, dramArbs_0_io_debugSignals_16}; // @[Fringe.scala 179:22:@61505.4]
  assign regs_io_argOuts_34_bits = {{32'd0}, dramArbs_0_io_debugSignals_17}; // @[Fringe.scala 179:22:@61507.4]
  assign regs_io_argOuts_35_bits = {{32'd0}, dramArbs_0_io_debugSignals_18}; // @[Fringe.scala 179:22:@61509.4]
  assign regs_io_argOuts_36_bits = {{32'd0}, dramArbs_0_io_debugSignals_19}; // @[Fringe.scala 179:22:@61511.4]
  assign regs_io_argOuts_37_bits = {{32'd0}, dramArbs_0_io_debugSignals_20}; // @[Fringe.scala 179:22:@61513.4]
  assign regs_io_argOuts_38_bits = {{32'd0}, dramArbs_0_io_debugSignals_21}; // @[Fringe.scala 179:22:@61515.4]
  assign regs_io_argOuts_39_bits = {{32'd0}, dramArbs_0_io_debugSignals_22}; // @[Fringe.scala 179:22:@61517.4]
  assign regs_io_argOuts_40_bits = {{32'd0}, dramArbs_0_io_debugSignals_23}; // @[Fringe.scala 179:22:@61519.4]
  assign regs_io_argOuts_41_bits = {{32'd0}, dramArbs_0_io_debugSignals_24}; // @[Fringe.scala 179:22:@61521.4]
  assign regs_io_argOuts_42_bits = {{32'd0}, dramArbs_0_io_debugSignals_25}; // @[Fringe.scala 179:22:@61523.4]
  assign regs_io_argOuts_43_bits = {{32'd0}, dramArbs_0_io_debugSignals_26}; // @[Fringe.scala 179:22:@61525.4]
  assign regs_io_argOuts_44_bits = {{32'd0}, dramArbs_0_io_debugSignals_27}; // @[Fringe.scala 179:22:@61527.4]
  assign regs_io_argOuts_45_bits = {{32'd0}, dramArbs_0_io_debugSignals_28}; // @[Fringe.scala 179:22:@61529.4]
  assign regs_io_argOuts_46_bits = {{32'd0}, dramArbs_0_io_debugSignals_29}; // @[Fringe.scala 179:22:@61531.4]
  assign regs_io_argOuts_57_bits = {{32'd0}, dramArbs_0_io_debugSignals_40}; // @[Fringe.scala 179:22:@61553.4]
  assign timeoutCtr_clock = clock; // @[:@61373.4]
  assign timeoutCtr_reset = reset; // @[:@61374.4]
  assign timeoutCtr_io_enable = _T_921 & _T_925; // @[Fringe.scala 149:24:@61388.4]
  assign depulser_clock = clock; // @[:@61391.4]
  assign depulser_reset = reset; // @[:@61392.4]
  assign depulser_io_in = io_done | timeoutCtr_io_done; // @[Fringe.scala 155:18:@61397.4]
  assign depulser_io_rst = _T_936[0]; // @[Fringe.scala 156:19:@61399.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_943 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1468 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_943 <= 1'h0;
    end else begin
      _T_943 <= heap_io_host_0_req_valid;
    end
    if (reset) begin
      _T_1468 <= 1'h0;
    end else begin
      _T_1468 <= _T_1465;
    end
  end
endmodule
module AXI4LiteToRFBridgeKCU1500( // @[:@62776.2]
  input         clock, // @[:@62777.4]
  input         reset, // @[:@62778.4]
  input  [31:0] io_S_AXI_AWADDR, // @[:@62779.4]
  input  [2:0]  io_S_AXI_AWPROT, // @[:@62779.4]
  input         io_S_AXI_AWVALID, // @[:@62779.4]
  output        io_S_AXI_AWREADY, // @[:@62779.4]
  input  [31:0] io_S_AXI_ARADDR, // @[:@62779.4]
  input  [2:0]  io_S_AXI_ARPROT, // @[:@62779.4]
  input         io_S_AXI_ARVALID, // @[:@62779.4]
  output        io_S_AXI_ARREADY, // @[:@62779.4]
  input  [31:0] io_S_AXI_WDATA, // @[:@62779.4]
  input  [3:0]  io_S_AXI_WSTRB, // @[:@62779.4]
  input         io_S_AXI_WVALID, // @[:@62779.4]
  output        io_S_AXI_WREADY, // @[:@62779.4]
  output [31:0] io_S_AXI_RDATA, // @[:@62779.4]
  output [1:0]  io_S_AXI_RRESP, // @[:@62779.4]
  output        io_S_AXI_RVALID, // @[:@62779.4]
  input         io_S_AXI_RREADY, // @[:@62779.4]
  output [1:0]  io_S_AXI_BRESP, // @[:@62779.4]
  output        io_S_AXI_BVALID, // @[:@62779.4]
  input         io_S_AXI_BREADY, // @[:@62779.4]
  output [31:0] io_raddr, // @[:@62779.4]
  output        io_wen, // @[:@62779.4]
  output [31:0] io_waddr, // @[:@62779.4]
  output [31:0] io_wdata, // @[:@62779.4]
  input  [31:0] io_rdata // @[:@62779.4]
);
  wire [31:0] d_rf_rdata; // @[AXI4LiteToRFBridge.scala 109:17:@62781.4]
  wire [31:0] d_rf_wdata; // @[AXI4LiteToRFBridge.scala 109:17:@62781.4]
  wire [31:0] d_rf_waddr; // @[AXI4LiteToRFBridge.scala 109:17:@62781.4]
  wire  d_rf_wen; // @[AXI4LiteToRFBridge.scala 109:17:@62781.4]
  wire [31:0] d_rf_raddr; // @[AXI4LiteToRFBridge.scala 109:17:@62781.4]
  wire  d_S_AXI_ARESETN; // @[AXI4LiteToRFBridge.scala 109:17:@62781.4]
  wire  d_S_AXI_ACLK; // @[AXI4LiteToRFBridge.scala 109:17:@62781.4]
  wire [31:0] d_S_AXI_AWADDR; // @[AXI4LiteToRFBridge.scala 109:17:@62781.4]
  wire [2:0] d_S_AXI_AWPROT; // @[AXI4LiteToRFBridge.scala 109:17:@62781.4]
  wire  d_S_AXI_AWVALID; // @[AXI4LiteToRFBridge.scala 109:17:@62781.4]
  wire  d_S_AXI_AWREADY; // @[AXI4LiteToRFBridge.scala 109:17:@62781.4]
  wire [31:0] d_S_AXI_ARADDR; // @[AXI4LiteToRFBridge.scala 109:17:@62781.4]
  wire [2:0] d_S_AXI_ARPROT; // @[AXI4LiteToRFBridge.scala 109:17:@62781.4]
  wire  d_S_AXI_ARVALID; // @[AXI4LiteToRFBridge.scala 109:17:@62781.4]
  wire  d_S_AXI_ARREADY; // @[AXI4LiteToRFBridge.scala 109:17:@62781.4]
  wire [31:0] d_S_AXI_WDATA; // @[AXI4LiteToRFBridge.scala 109:17:@62781.4]
  wire [3:0] d_S_AXI_WSTRB; // @[AXI4LiteToRFBridge.scala 109:17:@62781.4]
  wire  d_S_AXI_WVALID; // @[AXI4LiteToRFBridge.scala 109:17:@62781.4]
  wire  d_S_AXI_WREADY; // @[AXI4LiteToRFBridge.scala 109:17:@62781.4]
  wire [31:0] d_S_AXI_RDATA; // @[AXI4LiteToRFBridge.scala 109:17:@62781.4]
  wire [1:0] d_S_AXI_RRESP; // @[AXI4LiteToRFBridge.scala 109:17:@62781.4]
  wire  d_S_AXI_RVALID; // @[AXI4LiteToRFBridge.scala 109:17:@62781.4]
  wire  d_S_AXI_RREADY; // @[AXI4LiteToRFBridge.scala 109:17:@62781.4]
  wire [1:0] d_S_AXI_BRESP; // @[AXI4LiteToRFBridge.scala 109:17:@62781.4]
  wire  d_S_AXI_BVALID; // @[AXI4LiteToRFBridge.scala 109:17:@62781.4]
  wire  d_S_AXI_BREADY; // @[AXI4LiteToRFBridge.scala 109:17:@62781.4]
  AXI4LiteToRFBridgeVerilog d ( // @[AXI4LiteToRFBridge.scala 109:17:@62781.4]
    .rf_rdata(d_rf_rdata),
    .rf_wdata(d_rf_wdata),
    .rf_waddr(d_rf_waddr),
    .rf_wen(d_rf_wen),
    .rf_raddr(d_rf_raddr),
    .S_AXI_ARESETN(d_S_AXI_ARESETN),
    .S_AXI_ACLK(d_S_AXI_ACLK),
    .S_AXI_AWADDR(d_S_AXI_AWADDR),
    .S_AXI_AWPROT(d_S_AXI_AWPROT),
    .S_AXI_AWVALID(d_S_AXI_AWVALID),
    .S_AXI_AWREADY(d_S_AXI_AWREADY),
    .S_AXI_ARADDR(d_S_AXI_ARADDR),
    .S_AXI_ARPROT(d_S_AXI_ARPROT),
    .S_AXI_ARVALID(d_S_AXI_ARVALID),
    .S_AXI_ARREADY(d_S_AXI_ARREADY),
    .S_AXI_WDATA(d_S_AXI_WDATA),
    .S_AXI_WSTRB(d_S_AXI_WSTRB),
    .S_AXI_WVALID(d_S_AXI_WVALID),
    .S_AXI_WREADY(d_S_AXI_WREADY),
    .S_AXI_RDATA(d_S_AXI_RDATA),
    .S_AXI_RRESP(d_S_AXI_RRESP),
    .S_AXI_RVALID(d_S_AXI_RVALID),
    .S_AXI_RREADY(d_S_AXI_RREADY),
    .S_AXI_BRESP(d_S_AXI_BRESP),
    .S_AXI_BVALID(d_S_AXI_BVALID),
    .S_AXI_BREADY(d_S_AXI_BREADY)
  );
  assign io_S_AXI_AWREADY = d_S_AXI_AWREADY; // @[AXI4LiteToRFBridge.scala 111:14:@62805.4]
  assign io_S_AXI_ARREADY = d_S_AXI_ARREADY; // @[AXI4LiteToRFBridge.scala 111:14:@62801.4]
  assign io_S_AXI_WREADY = d_S_AXI_WREADY; // @[AXI4LiteToRFBridge.scala 111:14:@62797.4]
  assign io_S_AXI_RDATA = d_S_AXI_RDATA; // @[AXI4LiteToRFBridge.scala 111:14:@62796.4]
  assign io_S_AXI_RRESP = d_S_AXI_RRESP; // @[AXI4LiteToRFBridge.scala 111:14:@62795.4]
  assign io_S_AXI_RVALID = d_S_AXI_RVALID; // @[AXI4LiteToRFBridge.scala 111:14:@62794.4]
  assign io_S_AXI_BRESP = d_S_AXI_BRESP; // @[AXI4LiteToRFBridge.scala 111:14:@62792.4]
  assign io_S_AXI_BVALID = d_S_AXI_BVALID; // @[AXI4LiteToRFBridge.scala 111:14:@62791.4]
  assign io_raddr = d_rf_raddr; // @[AXI4LiteToRFBridge.scala 115:12:@62813.4]
  assign io_wen = d_rf_wen; // @[AXI4LiteToRFBridge.scala 118:12:@62816.4]
  assign io_waddr = d_rf_waddr; // @[AXI4LiteToRFBridge.scala 116:12:@62814.4]
  assign io_wdata = d_rf_wdata; // @[AXI4LiteToRFBridge.scala 117:12:@62815.4]
  assign d_rf_rdata = io_rdata; // @[AXI4LiteToRFBridge.scala 119:17:@62817.4]
  assign d_S_AXI_ARESETN = ~ reset; // @[AXI4LiteToRFBridge.scala 113:22:@62812.4]
  assign d_S_AXI_ACLK = clock; // @[AXI4LiteToRFBridge.scala 112:19:@62809.4]
  assign d_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[AXI4LiteToRFBridge.scala 111:14:@62808.4]
  assign d_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[AXI4LiteToRFBridge.scala 111:14:@62807.4]
  assign d_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[AXI4LiteToRFBridge.scala 111:14:@62806.4]
  assign d_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[AXI4LiteToRFBridge.scala 111:14:@62804.4]
  assign d_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[AXI4LiteToRFBridge.scala 111:14:@62803.4]
  assign d_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[AXI4LiteToRFBridge.scala 111:14:@62802.4]
  assign d_S_AXI_WDATA = io_S_AXI_WDATA; // @[AXI4LiteToRFBridge.scala 111:14:@62800.4]
  assign d_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[AXI4LiteToRFBridge.scala 111:14:@62799.4]
  assign d_S_AXI_WVALID = io_S_AXI_WVALID; // @[AXI4LiteToRFBridge.scala 111:14:@62798.4]
  assign d_S_AXI_RREADY = io_S_AXI_RREADY; // @[AXI4LiteToRFBridge.scala 111:14:@62793.4]
  assign d_S_AXI_BREADY = io_S_AXI_BREADY; // @[AXI4LiteToRFBridge.scala 111:14:@62790.4]
endmodule
module MAGToAXI4Bridge( // @[:@62819.2]
  output         io_in_cmd_ready, // @[:@62822.4]
  input          io_in_cmd_valid, // @[:@62822.4]
  input  [63:0]  io_in_cmd_bits_addr, // @[:@62822.4]
  input  [31:0]  io_in_cmd_bits_size, // @[:@62822.4]
  input  [31:0]  io_in_cmd_bits_tag, // @[:@62822.4]
  output         io_in_wdata_ready, // @[:@62822.4]
  input          io_in_wdata_bits_wlast, // @[:@62822.4]
  input          io_in_rresp_ready, // @[:@62822.4]
  output         io_in_rresp_valid, // @[:@62822.4]
  output [31:0]  io_in_rresp_bits_rdata_0, // @[:@62822.4]
  output [31:0]  io_in_rresp_bits_rdata_1, // @[:@62822.4]
  output [31:0]  io_in_rresp_bits_rdata_2, // @[:@62822.4]
  output [31:0]  io_in_rresp_bits_rdata_3, // @[:@62822.4]
  output [31:0]  io_in_rresp_bits_rdata_4, // @[:@62822.4]
  output [31:0]  io_in_rresp_bits_rdata_5, // @[:@62822.4]
  output [31:0]  io_in_rresp_bits_rdata_6, // @[:@62822.4]
  output [31:0]  io_in_rresp_bits_rdata_7, // @[:@62822.4]
  output [31:0]  io_in_rresp_bits_rdata_8, // @[:@62822.4]
  output [31:0]  io_in_rresp_bits_rdata_9, // @[:@62822.4]
  output [31:0]  io_in_rresp_bits_rdata_10, // @[:@62822.4]
  output [31:0]  io_in_rresp_bits_rdata_11, // @[:@62822.4]
  output [31:0]  io_in_rresp_bits_rdata_12, // @[:@62822.4]
  output [31:0]  io_in_rresp_bits_rdata_13, // @[:@62822.4]
  output [31:0]  io_in_rresp_bits_rdata_14, // @[:@62822.4]
  output [31:0]  io_in_rresp_bits_rdata_15, // @[:@62822.4]
  output [31:0]  io_in_rresp_bits_tag, // @[:@62822.4]
  input          io_in_wresp_ready, // @[:@62822.4]
  output         io_in_wresp_valid, // @[:@62822.4]
  output [31:0]  io_in_wresp_bits_tag, // @[:@62822.4]
  output [3:0]   io_M_AXI_AWID, // @[:@62822.4]
  output [31:0]  io_M_AXI_AWADDR, // @[:@62822.4]
  output [7:0]   io_M_AXI_AWLEN, // @[:@62822.4]
  output [3:0]   io_M_AXI_ARID, // @[:@62822.4]
  output [31:0]  io_M_AXI_ARADDR, // @[:@62822.4]
  output [7:0]   io_M_AXI_ARLEN, // @[:@62822.4]
  output         io_M_AXI_ARVALID, // @[:@62822.4]
  input          io_M_AXI_ARREADY, // @[:@62822.4]
  output         io_M_AXI_WLAST, // @[:@62822.4]
  input          io_M_AXI_WREADY, // @[:@62822.4]
  input  [3:0]   io_M_AXI_RID, // @[:@62822.4]
  input  [511:0] io_M_AXI_RDATA, // @[:@62822.4]
  input          io_M_AXI_RVALID, // @[:@62822.4]
  output         io_M_AXI_RREADY, // @[:@62822.4]
  input  [3:0]   io_M_AXI_BID, // @[:@62822.4]
  input          io_M_AXI_BVALID, // @[:@62822.4]
  output         io_M_AXI_BREADY // @[:@62822.4]
);
  wire [32:0] _T_218; // @[MAGToAXI4Bridge.scala 27:29:@62979.4]
  wire [32:0] _T_219; // @[MAGToAXI4Bridge.scala 27:29:@62980.4]
  wire [31:0] _T_220; // @[MAGToAXI4Bridge.scala 27:29:@62981.4]
  assign _T_218 = io_in_cmd_bits_size - 32'h1; // @[MAGToAXI4Bridge.scala 27:29:@62979.4]
  assign _T_219 = $unsigned(_T_218); // @[MAGToAXI4Bridge.scala 27:29:@62980.4]
  assign _T_220 = _T_219[31:0]; // @[MAGToAXI4Bridge.scala 27:29:@62981.4]
  assign io_in_cmd_ready = io_M_AXI_ARREADY; // @[MAGToAXI4Bridge.scala 36:21:@62993.4]
  assign io_in_wdata_ready = io_M_AXI_WREADY; // @[MAGToAXI4Bridge.scala 56:21:@63090.4]
  assign io_in_rresp_valid = io_M_AXI_RVALID; // @[MAGToAXI4Bridge.scala 70:21:@63142.4]
  assign io_in_rresp_bits_rdata_0 = io_M_AXI_RDATA[31:0]; // @[MAGToAXI4Bridge.scala 62:26:@63124.4]
  assign io_in_rresp_bits_rdata_1 = io_M_AXI_RDATA[63:32]; // @[MAGToAXI4Bridge.scala 62:26:@63125.4]
  assign io_in_rresp_bits_rdata_2 = io_M_AXI_RDATA[95:64]; // @[MAGToAXI4Bridge.scala 62:26:@63126.4]
  assign io_in_rresp_bits_rdata_3 = io_M_AXI_RDATA[127:96]; // @[MAGToAXI4Bridge.scala 62:26:@63127.4]
  assign io_in_rresp_bits_rdata_4 = io_M_AXI_RDATA[159:128]; // @[MAGToAXI4Bridge.scala 62:26:@63128.4]
  assign io_in_rresp_bits_rdata_5 = io_M_AXI_RDATA[191:160]; // @[MAGToAXI4Bridge.scala 62:26:@63129.4]
  assign io_in_rresp_bits_rdata_6 = io_M_AXI_RDATA[223:192]; // @[MAGToAXI4Bridge.scala 62:26:@63130.4]
  assign io_in_rresp_bits_rdata_7 = io_M_AXI_RDATA[255:224]; // @[MAGToAXI4Bridge.scala 62:26:@63131.4]
  assign io_in_rresp_bits_rdata_8 = io_M_AXI_RDATA[287:256]; // @[MAGToAXI4Bridge.scala 62:26:@63132.4]
  assign io_in_rresp_bits_rdata_9 = io_M_AXI_RDATA[319:288]; // @[MAGToAXI4Bridge.scala 62:26:@63133.4]
  assign io_in_rresp_bits_rdata_10 = io_M_AXI_RDATA[351:320]; // @[MAGToAXI4Bridge.scala 62:26:@63134.4]
  assign io_in_rresp_bits_rdata_11 = io_M_AXI_RDATA[383:352]; // @[MAGToAXI4Bridge.scala 62:26:@63135.4]
  assign io_in_rresp_bits_rdata_12 = io_M_AXI_RDATA[415:384]; // @[MAGToAXI4Bridge.scala 62:26:@63136.4]
  assign io_in_rresp_bits_rdata_13 = io_M_AXI_RDATA[447:416]; // @[MAGToAXI4Bridge.scala 62:26:@63137.4]
  assign io_in_rresp_bits_rdata_14 = io_M_AXI_RDATA[479:448]; // @[MAGToAXI4Bridge.scala 62:26:@63138.4]
  assign io_in_rresp_bits_rdata_15 = io_M_AXI_RDATA[511:480]; // @[MAGToAXI4Bridge.scala 62:26:@63139.4]
  assign io_in_rresp_bits_tag = {{28'd0}, io_M_AXI_RID}; // @[MAGToAXI4Bridge.scala 73:24:@63144.4]
  assign io_in_wresp_valid = io_M_AXI_BVALID; // @[MAGToAXI4Bridge.scala 71:21:@63143.4]
  assign io_in_wresp_bits_tag = {{28'd0}, io_M_AXI_BID}; // @[MAGToAXI4Bridge.scala 74:24:@63145.4]
  assign io_M_AXI_AWID = io_in_cmd_bits_tag[3:0]; // @[MAGToAXI4Bridge.scala 39:21:@62994.4]
  assign io_M_AXI_AWADDR = io_in_cmd_bits_addr[31:0]; // @[MAGToAXI4Bridge.scala 40:21:@62995.4]
  assign io_M_AXI_AWLEN = _T_220[7:0]; // @[MAGToAXI4Bridge.scala 41:21:@62999.4]
  assign io_M_AXI_ARID = io_in_cmd_bits_tag[3:0]; // @[MAGToAXI4Bridge.scala 25:21:@62977.4]
  assign io_M_AXI_ARADDR = io_in_cmd_bits_addr[31:0]; // @[MAGToAXI4Bridge.scala 26:21:@62978.4]
  assign io_M_AXI_ARLEN = _T_220[7:0]; // @[MAGToAXI4Bridge.scala 27:21:@62982.4]
  assign io_M_AXI_ARVALID = io_in_cmd_valid; // @[MAGToAXI4Bridge.scala 35:21:@62991.4]
  assign io_M_AXI_WLAST = io_in_wdata_bits_wlast; // @[MAGToAXI4Bridge.scala 54:21:@63088.4]
  assign io_M_AXI_RREADY = io_in_rresp_ready; // @[MAGToAXI4Bridge.scala 64:19:@63140.4]
  assign io_M_AXI_BREADY = io_in_wresp_ready; // @[MAGToAXI4Bridge.scala 67:19:@63141.4]
endmodule
module FringeZynq( // @[:@63147.2]
  input          clock, // @[:@63148.4]
  input          reset, // @[:@63149.4]
  input  [31:0]  io_S_AXI_AWADDR, // @[:@63150.4]
  input  [2:0]   io_S_AXI_AWPROT, // @[:@63150.4]
  input          io_S_AXI_AWVALID, // @[:@63150.4]
  output         io_S_AXI_AWREADY, // @[:@63150.4]
  input  [31:0]  io_S_AXI_ARADDR, // @[:@63150.4]
  input  [2:0]   io_S_AXI_ARPROT, // @[:@63150.4]
  input          io_S_AXI_ARVALID, // @[:@63150.4]
  output         io_S_AXI_ARREADY, // @[:@63150.4]
  input  [31:0]  io_S_AXI_WDATA, // @[:@63150.4]
  input  [3:0]   io_S_AXI_WSTRB, // @[:@63150.4]
  input          io_S_AXI_WVALID, // @[:@63150.4]
  output         io_S_AXI_WREADY, // @[:@63150.4]
  output [31:0]  io_S_AXI_RDATA, // @[:@63150.4]
  output [1:0]   io_S_AXI_RRESP, // @[:@63150.4]
  output         io_S_AXI_RVALID, // @[:@63150.4]
  input          io_S_AXI_RREADY, // @[:@63150.4]
  output [1:0]   io_S_AXI_BRESP, // @[:@63150.4]
  output         io_S_AXI_BVALID, // @[:@63150.4]
  input          io_S_AXI_BREADY, // @[:@63150.4]
  output [3:0]   io_M_AXI_0_AWID, // @[:@63150.4]
  output [31:0]  io_M_AXI_0_AWADDR, // @[:@63150.4]
  output [7:0]   io_M_AXI_0_AWLEN, // @[:@63150.4]
  output [3:0]   io_M_AXI_0_ARID, // @[:@63150.4]
  output [31:0]  io_M_AXI_0_ARADDR, // @[:@63150.4]
  output [7:0]   io_M_AXI_0_ARLEN, // @[:@63150.4]
  output         io_M_AXI_0_ARVALID, // @[:@63150.4]
  input          io_M_AXI_0_ARREADY, // @[:@63150.4]
  output         io_M_AXI_0_WLAST, // @[:@63150.4]
  input          io_M_AXI_0_WREADY, // @[:@63150.4]
  input  [3:0]   io_M_AXI_0_RID, // @[:@63150.4]
  input  [511:0] io_M_AXI_0_RDATA, // @[:@63150.4]
  input          io_M_AXI_0_RVALID, // @[:@63150.4]
  output         io_M_AXI_0_RREADY, // @[:@63150.4]
  input  [3:0]   io_M_AXI_0_BID, // @[:@63150.4]
  input          io_M_AXI_0_BVALID, // @[:@63150.4]
  output         io_M_AXI_0_BREADY, // @[:@63150.4]
  output         io_enable, // @[:@63150.4]
  input          io_done, // @[:@63150.4]
  output         io_reset, // @[:@63150.4]
  output [63:0]  io_argIns_0, // @[:@63150.4]
  input          io_argOuts_0_valid, // @[:@63150.4]
  input  [63:0]  io_argOuts_0_bits, // @[:@63150.4]
  input          io_argOuts_1_valid, // @[:@63150.4]
  input  [63:0]  io_argOuts_1_bits, // @[:@63150.4]
  input          io_argOuts_2_valid, // @[:@63150.4]
  input  [63:0]  io_argOuts_2_bits, // @[:@63150.4]
  input          io_argOuts_3_valid, // @[:@63150.4]
  input  [63:0]  io_argOuts_3_bits, // @[:@63150.4]
  input          io_argOuts_4_valid, // @[:@63150.4]
  input  [63:0]  io_argOuts_4_bits, // @[:@63150.4]
  input          io_argOuts_5_valid, // @[:@63150.4]
  input  [63:0]  io_argOuts_5_bits, // @[:@63150.4]
  input          io_argOuts_6_valid, // @[:@63150.4]
  input  [63:0]  io_argOuts_6_bits, // @[:@63150.4]
  input          io_argOuts_7_valid, // @[:@63150.4]
  input  [63:0]  io_argOuts_7_bits, // @[:@63150.4]
  input          io_argOuts_8_valid, // @[:@63150.4]
  input  [63:0]  io_argOuts_8_bits, // @[:@63150.4]
  input          io_argOuts_9_valid, // @[:@63150.4]
  input  [63:0]  io_argOuts_9_bits, // @[:@63150.4]
  input          io_argOuts_10_valid, // @[:@63150.4]
  input  [63:0]  io_argOuts_10_bits, // @[:@63150.4]
  input          io_argOuts_11_valid, // @[:@63150.4]
  input  [63:0]  io_argOuts_11_bits, // @[:@63150.4]
  input          io_argOuts_12_valid, // @[:@63150.4]
  input  [63:0]  io_argOuts_12_bits, // @[:@63150.4]
  input          io_argOuts_13_valid, // @[:@63150.4]
  input  [63:0]  io_argOuts_13_bits, // @[:@63150.4]
  input          io_argOuts_14_valid, // @[:@63150.4]
  input  [63:0]  io_argOuts_14_bits, // @[:@63150.4]
  input          io_argOuts_15_valid, // @[:@63150.4]
  input  [63:0]  io_argOuts_15_bits, // @[:@63150.4]
  output         io_memStreams_loads_0_cmd_ready, // @[:@63150.4]
  input          io_memStreams_loads_0_cmd_valid, // @[:@63150.4]
  input  [63:0]  io_memStreams_loads_0_cmd_bits_addr, // @[:@63150.4]
  input  [31:0]  io_memStreams_loads_0_cmd_bits_size, // @[:@63150.4]
  input          io_memStreams_loads_0_data_ready, // @[:@63150.4]
  output         io_memStreams_loads_0_data_valid, // @[:@63150.4]
  output [31:0]  io_memStreams_loads_0_data_bits_rdata_0, // @[:@63150.4]
  input          io_memStreams_stores_0_cmd_valid, // @[:@63150.4]
  input  [63:0]  io_memStreams_stores_0_cmd_bits_addr, // @[:@63150.4]
  input  [31:0]  io_memStreams_stores_0_cmd_bits_size, // @[:@63150.4]
  input          io_memStreams_stores_0_data_valid, // @[:@63150.4]
  input  [31:0]  io_memStreams_stores_0_data_bits_wdata_0, // @[:@63150.4]
  input  [15:0]  io_memStreams_stores_0_data_bits_wstrb, // @[:@63150.4]
  input          io_heap_0_req_valid, // @[:@63150.4]
  input          io_heap_0_req_bits_allocDealloc, // @[:@63150.4]
  input  [63:0]  io_heap_0_req_bits_sizeAddr, // @[:@63150.4]
  output         io_heap_0_resp_valid, // @[:@63150.4]
  output         io_heap_0_resp_bits_allocDealloc, // @[:@63150.4]
  output [63:0]  io_heap_0_resp_bits_sizeAddr // @[:@63150.4]
);
  wire  fringeCommon_clock; // @[FringeZynq.scala 68:28:@63557.4]
  wire  fringeCommon_reset; // @[FringeZynq.scala 68:28:@63557.4]
  wire [31:0] fringeCommon_io_raddr; // @[FringeZynq.scala 68:28:@63557.4]
  wire  fringeCommon_io_wen; // @[FringeZynq.scala 68:28:@63557.4]
  wire [31:0] fringeCommon_io_waddr; // @[FringeZynq.scala 68:28:@63557.4]
  wire [63:0] fringeCommon_io_wdata; // @[FringeZynq.scala 68:28:@63557.4]
  wire [63:0] fringeCommon_io_rdata; // @[FringeZynq.scala 68:28:@63557.4]
  wire  fringeCommon_io_enable; // @[FringeZynq.scala 68:28:@63557.4]
  wire  fringeCommon_io_done; // @[FringeZynq.scala 68:28:@63557.4]
  wire  fringeCommon_io_reset; // @[FringeZynq.scala 68:28:@63557.4]
  wire [63:0] fringeCommon_io_argIns_0; // @[FringeZynq.scala 68:28:@63557.4]
  wire  fringeCommon_io_argOuts_0_valid; // @[FringeZynq.scala 68:28:@63557.4]
  wire [63:0] fringeCommon_io_argOuts_0_bits; // @[FringeZynq.scala 68:28:@63557.4]
  wire  fringeCommon_io_argOuts_1_valid; // @[FringeZynq.scala 68:28:@63557.4]
  wire [63:0] fringeCommon_io_argOuts_1_bits; // @[FringeZynq.scala 68:28:@63557.4]
  wire  fringeCommon_io_argOuts_2_valid; // @[FringeZynq.scala 68:28:@63557.4]
  wire [63:0] fringeCommon_io_argOuts_2_bits; // @[FringeZynq.scala 68:28:@63557.4]
  wire  fringeCommon_io_argOuts_3_valid; // @[FringeZynq.scala 68:28:@63557.4]
  wire [63:0] fringeCommon_io_argOuts_3_bits; // @[FringeZynq.scala 68:28:@63557.4]
  wire  fringeCommon_io_argOuts_4_valid; // @[FringeZynq.scala 68:28:@63557.4]
  wire [63:0] fringeCommon_io_argOuts_4_bits; // @[FringeZynq.scala 68:28:@63557.4]
  wire  fringeCommon_io_argOuts_5_valid; // @[FringeZynq.scala 68:28:@63557.4]
  wire [63:0] fringeCommon_io_argOuts_5_bits; // @[FringeZynq.scala 68:28:@63557.4]
  wire  fringeCommon_io_argOuts_6_valid; // @[FringeZynq.scala 68:28:@63557.4]
  wire [63:0] fringeCommon_io_argOuts_6_bits; // @[FringeZynq.scala 68:28:@63557.4]
  wire  fringeCommon_io_argOuts_7_valid; // @[FringeZynq.scala 68:28:@63557.4]
  wire [63:0] fringeCommon_io_argOuts_7_bits; // @[FringeZynq.scala 68:28:@63557.4]
  wire  fringeCommon_io_argOuts_8_valid; // @[FringeZynq.scala 68:28:@63557.4]
  wire [63:0] fringeCommon_io_argOuts_8_bits; // @[FringeZynq.scala 68:28:@63557.4]
  wire  fringeCommon_io_argOuts_9_valid; // @[FringeZynq.scala 68:28:@63557.4]
  wire [63:0] fringeCommon_io_argOuts_9_bits; // @[FringeZynq.scala 68:28:@63557.4]
  wire  fringeCommon_io_argOuts_10_valid; // @[FringeZynq.scala 68:28:@63557.4]
  wire [63:0] fringeCommon_io_argOuts_10_bits; // @[FringeZynq.scala 68:28:@63557.4]
  wire  fringeCommon_io_argOuts_11_valid; // @[FringeZynq.scala 68:28:@63557.4]
  wire [63:0] fringeCommon_io_argOuts_11_bits; // @[FringeZynq.scala 68:28:@63557.4]
  wire  fringeCommon_io_argOuts_12_valid; // @[FringeZynq.scala 68:28:@63557.4]
  wire [63:0] fringeCommon_io_argOuts_12_bits; // @[FringeZynq.scala 68:28:@63557.4]
  wire  fringeCommon_io_argOuts_13_valid; // @[FringeZynq.scala 68:28:@63557.4]
  wire [63:0] fringeCommon_io_argOuts_13_bits; // @[FringeZynq.scala 68:28:@63557.4]
  wire  fringeCommon_io_argOuts_14_valid; // @[FringeZynq.scala 68:28:@63557.4]
  wire [63:0] fringeCommon_io_argOuts_14_bits; // @[FringeZynq.scala 68:28:@63557.4]
  wire  fringeCommon_io_argOuts_15_valid; // @[FringeZynq.scala 68:28:@63557.4]
  wire [63:0] fringeCommon_io_argOuts_15_bits; // @[FringeZynq.scala 68:28:@63557.4]
  wire  fringeCommon_io_memStreams_loads_0_cmd_ready; // @[FringeZynq.scala 68:28:@63557.4]
  wire  fringeCommon_io_memStreams_loads_0_cmd_valid; // @[FringeZynq.scala 68:28:@63557.4]
  wire [63:0] fringeCommon_io_memStreams_loads_0_cmd_bits_addr; // @[FringeZynq.scala 68:28:@63557.4]
  wire [31:0] fringeCommon_io_memStreams_loads_0_cmd_bits_size; // @[FringeZynq.scala 68:28:@63557.4]
  wire  fringeCommon_io_memStreams_loads_0_data_ready; // @[FringeZynq.scala 68:28:@63557.4]
  wire  fringeCommon_io_memStreams_loads_0_data_valid; // @[FringeZynq.scala 68:28:@63557.4]
  wire [31:0] fringeCommon_io_memStreams_loads_0_data_bits_rdata_0; // @[FringeZynq.scala 68:28:@63557.4]
  wire  fringeCommon_io_memStreams_stores_0_cmd_valid; // @[FringeZynq.scala 68:28:@63557.4]
  wire [63:0] fringeCommon_io_memStreams_stores_0_cmd_bits_addr; // @[FringeZynq.scala 68:28:@63557.4]
  wire [31:0] fringeCommon_io_memStreams_stores_0_cmd_bits_size; // @[FringeZynq.scala 68:28:@63557.4]
  wire  fringeCommon_io_memStreams_stores_0_data_valid; // @[FringeZynq.scala 68:28:@63557.4]
  wire [31:0] fringeCommon_io_memStreams_stores_0_data_bits_wdata_0; // @[FringeZynq.scala 68:28:@63557.4]
  wire [15:0] fringeCommon_io_memStreams_stores_0_data_bits_wstrb; // @[FringeZynq.scala 68:28:@63557.4]
  wire  fringeCommon_io_dram_0_cmd_ready; // @[FringeZynq.scala 68:28:@63557.4]
  wire  fringeCommon_io_dram_0_cmd_valid; // @[FringeZynq.scala 68:28:@63557.4]
  wire [63:0] fringeCommon_io_dram_0_cmd_bits_addr; // @[FringeZynq.scala 68:28:@63557.4]
  wire [31:0] fringeCommon_io_dram_0_cmd_bits_size; // @[FringeZynq.scala 68:28:@63557.4]
  wire [31:0] fringeCommon_io_dram_0_cmd_bits_tag; // @[FringeZynq.scala 68:28:@63557.4]
  wire  fringeCommon_io_dram_0_wdata_ready; // @[FringeZynq.scala 68:28:@63557.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wlast; // @[FringeZynq.scala 68:28:@63557.4]
  wire  fringeCommon_io_dram_0_rresp_ready; // @[FringeZynq.scala 68:28:@63557.4]
  wire  fringeCommon_io_dram_0_rresp_valid; // @[FringeZynq.scala 68:28:@63557.4]
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_rdata_0; // @[FringeZynq.scala 68:28:@63557.4]
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_rdata_1; // @[FringeZynq.scala 68:28:@63557.4]
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_rdata_2; // @[FringeZynq.scala 68:28:@63557.4]
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_rdata_3; // @[FringeZynq.scala 68:28:@63557.4]
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_rdata_4; // @[FringeZynq.scala 68:28:@63557.4]
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_rdata_5; // @[FringeZynq.scala 68:28:@63557.4]
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_rdata_6; // @[FringeZynq.scala 68:28:@63557.4]
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_rdata_7; // @[FringeZynq.scala 68:28:@63557.4]
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_rdata_8; // @[FringeZynq.scala 68:28:@63557.4]
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_rdata_9; // @[FringeZynq.scala 68:28:@63557.4]
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_rdata_10; // @[FringeZynq.scala 68:28:@63557.4]
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_rdata_11; // @[FringeZynq.scala 68:28:@63557.4]
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_rdata_12; // @[FringeZynq.scala 68:28:@63557.4]
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_rdata_13; // @[FringeZynq.scala 68:28:@63557.4]
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_rdata_14; // @[FringeZynq.scala 68:28:@63557.4]
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_rdata_15; // @[FringeZynq.scala 68:28:@63557.4]
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_tag; // @[FringeZynq.scala 68:28:@63557.4]
  wire  fringeCommon_io_dram_0_wresp_ready; // @[FringeZynq.scala 68:28:@63557.4]
  wire  fringeCommon_io_dram_0_wresp_valid; // @[FringeZynq.scala 68:28:@63557.4]
  wire [31:0] fringeCommon_io_dram_0_wresp_bits_tag; // @[FringeZynq.scala 68:28:@63557.4]
  wire  fringeCommon_io_heap_0_req_valid; // @[FringeZynq.scala 68:28:@63557.4]
  wire  fringeCommon_io_heap_0_req_bits_allocDealloc; // @[FringeZynq.scala 68:28:@63557.4]
  wire [63:0] fringeCommon_io_heap_0_req_bits_sizeAddr; // @[FringeZynq.scala 68:28:@63557.4]
  wire  fringeCommon_io_heap_0_resp_valid; // @[FringeZynq.scala 68:28:@63557.4]
  wire  fringeCommon_io_heap_0_resp_bits_allocDealloc; // @[FringeZynq.scala 68:28:@63557.4]
  wire [63:0] fringeCommon_io_heap_0_resp_bits_sizeAddr; // @[FringeZynq.scala 68:28:@63557.4]
  wire  AXI4LiteToRFBridgeKCU1500_clock; // @[FringeZynq.scala 78:31:@64186.4]
  wire  AXI4LiteToRFBridgeKCU1500_reset; // @[FringeZynq.scala 78:31:@64186.4]
  wire [31:0] AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWADDR; // @[FringeZynq.scala 78:31:@64186.4]
  wire [2:0] AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWPROT; // @[FringeZynq.scala 78:31:@64186.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWVALID; // @[FringeZynq.scala 78:31:@64186.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWREADY; // @[FringeZynq.scala 78:31:@64186.4]
  wire [31:0] AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARADDR; // @[FringeZynq.scala 78:31:@64186.4]
  wire [2:0] AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARPROT; // @[FringeZynq.scala 78:31:@64186.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARVALID; // @[FringeZynq.scala 78:31:@64186.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARREADY; // @[FringeZynq.scala 78:31:@64186.4]
  wire [31:0] AXI4LiteToRFBridgeKCU1500_io_S_AXI_WDATA; // @[FringeZynq.scala 78:31:@64186.4]
  wire [3:0] AXI4LiteToRFBridgeKCU1500_io_S_AXI_WSTRB; // @[FringeZynq.scala 78:31:@64186.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_WVALID; // @[FringeZynq.scala 78:31:@64186.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_WREADY; // @[FringeZynq.scala 78:31:@64186.4]
  wire [31:0] AXI4LiteToRFBridgeKCU1500_io_S_AXI_RDATA; // @[FringeZynq.scala 78:31:@64186.4]
  wire [1:0] AXI4LiteToRFBridgeKCU1500_io_S_AXI_RRESP; // @[FringeZynq.scala 78:31:@64186.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_RVALID; // @[FringeZynq.scala 78:31:@64186.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_RREADY; // @[FringeZynq.scala 78:31:@64186.4]
  wire [1:0] AXI4LiteToRFBridgeKCU1500_io_S_AXI_BRESP; // @[FringeZynq.scala 78:31:@64186.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_BVALID; // @[FringeZynq.scala 78:31:@64186.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_BREADY; // @[FringeZynq.scala 78:31:@64186.4]
  wire [31:0] AXI4LiteToRFBridgeKCU1500_io_raddr; // @[FringeZynq.scala 78:31:@64186.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_wen; // @[FringeZynq.scala 78:31:@64186.4]
  wire [31:0] AXI4LiteToRFBridgeKCU1500_io_waddr; // @[FringeZynq.scala 78:31:@64186.4]
  wire [31:0] AXI4LiteToRFBridgeKCU1500_io_wdata; // @[FringeZynq.scala 78:31:@64186.4]
  wire [31:0] AXI4LiteToRFBridgeKCU1500_io_rdata; // @[FringeZynq.scala 78:31:@64186.4]
  wire  MAGToAXI4Bridge_io_in_cmd_ready; // @[FringeZynq.scala 130:27:@64382.4]
  wire  MAGToAXI4Bridge_io_in_cmd_valid; // @[FringeZynq.scala 130:27:@64382.4]
  wire [63:0] MAGToAXI4Bridge_io_in_cmd_bits_addr; // @[FringeZynq.scala 130:27:@64382.4]
  wire [31:0] MAGToAXI4Bridge_io_in_cmd_bits_size; // @[FringeZynq.scala 130:27:@64382.4]
  wire [31:0] MAGToAXI4Bridge_io_in_cmd_bits_tag; // @[FringeZynq.scala 130:27:@64382.4]
  wire  MAGToAXI4Bridge_io_in_wdata_ready; // @[FringeZynq.scala 130:27:@64382.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wlast; // @[FringeZynq.scala 130:27:@64382.4]
  wire  MAGToAXI4Bridge_io_in_rresp_ready; // @[FringeZynq.scala 130:27:@64382.4]
  wire  MAGToAXI4Bridge_io_in_rresp_valid; // @[FringeZynq.scala 130:27:@64382.4]
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_0; // @[FringeZynq.scala 130:27:@64382.4]
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_1; // @[FringeZynq.scala 130:27:@64382.4]
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_2; // @[FringeZynq.scala 130:27:@64382.4]
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_3; // @[FringeZynq.scala 130:27:@64382.4]
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_4; // @[FringeZynq.scala 130:27:@64382.4]
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_5; // @[FringeZynq.scala 130:27:@64382.4]
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_6; // @[FringeZynq.scala 130:27:@64382.4]
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_7; // @[FringeZynq.scala 130:27:@64382.4]
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_8; // @[FringeZynq.scala 130:27:@64382.4]
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_9; // @[FringeZynq.scala 130:27:@64382.4]
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_10; // @[FringeZynq.scala 130:27:@64382.4]
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_11; // @[FringeZynq.scala 130:27:@64382.4]
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_12; // @[FringeZynq.scala 130:27:@64382.4]
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_13; // @[FringeZynq.scala 130:27:@64382.4]
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_14; // @[FringeZynq.scala 130:27:@64382.4]
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_15; // @[FringeZynq.scala 130:27:@64382.4]
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_tag; // @[FringeZynq.scala 130:27:@64382.4]
  wire  MAGToAXI4Bridge_io_in_wresp_ready; // @[FringeZynq.scala 130:27:@64382.4]
  wire  MAGToAXI4Bridge_io_in_wresp_valid; // @[FringeZynq.scala 130:27:@64382.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wresp_bits_tag; // @[FringeZynq.scala 130:27:@64382.4]
  wire [3:0] MAGToAXI4Bridge_io_M_AXI_AWID; // @[FringeZynq.scala 130:27:@64382.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_AWADDR; // @[FringeZynq.scala 130:27:@64382.4]
  wire [7:0] MAGToAXI4Bridge_io_M_AXI_AWLEN; // @[FringeZynq.scala 130:27:@64382.4]
  wire [3:0] MAGToAXI4Bridge_io_M_AXI_ARID; // @[FringeZynq.scala 130:27:@64382.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_ARADDR; // @[FringeZynq.scala 130:27:@64382.4]
  wire [7:0] MAGToAXI4Bridge_io_M_AXI_ARLEN; // @[FringeZynq.scala 130:27:@64382.4]
  wire  MAGToAXI4Bridge_io_M_AXI_ARVALID; // @[FringeZynq.scala 130:27:@64382.4]
  wire  MAGToAXI4Bridge_io_M_AXI_ARREADY; // @[FringeZynq.scala 130:27:@64382.4]
  wire  MAGToAXI4Bridge_io_M_AXI_WLAST; // @[FringeZynq.scala 130:27:@64382.4]
  wire  MAGToAXI4Bridge_io_M_AXI_WREADY; // @[FringeZynq.scala 130:27:@64382.4]
  wire [3:0] MAGToAXI4Bridge_io_M_AXI_RID; // @[FringeZynq.scala 130:27:@64382.4]
  wire [511:0] MAGToAXI4Bridge_io_M_AXI_RDATA; // @[FringeZynq.scala 130:27:@64382.4]
  wire  MAGToAXI4Bridge_io_M_AXI_RVALID; // @[FringeZynq.scala 130:27:@64382.4]
  wire  MAGToAXI4Bridge_io_M_AXI_RREADY; // @[FringeZynq.scala 130:27:@64382.4]
  wire [3:0] MAGToAXI4Bridge_io_M_AXI_BID; // @[FringeZynq.scala 130:27:@64382.4]
  wire  MAGToAXI4Bridge_io_M_AXI_BVALID; // @[FringeZynq.scala 130:27:@64382.4]
  wire  MAGToAXI4Bridge_io_M_AXI_BREADY; // @[FringeZynq.scala 130:27:@64382.4]
  Fringe fringeCommon ( // @[FringeZynq.scala 68:28:@63557.4]
    .clock(fringeCommon_clock),
    .reset(fringeCommon_reset),
    .io_raddr(fringeCommon_io_raddr),
    .io_wen(fringeCommon_io_wen),
    .io_waddr(fringeCommon_io_waddr),
    .io_wdata(fringeCommon_io_wdata),
    .io_rdata(fringeCommon_io_rdata),
    .io_enable(fringeCommon_io_enable),
    .io_done(fringeCommon_io_done),
    .io_reset(fringeCommon_io_reset),
    .io_argIns_0(fringeCommon_io_argIns_0),
    .io_argOuts_0_valid(fringeCommon_io_argOuts_0_valid),
    .io_argOuts_0_bits(fringeCommon_io_argOuts_0_bits),
    .io_argOuts_1_valid(fringeCommon_io_argOuts_1_valid),
    .io_argOuts_1_bits(fringeCommon_io_argOuts_1_bits),
    .io_argOuts_2_valid(fringeCommon_io_argOuts_2_valid),
    .io_argOuts_2_bits(fringeCommon_io_argOuts_2_bits),
    .io_argOuts_3_valid(fringeCommon_io_argOuts_3_valid),
    .io_argOuts_3_bits(fringeCommon_io_argOuts_3_bits),
    .io_argOuts_4_valid(fringeCommon_io_argOuts_4_valid),
    .io_argOuts_4_bits(fringeCommon_io_argOuts_4_bits),
    .io_argOuts_5_valid(fringeCommon_io_argOuts_5_valid),
    .io_argOuts_5_bits(fringeCommon_io_argOuts_5_bits),
    .io_argOuts_6_valid(fringeCommon_io_argOuts_6_valid),
    .io_argOuts_6_bits(fringeCommon_io_argOuts_6_bits),
    .io_argOuts_7_valid(fringeCommon_io_argOuts_7_valid),
    .io_argOuts_7_bits(fringeCommon_io_argOuts_7_bits),
    .io_argOuts_8_valid(fringeCommon_io_argOuts_8_valid),
    .io_argOuts_8_bits(fringeCommon_io_argOuts_8_bits),
    .io_argOuts_9_valid(fringeCommon_io_argOuts_9_valid),
    .io_argOuts_9_bits(fringeCommon_io_argOuts_9_bits),
    .io_argOuts_10_valid(fringeCommon_io_argOuts_10_valid),
    .io_argOuts_10_bits(fringeCommon_io_argOuts_10_bits),
    .io_argOuts_11_valid(fringeCommon_io_argOuts_11_valid),
    .io_argOuts_11_bits(fringeCommon_io_argOuts_11_bits),
    .io_argOuts_12_valid(fringeCommon_io_argOuts_12_valid),
    .io_argOuts_12_bits(fringeCommon_io_argOuts_12_bits),
    .io_argOuts_13_valid(fringeCommon_io_argOuts_13_valid),
    .io_argOuts_13_bits(fringeCommon_io_argOuts_13_bits),
    .io_argOuts_14_valid(fringeCommon_io_argOuts_14_valid),
    .io_argOuts_14_bits(fringeCommon_io_argOuts_14_bits),
    .io_argOuts_15_valid(fringeCommon_io_argOuts_15_valid),
    .io_argOuts_15_bits(fringeCommon_io_argOuts_15_bits),
    .io_memStreams_loads_0_cmd_ready(fringeCommon_io_memStreams_loads_0_cmd_ready),
    .io_memStreams_loads_0_cmd_valid(fringeCommon_io_memStreams_loads_0_cmd_valid),
    .io_memStreams_loads_0_cmd_bits_addr(fringeCommon_io_memStreams_loads_0_cmd_bits_addr),
    .io_memStreams_loads_0_cmd_bits_size(fringeCommon_io_memStreams_loads_0_cmd_bits_size),
    .io_memStreams_loads_0_data_ready(fringeCommon_io_memStreams_loads_0_data_ready),
    .io_memStreams_loads_0_data_valid(fringeCommon_io_memStreams_loads_0_data_valid),
    .io_memStreams_loads_0_data_bits_rdata_0(fringeCommon_io_memStreams_loads_0_data_bits_rdata_0),
    .io_memStreams_stores_0_cmd_valid(fringeCommon_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(fringeCommon_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(fringeCommon_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_valid(fringeCommon_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(fringeCommon_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wstrb(fringeCommon_io_memStreams_stores_0_data_bits_wstrb),
    .io_dram_0_cmd_ready(fringeCommon_io_dram_0_cmd_ready),
    .io_dram_0_cmd_valid(fringeCommon_io_dram_0_cmd_valid),
    .io_dram_0_cmd_bits_addr(fringeCommon_io_dram_0_cmd_bits_addr),
    .io_dram_0_cmd_bits_size(fringeCommon_io_dram_0_cmd_bits_size),
    .io_dram_0_cmd_bits_tag(fringeCommon_io_dram_0_cmd_bits_tag),
    .io_dram_0_wdata_ready(fringeCommon_io_dram_0_wdata_ready),
    .io_dram_0_wdata_bits_wlast(fringeCommon_io_dram_0_wdata_bits_wlast),
    .io_dram_0_rresp_ready(fringeCommon_io_dram_0_rresp_ready),
    .io_dram_0_rresp_valid(fringeCommon_io_dram_0_rresp_valid),
    .io_dram_0_rresp_bits_rdata_0(fringeCommon_io_dram_0_rresp_bits_rdata_0),
    .io_dram_0_rresp_bits_rdata_1(fringeCommon_io_dram_0_rresp_bits_rdata_1),
    .io_dram_0_rresp_bits_rdata_2(fringeCommon_io_dram_0_rresp_bits_rdata_2),
    .io_dram_0_rresp_bits_rdata_3(fringeCommon_io_dram_0_rresp_bits_rdata_3),
    .io_dram_0_rresp_bits_rdata_4(fringeCommon_io_dram_0_rresp_bits_rdata_4),
    .io_dram_0_rresp_bits_rdata_5(fringeCommon_io_dram_0_rresp_bits_rdata_5),
    .io_dram_0_rresp_bits_rdata_6(fringeCommon_io_dram_0_rresp_bits_rdata_6),
    .io_dram_0_rresp_bits_rdata_7(fringeCommon_io_dram_0_rresp_bits_rdata_7),
    .io_dram_0_rresp_bits_rdata_8(fringeCommon_io_dram_0_rresp_bits_rdata_8),
    .io_dram_0_rresp_bits_rdata_9(fringeCommon_io_dram_0_rresp_bits_rdata_9),
    .io_dram_0_rresp_bits_rdata_10(fringeCommon_io_dram_0_rresp_bits_rdata_10),
    .io_dram_0_rresp_bits_rdata_11(fringeCommon_io_dram_0_rresp_bits_rdata_11),
    .io_dram_0_rresp_bits_rdata_12(fringeCommon_io_dram_0_rresp_bits_rdata_12),
    .io_dram_0_rresp_bits_rdata_13(fringeCommon_io_dram_0_rresp_bits_rdata_13),
    .io_dram_0_rresp_bits_rdata_14(fringeCommon_io_dram_0_rresp_bits_rdata_14),
    .io_dram_0_rresp_bits_rdata_15(fringeCommon_io_dram_0_rresp_bits_rdata_15),
    .io_dram_0_rresp_bits_tag(fringeCommon_io_dram_0_rresp_bits_tag),
    .io_dram_0_wresp_ready(fringeCommon_io_dram_0_wresp_ready),
    .io_dram_0_wresp_valid(fringeCommon_io_dram_0_wresp_valid),
    .io_dram_0_wresp_bits_tag(fringeCommon_io_dram_0_wresp_bits_tag),
    .io_heap_0_req_valid(fringeCommon_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(fringeCommon_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(fringeCommon_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(fringeCommon_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(fringeCommon_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(fringeCommon_io_heap_0_resp_bits_sizeAddr)
  );
  AXI4LiteToRFBridgeKCU1500 AXI4LiteToRFBridgeKCU1500 ( // @[FringeZynq.scala 78:31:@64186.4]
    .clock(AXI4LiteToRFBridgeKCU1500_clock),
    .reset(AXI4LiteToRFBridgeKCU1500_reset),
    .io_S_AXI_AWADDR(AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWADDR),
    .io_S_AXI_AWPROT(AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWPROT),
    .io_S_AXI_AWVALID(AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWVALID),
    .io_S_AXI_AWREADY(AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWREADY),
    .io_S_AXI_ARADDR(AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARADDR),
    .io_S_AXI_ARPROT(AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARPROT),
    .io_S_AXI_ARVALID(AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARVALID),
    .io_S_AXI_ARREADY(AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARREADY),
    .io_S_AXI_WDATA(AXI4LiteToRFBridgeKCU1500_io_S_AXI_WDATA),
    .io_S_AXI_WSTRB(AXI4LiteToRFBridgeKCU1500_io_S_AXI_WSTRB),
    .io_S_AXI_WVALID(AXI4LiteToRFBridgeKCU1500_io_S_AXI_WVALID),
    .io_S_AXI_WREADY(AXI4LiteToRFBridgeKCU1500_io_S_AXI_WREADY),
    .io_S_AXI_RDATA(AXI4LiteToRFBridgeKCU1500_io_S_AXI_RDATA),
    .io_S_AXI_RRESP(AXI4LiteToRFBridgeKCU1500_io_S_AXI_RRESP),
    .io_S_AXI_RVALID(AXI4LiteToRFBridgeKCU1500_io_S_AXI_RVALID),
    .io_S_AXI_RREADY(AXI4LiteToRFBridgeKCU1500_io_S_AXI_RREADY),
    .io_S_AXI_BRESP(AXI4LiteToRFBridgeKCU1500_io_S_AXI_BRESP),
    .io_S_AXI_BVALID(AXI4LiteToRFBridgeKCU1500_io_S_AXI_BVALID),
    .io_S_AXI_BREADY(AXI4LiteToRFBridgeKCU1500_io_S_AXI_BREADY),
    .io_raddr(AXI4LiteToRFBridgeKCU1500_io_raddr),
    .io_wen(AXI4LiteToRFBridgeKCU1500_io_wen),
    .io_waddr(AXI4LiteToRFBridgeKCU1500_io_waddr),
    .io_wdata(AXI4LiteToRFBridgeKCU1500_io_wdata),
    .io_rdata(AXI4LiteToRFBridgeKCU1500_io_rdata)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge ( // @[FringeZynq.scala 130:27:@64382.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_io_in_cmd_bits_size),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_io_in_wdata_ready),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_io_in_rresp_ready),
    .io_in_rresp_valid(MAGToAXI4Bridge_io_in_rresp_valid),
    .io_in_rresp_bits_rdata_0(MAGToAXI4Bridge_io_in_rresp_bits_rdata_0),
    .io_in_rresp_bits_rdata_1(MAGToAXI4Bridge_io_in_rresp_bits_rdata_1),
    .io_in_rresp_bits_rdata_2(MAGToAXI4Bridge_io_in_rresp_bits_rdata_2),
    .io_in_rresp_bits_rdata_3(MAGToAXI4Bridge_io_in_rresp_bits_rdata_3),
    .io_in_rresp_bits_rdata_4(MAGToAXI4Bridge_io_in_rresp_bits_rdata_4),
    .io_in_rresp_bits_rdata_5(MAGToAXI4Bridge_io_in_rresp_bits_rdata_5),
    .io_in_rresp_bits_rdata_6(MAGToAXI4Bridge_io_in_rresp_bits_rdata_6),
    .io_in_rresp_bits_rdata_7(MAGToAXI4Bridge_io_in_rresp_bits_rdata_7),
    .io_in_rresp_bits_rdata_8(MAGToAXI4Bridge_io_in_rresp_bits_rdata_8),
    .io_in_rresp_bits_rdata_9(MAGToAXI4Bridge_io_in_rresp_bits_rdata_9),
    .io_in_rresp_bits_rdata_10(MAGToAXI4Bridge_io_in_rresp_bits_rdata_10),
    .io_in_rresp_bits_rdata_11(MAGToAXI4Bridge_io_in_rresp_bits_rdata_11),
    .io_in_rresp_bits_rdata_12(MAGToAXI4Bridge_io_in_rresp_bits_rdata_12),
    .io_in_rresp_bits_rdata_13(MAGToAXI4Bridge_io_in_rresp_bits_rdata_13),
    .io_in_rresp_bits_rdata_14(MAGToAXI4Bridge_io_in_rresp_bits_rdata_14),
    .io_in_rresp_bits_rdata_15(MAGToAXI4Bridge_io_in_rresp_bits_rdata_15),
    .io_in_rresp_bits_tag(MAGToAXI4Bridge_io_in_rresp_bits_tag),
    .io_in_wresp_ready(MAGToAXI4Bridge_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_io_M_AXI_AWLEN),
    .io_M_AXI_ARID(MAGToAXI4Bridge_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_io_M_AXI_ARREADY),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_io_M_AXI_WLAST),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_io_M_AXI_WREADY),
    .io_M_AXI_RID(MAGToAXI4Bridge_io_M_AXI_RID),
    .io_M_AXI_RDATA(MAGToAXI4Bridge_io_M_AXI_RDATA),
    .io_M_AXI_RVALID(MAGToAXI4Bridge_io_M_AXI_RVALID),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_io_M_AXI_BREADY)
  );
  assign io_S_AXI_AWREADY = AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWREADY; // @[FringeZynq.scala 79:28:@64204.4]
  assign io_S_AXI_ARREADY = AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARREADY; // @[FringeZynq.scala 79:28:@64200.4]
  assign io_S_AXI_WREADY = AXI4LiteToRFBridgeKCU1500_io_S_AXI_WREADY; // @[FringeZynq.scala 79:28:@64196.4]
  assign io_S_AXI_RDATA = AXI4LiteToRFBridgeKCU1500_io_S_AXI_RDATA; // @[FringeZynq.scala 79:28:@64195.4]
  assign io_S_AXI_RRESP = AXI4LiteToRFBridgeKCU1500_io_S_AXI_RRESP; // @[FringeZynq.scala 79:28:@64194.4]
  assign io_S_AXI_RVALID = AXI4LiteToRFBridgeKCU1500_io_S_AXI_RVALID; // @[FringeZynq.scala 79:28:@64193.4]
  assign io_S_AXI_BRESP = AXI4LiteToRFBridgeKCU1500_io_S_AXI_BRESP; // @[FringeZynq.scala 79:28:@64191.4]
  assign io_S_AXI_BVALID = AXI4LiteToRFBridgeKCU1500_io_S_AXI_BVALID; // @[FringeZynq.scala 79:28:@64190.4]
  assign io_M_AXI_0_AWID = MAGToAXI4Bridge_io_M_AXI_AWID; // @[FringeZynq.scala 132:10:@64537.4]
  assign io_M_AXI_0_AWADDR = MAGToAXI4Bridge_io_M_AXI_AWADDR; // @[FringeZynq.scala 132:10:@64535.4]
  assign io_M_AXI_0_AWLEN = MAGToAXI4Bridge_io_M_AXI_AWLEN; // @[FringeZynq.scala 132:10:@64534.4]
  assign io_M_AXI_0_ARID = MAGToAXI4Bridge_io_M_AXI_ARID; // @[FringeZynq.scala 132:10:@64525.4]
  assign io_M_AXI_0_ARADDR = MAGToAXI4Bridge_io_M_AXI_ARADDR; // @[FringeZynq.scala 132:10:@64523.4]
  assign io_M_AXI_0_ARLEN = MAGToAXI4Bridge_io_M_AXI_ARLEN; // @[FringeZynq.scala 132:10:@64522.4]
  assign io_M_AXI_0_ARVALID = MAGToAXI4Bridge_io_M_AXI_ARVALID; // @[FringeZynq.scala 132:10:@64515.4]
  assign io_M_AXI_0_WLAST = MAGToAXI4Bridge_io_M_AXI_WLAST; // @[FringeZynq.scala 132:10:@64511.4]
  assign io_M_AXI_0_RREADY = MAGToAXI4Bridge_io_M_AXI_RREADY; // @[FringeZynq.scala 132:10:@64502.4]
  assign io_M_AXI_0_BREADY = MAGToAXI4Bridge_io_M_AXI_BREADY; // @[FringeZynq.scala 132:10:@64497.4]
  assign io_enable = fringeCommon_io_enable; // @[FringeZynq.scala 114:13:@64216.4]
  assign io_reset = fringeCommon_io_reset; // @[FringeZynq.scala 118:12:@64220.4]
  assign io_argIns_0 = fringeCommon_io_argIns_0; // @[FringeZynq.scala 120:13:@64221.4]
  assign io_memStreams_loads_0_cmd_ready = fringeCommon_io_memStreams_loads_0_cmd_ready; // @[FringeZynq.scala 125:17:@64375.4]
  assign io_memStreams_loads_0_data_valid = fringeCommon_io_memStreams_loads_0_data_valid; // @[FringeZynq.scala 125:17:@64370.4]
  assign io_memStreams_loads_0_data_bits_rdata_0 = fringeCommon_io_memStreams_loads_0_data_bits_rdata_0; // @[FringeZynq.scala 125:17:@64369.4]
  assign io_heap_0_resp_valid = fringeCommon_io_heap_0_resp_valid; // @[FringeZynq.scala 126:11:@64378.4]
  assign io_heap_0_resp_bits_allocDealloc = fringeCommon_io_heap_0_resp_bits_allocDealloc; // @[FringeZynq.scala 126:11:@64377.4]
  assign io_heap_0_resp_bits_sizeAddr = fringeCommon_io_heap_0_resp_bits_sizeAddr; // @[FringeZynq.scala 126:11:@64376.4]
  assign fringeCommon_clock = clock; // @[:@63558.4]
  assign fringeCommon_reset = reset; // @[:@63559.4 FringeZynq.scala 81:24:@64209.4 FringeZynq.scala 116:22:@64219.4]
  assign fringeCommon_io_raddr = AXI4LiteToRFBridgeKCU1500_io_raddr; // @[FringeZynq.scala 82:27:@64210.4]
  assign fringeCommon_io_wen = AXI4LiteToRFBridgeKCU1500_io_wen; // @[FringeZynq.scala 83:27:@64211.4]
  assign fringeCommon_io_waddr = AXI4LiteToRFBridgeKCU1500_io_waddr; // @[FringeZynq.scala 84:27:@64212.4]
  assign fringeCommon_io_wdata = {{32'd0}, AXI4LiteToRFBridgeKCU1500_io_wdata}; // @[FringeZynq.scala 85:27:@64213.4]
  assign fringeCommon_io_done = io_done; // @[FringeZynq.scala 115:24:@64217.4]
  assign fringeCommon_io_argOuts_0_valid = io_argOuts_0_valid; // @[FringeZynq.scala 121:27:@64223.4]
  assign fringeCommon_io_argOuts_0_bits = io_argOuts_0_bits; // @[FringeZynq.scala 121:27:@64222.4]
  assign fringeCommon_io_argOuts_1_valid = io_argOuts_1_valid; // @[FringeZynq.scala 121:27:@64226.4]
  assign fringeCommon_io_argOuts_1_bits = io_argOuts_1_bits; // @[FringeZynq.scala 121:27:@64225.4]
  assign fringeCommon_io_argOuts_2_valid = io_argOuts_2_valid; // @[FringeZynq.scala 121:27:@64229.4]
  assign fringeCommon_io_argOuts_2_bits = io_argOuts_2_bits; // @[FringeZynq.scala 121:27:@64228.4]
  assign fringeCommon_io_argOuts_3_valid = io_argOuts_3_valid; // @[FringeZynq.scala 121:27:@64232.4]
  assign fringeCommon_io_argOuts_3_bits = io_argOuts_3_bits; // @[FringeZynq.scala 121:27:@64231.4]
  assign fringeCommon_io_argOuts_4_valid = io_argOuts_4_valid; // @[FringeZynq.scala 121:27:@64235.4]
  assign fringeCommon_io_argOuts_4_bits = io_argOuts_4_bits; // @[FringeZynq.scala 121:27:@64234.4]
  assign fringeCommon_io_argOuts_5_valid = io_argOuts_5_valid; // @[FringeZynq.scala 121:27:@64238.4]
  assign fringeCommon_io_argOuts_5_bits = io_argOuts_5_bits; // @[FringeZynq.scala 121:27:@64237.4]
  assign fringeCommon_io_argOuts_6_valid = io_argOuts_6_valid; // @[FringeZynq.scala 121:27:@64241.4]
  assign fringeCommon_io_argOuts_6_bits = io_argOuts_6_bits; // @[FringeZynq.scala 121:27:@64240.4]
  assign fringeCommon_io_argOuts_7_valid = io_argOuts_7_valid; // @[FringeZynq.scala 121:27:@64244.4]
  assign fringeCommon_io_argOuts_7_bits = io_argOuts_7_bits; // @[FringeZynq.scala 121:27:@64243.4]
  assign fringeCommon_io_argOuts_8_valid = io_argOuts_8_valid; // @[FringeZynq.scala 121:27:@64247.4]
  assign fringeCommon_io_argOuts_8_bits = io_argOuts_8_bits; // @[FringeZynq.scala 121:27:@64246.4]
  assign fringeCommon_io_argOuts_9_valid = io_argOuts_9_valid; // @[FringeZynq.scala 121:27:@64250.4]
  assign fringeCommon_io_argOuts_9_bits = io_argOuts_9_bits; // @[FringeZynq.scala 121:27:@64249.4]
  assign fringeCommon_io_argOuts_10_valid = io_argOuts_10_valid; // @[FringeZynq.scala 121:27:@64253.4]
  assign fringeCommon_io_argOuts_10_bits = io_argOuts_10_bits; // @[FringeZynq.scala 121:27:@64252.4]
  assign fringeCommon_io_argOuts_11_valid = io_argOuts_11_valid; // @[FringeZynq.scala 121:27:@64256.4]
  assign fringeCommon_io_argOuts_11_bits = io_argOuts_11_bits; // @[FringeZynq.scala 121:27:@64255.4]
  assign fringeCommon_io_argOuts_12_valid = io_argOuts_12_valid; // @[FringeZynq.scala 121:27:@64259.4]
  assign fringeCommon_io_argOuts_12_bits = io_argOuts_12_bits; // @[FringeZynq.scala 121:27:@64258.4]
  assign fringeCommon_io_argOuts_13_valid = io_argOuts_13_valid; // @[FringeZynq.scala 121:27:@64262.4]
  assign fringeCommon_io_argOuts_13_bits = io_argOuts_13_bits; // @[FringeZynq.scala 121:27:@64261.4]
  assign fringeCommon_io_argOuts_14_valid = io_argOuts_14_valid; // @[FringeZynq.scala 121:27:@64265.4]
  assign fringeCommon_io_argOuts_14_bits = io_argOuts_14_bits; // @[FringeZynq.scala 121:27:@64264.4]
  assign fringeCommon_io_argOuts_15_valid = io_argOuts_15_valid; // @[FringeZynq.scala 121:27:@64268.4]
  assign fringeCommon_io_argOuts_15_bits = io_argOuts_15_bits; // @[FringeZynq.scala 121:27:@64267.4]
  assign fringeCommon_io_memStreams_loads_0_cmd_valid = io_memStreams_loads_0_cmd_valid; // @[FringeZynq.scala 125:17:@64374.4]
  assign fringeCommon_io_memStreams_loads_0_cmd_bits_addr = io_memStreams_loads_0_cmd_bits_addr; // @[FringeZynq.scala 125:17:@64373.4]
  assign fringeCommon_io_memStreams_loads_0_cmd_bits_size = io_memStreams_loads_0_cmd_bits_size; // @[FringeZynq.scala 125:17:@64372.4]
  assign fringeCommon_io_memStreams_loads_0_data_ready = io_memStreams_loads_0_data_ready; // @[FringeZynq.scala 125:17:@64371.4]
  assign fringeCommon_io_memStreams_stores_0_cmd_valid = io_memStreams_stores_0_cmd_valid; // @[FringeZynq.scala 125:17:@64367.4]
  assign fringeCommon_io_memStreams_stores_0_cmd_bits_addr = io_memStreams_stores_0_cmd_bits_addr; // @[FringeZynq.scala 125:17:@64366.4]
  assign fringeCommon_io_memStreams_stores_0_cmd_bits_size = io_memStreams_stores_0_cmd_bits_size; // @[FringeZynq.scala 125:17:@64365.4]
  assign fringeCommon_io_memStreams_stores_0_data_valid = io_memStreams_stores_0_data_valid; // @[FringeZynq.scala 125:17:@64363.4]
  assign fringeCommon_io_memStreams_stores_0_data_bits_wdata_0 = io_memStreams_stores_0_data_bits_wdata_0; // @[FringeZynq.scala 125:17:@64347.4]
  assign fringeCommon_io_memStreams_stores_0_data_bits_wstrb = io_memStreams_stores_0_data_bits_wstrb; // @[FringeZynq.scala 125:17:@64346.4]
  assign fringeCommon_io_dram_0_cmd_ready = MAGToAXI4Bridge_io_in_cmd_ready; // @[FringeZynq.scala 131:21:@64496.4]
  assign fringeCommon_io_dram_0_wdata_ready = MAGToAXI4Bridge_io_in_wdata_ready; // @[FringeZynq.scala 131:21:@64489.4]
  assign fringeCommon_io_dram_0_rresp_valid = MAGToAXI4Bridge_io_in_rresp_valid; // @[FringeZynq.scala 131:21:@64405.4]
  assign fringeCommon_io_dram_0_rresp_bits_rdata_0 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_0; // @[FringeZynq.scala 131:21:@64389.4]
  assign fringeCommon_io_dram_0_rresp_bits_rdata_1 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_1; // @[FringeZynq.scala 131:21:@64390.4]
  assign fringeCommon_io_dram_0_rresp_bits_rdata_2 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_2; // @[FringeZynq.scala 131:21:@64391.4]
  assign fringeCommon_io_dram_0_rresp_bits_rdata_3 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_3; // @[FringeZynq.scala 131:21:@64392.4]
  assign fringeCommon_io_dram_0_rresp_bits_rdata_4 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_4; // @[FringeZynq.scala 131:21:@64393.4]
  assign fringeCommon_io_dram_0_rresp_bits_rdata_5 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_5; // @[FringeZynq.scala 131:21:@64394.4]
  assign fringeCommon_io_dram_0_rresp_bits_rdata_6 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_6; // @[FringeZynq.scala 131:21:@64395.4]
  assign fringeCommon_io_dram_0_rresp_bits_rdata_7 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_7; // @[FringeZynq.scala 131:21:@64396.4]
  assign fringeCommon_io_dram_0_rresp_bits_rdata_8 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_8; // @[FringeZynq.scala 131:21:@64397.4]
  assign fringeCommon_io_dram_0_rresp_bits_rdata_9 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_9; // @[FringeZynq.scala 131:21:@64398.4]
  assign fringeCommon_io_dram_0_rresp_bits_rdata_10 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_10; // @[FringeZynq.scala 131:21:@64399.4]
  assign fringeCommon_io_dram_0_rresp_bits_rdata_11 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_11; // @[FringeZynq.scala 131:21:@64400.4]
  assign fringeCommon_io_dram_0_rresp_bits_rdata_12 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_12; // @[FringeZynq.scala 131:21:@64401.4]
  assign fringeCommon_io_dram_0_rresp_bits_rdata_13 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_13; // @[FringeZynq.scala 131:21:@64402.4]
  assign fringeCommon_io_dram_0_rresp_bits_rdata_14 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_14; // @[FringeZynq.scala 131:21:@64403.4]
  assign fringeCommon_io_dram_0_rresp_bits_rdata_15 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_15; // @[FringeZynq.scala 131:21:@64404.4]
  assign fringeCommon_io_dram_0_rresp_bits_tag = MAGToAXI4Bridge_io_in_rresp_bits_tag; // @[FringeZynq.scala 131:21:@64388.4]
  assign fringeCommon_io_dram_0_wresp_valid = MAGToAXI4Bridge_io_in_wresp_valid; // @[FringeZynq.scala 131:21:@64386.4]
  assign fringeCommon_io_dram_0_wresp_bits_tag = MAGToAXI4Bridge_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:21:@64385.4]
  assign fringeCommon_io_heap_0_req_valid = io_heap_0_req_valid; // @[FringeZynq.scala 126:11:@64381.4]
  assign fringeCommon_io_heap_0_req_bits_allocDealloc = io_heap_0_req_bits_allocDealloc; // @[FringeZynq.scala 126:11:@64380.4]
  assign fringeCommon_io_heap_0_req_bits_sizeAddr = io_heap_0_req_bits_sizeAddr; // @[FringeZynq.scala 126:11:@64379.4]
  assign AXI4LiteToRFBridgeKCU1500_clock = clock; // @[:@64187.4]
  assign AXI4LiteToRFBridgeKCU1500_reset = reset; // @[:@64188.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[FringeZynq.scala 79:28:@64207.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[FringeZynq.scala 79:28:@64206.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[FringeZynq.scala 79:28:@64205.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[FringeZynq.scala 79:28:@64203.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[FringeZynq.scala 79:28:@64202.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[FringeZynq.scala 79:28:@64201.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_WDATA = io_S_AXI_WDATA; // @[FringeZynq.scala 79:28:@64199.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[FringeZynq.scala 79:28:@64198.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_WVALID = io_S_AXI_WVALID; // @[FringeZynq.scala 79:28:@64197.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_RREADY = io_S_AXI_RREADY; // @[FringeZynq.scala 79:28:@64192.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_BREADY = io_S_AXI_BREADY; // @[FringeZynq.scala 79:28:@64189.4]
  assign AXI4LiteToRFBridgeKCU1500_io_rdata = fringeCommon_io_rdata[31:0]; // @[FringeZynq.scala 86:28:@64214.4]
  assign MAGToAXI4Bridge_io_in_cmd_valid = fringeCommon_io_dram_0_cmd_valid; // @[FringeZynq.scala 131:21:@64495.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_addr = fringeCommon_io_dram_0_cmd_bits_addr; // @[FringeZynq.scala 131:21:@64494.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_size = fringeCommon_io_dram_0_cmd_bits_size; // @[FringeZynq.scala 131:21:@64493.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_tag = fringeCommon_io_dram_0_cmd_bits_tag; // @[FringeZynq.scala 131:21:@64490.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wlast = fringeCommon_io_dram_0_wdata_bits_wlast; // @[FringeZynq.scala 131:21:@64407.4]
  assign MAGToAXI4Bridge_io_in_rresp_ready = fringeCommon_io_dram_0_rresp_ready; // @[FringeZynq.scala 131:21:@64406.4]
  assign MAGToAXI4Bridge_io_in_wresp_ready = fringeCommon_io_dram_0_wresp_ready; // @[FringeZynq.scala 131:21:@64387.4]
  assign MAGToAXI4Bridge_io_M_AXI_ARREADY = io_M_AXI_0_ARREADY; // @[FringeZynq.scala 132:10:@64514.4]
  assign MAGToAXI4Bridge_io_M_AXI_WREADY = io_M_AXI_0_WREADY; // @[FringeZynq.scala 132:10:@64509.4]
  assign MAGToAXI4Bridge_io_M_AXI_RID = io_M_AXI_0_RID; // @[FringeZynq.scala 132:10:@64508.4]
  assign MAGToAXI4Bridge_io_M_AXI_RDATA = io_M_AXI_0_RDATA; // @[FringeZynq.scala 132:10:@64506.4]
  assign MAGToAXI4Bridge_io_M_AXI_RVALID = io_M_AXI_0_RVALID; // @[FringeZynq.scala 132:10:@64503.4]
  assign MAGToAXI4Bridge_io_M_AXI_BID = io_M_AXI_0_BID; // @[FringeZynq.scala 132:10:@64501.4]
  assign MAGToAXI4Bridge_io_M_AXI_BVALID = io_M_AXI_0_BVALID; // @[FringeZynq.scala 132:10:@64498.4]
endmodule
module Top( // @[:@64539.2]
  input          clock, // @[:@64540.4]
  input          reset, // @[:@64541.4]
  input          io_raddr, // @[:@64542.4]
  input          io_wen, // @[:@64542.4]
  input          io_waddr, // @[:@64542.4]
  input          io_wdata, // @[:@64542.4]
  output         io_rdata, // @[:@64542.4]
  input  [31:0]  io_S_AXI_AWADDR, // @[:@64542.4]
  input  [2:0]   io_S_AXI_AWPROT, // @[:@64542.4]
  input          io_S_AXI_AWVALID, // @[:@64542.4]
  output         io_S_AXI_AWREADY, // @[:@64542.4]
  input  [31:0]  io_S_AXI_ARADDR, // @[:@64542.4]
  input  [2:0]   io_S_AXI_ARPROT, // @[:@64542.4]
  input          io_S_AXI_ARVALID, // @[:@64542.4]
  output         io_S_AXI_ARREADY, // @[:@64542.4]
  input  [31:0]  io_S_AXI_WDATA, // @[:@64542.4]
  input  [3:0]   io_S_AXI_WSTRB, // @[:@64542.4]
  input          io_S_AXI_WVALID, // @[:@64542.4]
  output         io_S_AXI_WREADY, // @[:@64542.4]
  output [31:0]  io_S_AXI_RDATA, // @[:@64542.4]
  output [1:0]   io_S_AXI_RRESP, // @[:@64542.4]
  output         io_S_AXI_RVALID, // @[:@64542.4]
  input          io_S_AXI_RREADY, // @[:@64542.4]
  output [1:0]   io_S_AXI_BRESP, // @[:@64542.4]
  output         io_S_AXI_BVALID, // @[:@64542.4]
  input          io_S_AXI_BREADY, // @[:@64542.4]
  output [3:0]   io_M_AXI_0_AWID, // @[:@64542.4]
  output [3:0]   io_M_AXI_0_AWUSER, // @[:@64542.4]
  output [31:0]  io_M_AXI_0_AWADDR, // @[:@64542.4]
  output [7:0]   io_M_AXI_0_AWLEN, // @[:@64542.4]
  output [2:0]   io_M_AXI_0_AWSIZE, // @[:@64542.4]
  output [1:0]   io_M_AXI_0_AWBURST, // @[:@64542.4]
  output         io_M_AXI_0_AWLOCK, // @[:@64542.4]
  output [3:0]   io_M_AXI_0_AWCACHE, // @[:@64542.4]
  output [2:0]   io_M_AXI_0_AWPROT, // @[:@64542.4]
  output [3:0]   io_M_AXI_0_AWQOS, // @[:@64542.4]
  output         io_M_AXI_0_AWVALID, // @[:@64542.4]
  input          io_M_AXI_0_AWREADY, // @[:@64542.4]
  output [3:0]   io_M_AXI_0_ARID, // @[:@64542.4]
  output [3:0]   io_M_AXI_0_ARUSER, // @[:@64542.4]
  output [31:0]  io_M_AXI_0_ARADDR, // @[:@64542.4]
  output [7:0]   io_M_AXI_0_ARLEN, // @[:@64542.4]
  output [2:0]   io_M_AXI_0_ARSIZE, // @[:@64542.4]
  output [1:0]   io_M_AXI_0_ARBURST, // @[:@64542.4]
  output         io_M_AXI_0_ARLOCK, // @[:@64542.4]
  output [3:0]   io_M_AXI_0_ARCACHE, // @[:@64542.4]
  output [2:0]   io_M_AXI_0_ARPROT, // @[:@64542.4]
  output [3:0]   io_M_AXI_0_ARQOS, // @[:@64542.4]
  output         io_M_AXI_0_ARVALID, // @[:@64542.4]
  input          io_M_AXI_0_ARREADY, // @[:@64542.4]
  output [511:0] io_M_AXI_0_WDATA, // @[:@64542.4]
  output [63:0]  io_M_AXI_0_WSTRB, // @[:@64542.4]
  output         io_M_AXI_0_WLAST, // @[:@64542.4]
  output         io_M_AXI_0_WVALID, // @[:@64542.4]
  input          io_M_AXI_0_WREADY, // @[:@64542.4]
  input  [3:0]   io_M_AXI_0_RID, // @[:@64542.4]
  input  [31:0]  io_M_AXI_0_RUSER, // @[:@64542.4]
  input  [511:0] io_M_AXI_0_RDATA, // @[:@64542.4]
  input  [1:0]   io_M_AXI_0_RRESP, // @[:@64542.4]
  input          io_M_AXI_0_RLAST, // @[:@64542.4]
  input          io_M_AXI_0_RVALID, // @[:@64542.4]
  output         io_M_AXI_0_RREADY, // @[:@64542.4]
  input  [3:0]   io_M_AXI_0_BID, // @[:@64542.4]
  input  [3:0]   io_M_AXI_0_BUSER, // @[:@64542.4]
  input  [1:0]   io_M_AXI_0_BRESP, // @[:@64542.4]
  input          io_M_AXI_0_BVALID, // @[:@64542.4]
  output         io_M_AXI_0_BREADY // @[:@64542.4]
);
  wire  accel_clock; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_reset; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_enable; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_done; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_reset; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_memStreams_loads_0_cmd_ready; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_memStreams_loads_0_cmd_valid; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_memStreams_loads_0_cmd_bits_addr; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_loads_0_cmd_bits_size; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_memStreams_loads_0_data_ready; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_memStreams_loads_0_data_valid; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_0; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_memStreams_stores_0_cmd_ready; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_memStreams_stores_0_cmd_valid; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_memStreams_stores_0_cmd_bits_addr; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_stores_0_cmd_bits_size; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_memStreams_stores_0_data_ready; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_memStreams_stores_0_data_valid; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_0; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_1; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_2; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_3; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_4; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_5; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_6; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_7; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_8; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_9; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_10; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_11; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_12; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_13; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_14; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_15; // @[Instantiator.scala 68:38:@64544.4]
  wire [15:0] accel_io_memStreams_stores_0_data_bits_wstrb; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_memStreams_stores_0_wresp_ready; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_memStreams_stores_0_wresp_valid; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_memStreams_stores_0_wresp_bits; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_memStreams_gathers_0_cmd_ready; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_memStreams_gathers_0_cmd_valid; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_0; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_1; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_2; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_3; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_4; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_5; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_6; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_7; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_8; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_9; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_10; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_11; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_12; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_13; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_14; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_15; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_memStreams_gathers_0_data_ready; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_memStreams_gathers_0_data_valid; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_0; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_1; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_2; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_3; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_4; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_5; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_6; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_7; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_8; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_9; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_10; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_11; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_12; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_13; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_14; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_15; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_memStreams_scatters_0_cmd_ready; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_memStreams_scatters_0_cmd_valid; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_0; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_1; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_2; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_3; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_4; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_5; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_6; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_7; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_8; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_9; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_10; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_11; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_12; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_13; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_14; // @[Instantiator.scala 68:38:@64544.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_15; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_memStreams_scatters_0_wresp_ready; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_memStreams_scatters_0_wresp_valid; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_memStreams_scatters_0_wresp_bits; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_heap_0_req_valid; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_heap_0_req_bits_allocDealloc; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_heap_0_req_bits_sizeAddr; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_heap_0_resp_valid; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_heap_0_resp_bits_allocDealloc; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_heap_0_resp_bits_sizeAddr; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_argIns_0; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_argOuts_0_port_ready; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_argOuts_0_port_valid; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_argOuts_0_port_bits; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_argOuts_0_echo; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_argOuts_1_port_ready; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_argOuts_1_port_valid; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_argOuts_1_port_bits; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_argOuts_1_echo; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_argOuts_2_port_ready; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_argOuts_2_port_valid; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_argOuts_2_port_bits; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_argOuts_2_echo; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_argOuts_3_port_ready; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_argOuts_3_port_valid; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_argOuts_3_port_bits; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_argOuts_3_echo; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_argOuts_4_port_ready; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_argOuts_4_port_valid; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_argOuts_4_port_bits; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_argOuts_4_echo; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_argOuts_5_port_ready; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_argOuts_5_port_valid; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_argOuts_5_port_bits; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_argOuts_5_echo; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_argOuts_6_port_ready; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_argOuts_6_port_valid; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_argOuts_6_port_bits; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_argOuts_6_echo; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_argOuts_7_port_ready; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_argOuts_7_port_valid; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_argOuts_7_port_bits; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_argOuts_7_echo; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_argOuts_8_port_ready; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_argOuts_8_port_valid; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_argOuts_8_port_bits; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_argOuts_8_echo; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_argOuts_9_port_ready; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_argOuts_9_port_valid; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_argOuts_9_port_bits; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_argOuts_9_echo; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_argOuts_10_port_ready; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_argOuts_10_port_valid; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_argOuts_10_port_bits; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_argOuts_10_echo; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_argOuts_11_port_ready; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_argOuts_11_port_valid; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_argOuts_11_port_bits; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_argOuts_11_echo; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_argOuts_12_port_ready; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_argOuts_12_port_valid; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_argOuts_12_port_bits; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_argOuts_12_echo; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_argOuts_13_port_ready; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_argOuts_13_port_valid; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_argOuts_13_port_bits; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_argOuts_13_echo; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_argOuts_14_port_ready; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_argOuts_14_port_valid; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_argOuts_14_port_bits; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_argOuts_14_echo; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_argOuts_15_port_ready; // @[Instantiator.scala 68:38:@64544.4]
  wire  accel_io_argOuts_15_port_valid; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_argOuts_15_port_bits; // @[Instantiator.scala 68:38:@64544.4]
  wire [63:0] accel_io_argOuts_15_echo; // @[Instantiator.scala 68:38:@64544.4]
  wire  FringeZynq_clock; // @[KCU1500.scala 21:24:@64727.4]
  wire  FringeZynq_reset; // @[KCU1500.scala 21:24:@64727.4]
  wire [31:0] FringeZynq_io_S_AXI_AWADDR; // @[KCU1500.scala 21:24:@64727.4]
  wire [2:0] FringeZynq_io_S_AXI_AWPROT; // @[KCU1500.scala 21:24:@64727.4]
  wire  FringeZynq_io_S_AXI_AWVALID; // @[KCU1500.scala 21:24:@64727.4]
  wire  FringeZynq_io_S_AXI_AWREADY; // @[KCU1500.scala 21:24:@64727.4]
  wire [31:0] FringeZynq_io_S_AXI_ARADDR; // @[KCU1500.scala 21:24:@64727.4]
  wire [2:0] FringeZynq_io_S_AXI_ARPROT; // @[KCU1500.scala 21:24:@64727.4]
  wire  FringeZynq_io_S_AXI_ARVALID; // @[KCU1500.scala 21:24:@64727.4]
  wire  FringeZynq_io_S_AXI_ARREADY; // @[KCU1500.scala 21:24:@64727.4]
  wire [31:0] FringeZynq_io_S_AXI_WDATA; // @[KCU1500.scala 21:24:@64727.4]
  wire [3:0] FringeZynq_io_S_AXI_WSTRB; // @[KCU1500.scala 21:24:@64727.4]
  wire  FringeZynq_io_S_AXI_WVALID; // @[KCU1500.scala 21:24:@64727.4]
  wire  FringeZynq_io_S_AXI_WREADY; // @[KCU1500.scala 21:24:@64727.4]
  wire [31:0] FringeZynq_io_S_AXI_RDATA; // @[KCU1500.scala 21:24:@64727.4]
  wire [1:0] FringeZynq_io_S_AXI_RRESP; // @[KCU1500.scala 21:24:@64727.4]
  wire  FringeZynq_io_S_AXI_RVALID; // @[KCU1500.scala 21:24:@64727.4]
  wire  FringeZynq_io_S_AXI_RREADY; // @[KCU1500.scala 21:24:@64727.4]
  wire [1:0] FringeZynq_io_S_AXI_BRESP; // @[KCU1500.scala 21:24:@64727.4]
  wire  FringeZynq_io_S_AXI_BVALID; // @[KCU1500.scala 21:24:@64727.4]
  wire  FringeZynq_io_S_AXI_BREADY; // @[KCU1500.scala 21:24:@64727.4]
  wire [3:0] FringeZynq_io_M_AXI_0_AWID; // @[KCU1500.scala 21:24:@64727.4]
  wire [31:0] FringeZynq_io_M_AXI_0_AWADDR; // @[KCU1500.scala 21:24:@64727.4]
  wire [7:0] FringeZynq_io_M_AXI_0_AWLEN; // @[KCU1500.scala 21:24:@64727.4]
  wire [3:0] FringeZynq_io_M_AXI_0_ARID; // @[KCU1500.scala 21:24:@64727.4]
  wire [31:0] FringeZynq_io_M_AXI_0_ARADDR; // @[KCU1500.scala 21:24:@64727.4]
  wire [7:0] FringeZynq_io_M_AXI_0_ARLEN; // @[KCU1500.scala 21:24:@64727.4]
  wire  FringeZynq_io_M_AXI_0_ARVALID; // @[KCU1500.scala 21:24:@64727.4]
  wire  FringeZynq_io_M_AXI_0_ARREADY; // @[KCU1500.scala 21:24:@64727.4]
  wire  FringeZynq_io_M_AXI_0_WLAST; // @[KCU1500.scala 21:24:@64727.4]
  wire  FringeZynq_io_M_AXI_0_WREADY; // @[KCU1500.scala 21:24:@64727.4]
  wire [3:0] FringeZynq_io_M_AXI_0_RID; // @[KCU1500.scala 21:24:@64727.4]
  wire [511:0] FringeZynq_io_M_AXI_0_RDATA; // @[KCU1500.scala 21:24:@64727.4]
  wire  FringeZynq_io_M_AXI_0_RVALID; // @[KCU1500.scala 21:24:@64727.4]
  wire  FringeZynq_io_M_AXI_0_RREADY; // @[KCU1500.scala 21:24:@64727.4]
  wire [3:0] FringeZynq_io_M_AXI_0_BID; // @[KCU1500.scala 21:24:@64727.4]
  wire  FringeZynq_io_M_AXI_0_BVALID; // @[KCU1500.scala 21:24:@64727.4]
  wire  FringeZynq_io_M_AXI_0_BREADY; // @[KCU1500.scala 21:24:@64727.4]
  wire  FringeZynq_io_enable; // @[KCU1500.scala 21:24:@64727.4]
  wire  FringeZynq_io_done; // @[KCU1500.scala 21:24:@64727.4]
  wire  FringeZynq_io_reset; // @[KCU1500.scala 21:24:@64727.4]
  wire [63:0] FringeZynq_io_argIns_0; // @[KCU1500.scala 21:24:@64727.4]
  wire  FringeZynq_io_argOuts_0_valid; // @[KCU1500.scala 21:24:@64727.4]
  wire [63:0] FringeZynq_io_argOuts_0_bits; // @[KCU1500.scala 21:24:@64727.4]
  wire  FringeZynq_io_argOuts_1_valid; // @[KCU1500.scala 21:24:@64727.4]
  wire [63:0] FringeZynq_io_argOuts_1_bits; // @[KCU1500.scala 21:24:@64727.4]
  wire  FringeZynq_io_argOuts_2_valid; // @[KCU1500.scala 21:24:@64727.4]
  wire [63:0] FringeZynq_io_argOuts_2_bits; // @[KCU1500.scala 21:24:@64727.4]
  wire  FringeZynq_io_argOuts_3_valid; // @[KCU1500.scala 21:24:@64727.4]
  wire [63:0] FringeZynq_io_argOuts_3_bits; // @[KCU1500.scala 21:24:@64727.4]
  wire  FringeZynq_io_argOuts_4_valid; // @[KCU1500.scala 21:24:@64727.4]
  wire [63:0] FringeZynq_io_argOuts_4_bits; // @[KCU1500.scala 21:24:@64727.4]
  wire  FringeZynq_io_argOuts_5_valid; // @[KCU1500.scala 21:24:@64727.4]
  wire [63:0] FringeZynq_io_argOuts_5_bits; // @[KCU1500.scala 21:24:@64727.4]
  wire  FringeZynq_io_argOuts_6_valid; // @[KCU1500.scala 21:24:@64727.4]
  wire [63:0] FringeZynq_io_argOuts_6_bits; // @[KCU1500.scala 21:24:@64727.4]
  wire  FringeZynq_io_argOuts_7_valid; // @[KCU1500.scala 21:24:@64727.4]
  wire [63:0] FringeZynq_io_argOuts_7_bits; // @[KCU1500.scala 21:24:@64727.4]
  wire  FringeZynq_io_argOuts_8_valid; // @[KCU1500.scala 21:24:@64727.4]
  wire [63:0] FringeZynq_io_argOuts_8_bits; // @[KCU1500.scala 21:24:@64727.4]
  wire  FringeZynq_io_argOuts_9_valid; // @[KCU1500.scala 21:24:@64727.4]
  wire [63:0] FringeZynq_io_argOuts_9_bits; // @[KCU1500.scala 21:24:@64727.4]
  wire  FringeZynq_io_argOuts_10_valid; // @[KCU1500.scala 21:24:@64727.4]
  wire [63:0] FringeZynq_io_argOuts_10_bits; // @[KCU1500.scala 21:24:@64727.4]
  wire  FringeZynq_io_argOuts_11_valid; // @[KCU1500.scala 21:24:@64727.4]
  wire [63:0] FringeZynq_io_argOuts_11_bits; // @[KCU1500.scala 21:24:@64727.4]
  wire  FringeZynq_io_argOuts_12_valid; // @[KCU1500.scala 21:24:@64727.4]
  wire [63:0] FringeZynq_io_argOuts_12_bits; // @[KCU1500.scala 21:24:@64727.4]
  wire  FringeZynq_io_argOuts_13_valid; // @[KCU1500.scala 21:24:@64727.4]
  wire [63:0] FringeZynq_io_argOuts_13_bits; // @[KCU1500.scala 21:24:@64727.4]
  wire  FringeZynq_io_argOuts_14_valid; // @[KCU1500.scala 21:24:@64727.4]
  wire [63:0] FringeZynq_io_argOuts_14_bits; // @[KCU1500.scala 21:24:@64727.4]
  wire  FringeZynq_io_argOuts_15_valid; // @[KCU1500.scala 21:24:@64727.4]
  wire [63:0] FringeZynq_io_argOuts_15_bits; // @[KCU1500.scala 21:24:@64727.4]
  wire  FringeZynq_io_memStreams_loads_0_cmd_ready; // @[KCU1500.scala 21:24:@64727.4]
  wire  FringeZynq_io_memStreams_loads_0_cmd_valid; // @[KCU1500.scala 21:24:@64727.4]
  wire [63:0] FringeZynq_io_memStreams_loads_0_cmd_bits_addr; // @[KCU1500.scala 21:24:@64727.4]
  wire [31:0] FringeZynq_io_memStreams_loads_0_cmd_bits_size; // @[KCU1500.scala 21:24:@64727.4]
  wire  FringeZynq_io_memStreams_loads_0_data_ready; // @[KCU1500.scala 21:24:@64727.4]
  wire  FringeZynq_io_memStreams_loads_0_data_valid; // @[KCU1500.scala 21:24:@64727.4]
  wire [31:0] FringeZynq_io_memStreams_loads_0_data_bits_rdata_0; // @[KCU1500.scala 21:24:@64727.4]
  wire  FringeZynq_io_memStreams_stores_0_cmd_valid; // @[KCU1500.scala 21:24:@64727.4]
  wire [63:0] FringeZynq_io_memStreams_stores_0_cmd_bits_addr; // @[KCU1500.scala 21:24:@64727.4]
  wire [31:0] FringeZynq_io_memStreams_stores_0_cmd_bits_size; // @[KCU1500.scala 21:24:@64727.4]
  wire  FringeZynq_io_memStreams_stores_0_data_valid; // @[KCU1500.scala 21:24:@64727.4]
  wire [31:0] FringeZynq_io_memStreams_stores_0_data_bits_wdata_0; // @[KCU1500.scala 21:24:@64727.4]
  wire [15:0] FringeZynq_io_memStreams_stores_0_data_bits_wstrb; // @[KCU1500.scala 21:24:@64727.4]
  wire  FringeZynq_io_heap_0_req_valid; // @[KCU1500.scala 21:24:@64727.4]
  wire  FringeZynq_io_heap_0_req_bits_allocDealloc; // @[KCU1500.scala 21:24:@64727.4]
  wire [63:0] FringeZynq_io_heap_0_req_bits_sizeAddr; // @[KCU1500.scala 21:24:@64727.4]
  wire  FringeZynq_io_heap_0_resp_valid; // @[KCU1500.scala 21:24:@64727.4]
  wire  FringeZynq_io_heap_0_resp_bits_allocDealloc; // @[KCU1500.scala 21:24:@64727.4]
  wire [63:0] FringeZynq_io_heap_0_resp_bits_sizeAddr; // @[KCU1500.scala 21:24:@64727.4]
  AccelTop accel ( // @[Instantiator.scala 68:38:@64544.4]
    .clock(accel_clock),
    .reset(accel_reset),
    .io_enable(accel_io_enable),
    .io_done(accel_io_done),
    .io_reset(accel_io_reset),
    .io_memStreams_loads_0_cmd_ready(accel_io_memStreams_loads_0_cmd_ready),
    .io_memStreams_loads_0_cmd_valid(accel_io_memStreams_loads_0_cmd_valid),
    .io_memStreams_loads_0_cmd_bits_addr(accel_io_memStreams_loads_0_cmd_bits_addr),
    .io_memStreams_loads_0_cmd_bits_size(accel_io_memStreams_loads_0_cmd_bits_size),
    .io_memStreams_loads_0_data_ready(accel_io_memStreams_loads_0_data_ready),
    .io_memStreams_loads_0_data_valid(accel_io_memStreams_loads_0_data_valid),
    .io_memStreams_loads_0_data_bits_rdata_0(accel_io_memStreams_loads_0_data_bits_rdata_0),
    .io_memStreams_stores_0_cmd_ready(accel_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(accel_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(accel_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(accel_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(accel_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(accel_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(accel_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wdata_1(accel_io_memStreams_stores_0_data_bits_wdata_1),
    .io_memStreams_stores_0_data_bits_wdata_2(accel_io_memStreams_stores_0_data_bits_wdata_2),
    .io_memStreams_stores_0_data_bits_wdata_3(accel_io_memStreams_stores_0_data_bits_wdata_3),
    .io_memStreams_stores_0_data_bits_wdata_4(accel_io_memStreams_stores_0_data_bits_wdata_4),
    .io_memStreams_stores_0_data_bits_wdata_5(accel_io_memStreams_stores_0_data_bits_wdata_5),
    .io_memStreams_stores_0_data_bits_wdata_6(accel_io_memStreams_stores_0_data_bits_wdata_6),
    .io_memStreams_stores_0_data_bits_wdata_7(accel_io_memStreams_stores_0_data_bits_wdata_7),
    .io_memStreams_stores_0_data_bits_wdata_8(accel_io_memStreams_stores_0_data_bits_wdata_8),
    .io_memStreams_stores_0_data_bits_wdata_9(accel_io_memStreams_stores_0_data_bits_wdata_9),
    .io_memStreams_stores_0_data_bits_wdata_10(accel_io_memStreams_stores_0_data_bits_wdata_10),
    .io_memStreams_stores_0_data_bits_wdata_11(accel_io_memStreams_stores_0_data_bits_wdata_11),
    .io_memStreams_stores_0_data_bits_wdata_12(accel_io_memStreams_stores_0_data_bits_wdata_12),
    .io_memStreams_stores_0_data_bits_wdata_13(accel_io_memStreams_stores_0_data_bits_wdata_13),
    .io_memStreams_stores_0_data_bits_wdata_14(accel_io_memStreams_stores_0_data_bits_wdata_14),
    .io_memStreams_stores_0_data_bits_wdata_15(accel_io_memStreams_stores_0_data_bits_wdata_15),
    .io_memStreams_stores_0_data_bits_wstrb(accel_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(accel_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(accel_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(accel_io_memStreams_stores_0_wresp_bits),
    .io_memStreams_gathers_0_cmd_ready(accel_io_memStreams_gathers_0_cmd_ready),
    .io_memStreams_gathers_0_cmd_valid(accel_io_memStreams_gathers_0_cmd_valid),
    .io_memStreams_gathers_0_cmd_bits_addr_0(accel_io_memStreams_gathers_0_cmd_bits_addr_0),
    .io_memStreams_gathers_0_cmd_bits_addr_1(accel_io_memStreams_gathers_0_cmd_bits_addr_1),
    .io_memStreams_gathers_0_cmd_bits_addr_2(accel_io_memStreams_gathers_0_cmd_bits_addr_2),
    .io_memStreams_gathers_0_cmd_bits_addr_3(accel_io_memStreams_gathers_0_cmd_bits_addr_3),
    .io_memStreams_gathers_0_cmd_bits_addr_4(accel_io_memStreams_gathers_0_cmd_bits_addr_4),
    .io_memStreams_gathers_0_cmd_bits_addr_5(accel_io_memStreams_gathers_0_cmd_bits_addr_5),
    .io_memStreams_gathers_0_cmd_bits_addr_6(accel_io_memStreams_gathers_0_cmd_bits_addr_6),
    .io_memStreams_gathers_0_cmd_bits_addr_7(accel_io_memStreams_gathers_0_cmd_bits_addr_7),
    .io_memStreams_gathers_0_cmd_bits_addr_8(accel_io_memStreams_gathers_0_cmd_bits_addr_8),
    .io_memStreams_gathers_0_cmd_bits_addr_9(accel_io_memStreams_gathers_0_cmd_bits_addr_9),
    .io_memStreams_gathers_0_cmd_bits_addr_10(accel_io_memStreams_gathers_0_cmd_bits_addr_10),
    .io_memStreams_gathers_0_cmd_bits_addr_11(accel_io_memStreams_gathers_0_cmd_bits_addr_11),
    .io_memStreams_gathers_0_cmd_bits_addr_12(accel_io_memStreams_gathers_0_cmd_bits_addr_12),
    .io_memStreams_gathers_0_cmd_bits_addr_13(accel_io_memStreams_gathers_0_cmd_bits_addr_13),
    .io_memStreams_gathers_0_cmd_bits_addr_14(accel_io_memStreams_gathers_0_cmd_bits_addr_14),
    .io_memStreams_gathers_0_cmd_bits_addr_15(accel_io_memStreams_gathers_0_cmd_bits_addr_15),
    .io_memStreams_gathers_0_data_ready(accel_io_memStreams_gathers_0_data_ready),
    .io_memStreams_gathers_0_data_valid(accel_io_memStreams_gathers_0_data_valid),
    .io_memStreams_gathers_0_data_bits_0(accel_io_memStreams_gathers_0_data_bits_0),
    .io_memStreams_gathers_0_data_bits_1(accel_io_memStreams_gathers_0_data_bits_1),
    .io_memStreams_gathers_0_data_bits_2(accel_io_memStreams_gathers_0_data_bits_2),
    .io_memStreams_gathers_0_data_bits_3(accel_io_memStreams_gathers_0_data_bits_3),
    .io_memStreams_gathers_0_data_bits_4(accel_io_memStreams_gathers_0_data_bits_4),
    .io_memStreams_gathers_0_data_bits_5(accel_io_memStreams_gathers_0_data_bits_5),
    .io_memStreams_gathers_0_data_bits_6(accel_io_memStreams_gathers_0_data_bits_6),
    .io_memStreams_gathers_0_data_bits_7(accel_io_memStreams_gathers_0_data_bits_7),
    .io_memStreams_gathers_0_data_bits_8(accel_io_memStreams_gathers_0_data_bits_8),
    .io_memStreams_gathers_0_data_bits_9(accel_io_memStreams_gathers_0_data_bits_9),
    .io_memStreams_gathers_0_data_bits_10(accel_io_memStreams_gathers_0_data_bits_10),
    .io_memStreams_gathers_0_data_bits_11(accel_io_memStreams_gathers_0_data_bits_11),
    .io_memStreams_gathers_0_data_bits_12(accel_io_memStreams_gathers_0_data_bits_12),
    .io_memStreams_gathers_0_data_bits_13(accel_io_memStreams_gathers_0_data_bits_13),
    .io_memStreams_gathers_0_data_bits_14(accel_io_memStreams_gathers_0_data_bits_14),
    .io_memStreams_gathers_0_data_bits_15(accel_io_memStreams_gathers_0_data_bits_15),
    .io_memStreams_scatters_0_cmd_ready(accel_io_memStreams_scatters_0_cmd_ready),
    .io_memStreams_scatters_0_cmd_valid(accel_io_memStreams_scatters_0_cmd_valid),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_0(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_1(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_2(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_3(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_4(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_5(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_6(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_7(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_8(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_9(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_10(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_11(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_12(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_13(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_14(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_15(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15),
    .io_memStreams_scatters_0_cmd_bits_wdata_0(accel_io_memStreams_scatters_0_cmd_bits_wdata_0),
    .io_memStreams_scatters_0_cmd_bits_wdata_1(accel_io_memStreams_scatters_0_cmd_bits_wdata_1),
    .io_memStreams_scatters_0_cmd_bits_wdata_2(accel_io_memStreams_scatters_0_cmd_bits_wdata_2),
    .io_memStreams_scatters_0_cmd_bits_wdata_3(accel_io_memStreams_scatters_0_cmd_bits_wdata_3),
    .io_memStreams_scatters_0_cmd_bits_wdata_4(accel_io_memStreams_scatters_0_cmd_bits_wdata_4),
    .io_memStreams_scatters_0_cmd_bits_wdata_5(accel_io_memStreams_scatters_0_cmd_bits_wdata_5),
    .io_memStreams_scatters_0_cmd_bits_wdata_6(accel_io_memStreams_scatters_0_cmd_bits_wdata_6),
    .io_memStreams_scatters_0_cmd_bits_wdata_7(accel_io_memStreams_scatters_0_cmd_bits_wdata_7),
    .io_memStreams_scatters_0_cmd_bits_wdata_8(accel_io_memStreams_scatters_0_cmd_bits_wdata_8),
    .io_memStreams_scatters_0_cmd_bits_wdata_9(accel_io_memStreams_scatters_0_cmd_bits_wdata_9),
    .io_memStreams_scatters_0_cmd_bits_wdata_10(accel_io_memStreams_scatters_0_cmd_bits_wdata_10),
    .io_memStreams_scatters_0_cmd_bits_wdata_11(accel_io_memStreams_scatters_0_cmd_bits_wdata_11),
    .io_memStreams_scatters_0_cmd_bits_wdata_12(accel_io_memStreams_scatters_0_cmd_bits_wdata_12),
    .io_memStreams_scatters_0_cmd_bits_wdata_13(accel_io_memStreams_scatters_0_cmd_bits_wdata_13),
    .io_memStreams_scatters_0_cmd_bits_wdata_14(accel_io_memStreams_scatters_0_cmd_bits_wdata_14),
    .io_memStreams_scatters_0_cmd_bits_wdata_15(accel_io_memStreams_scatters_0_cmd_bits_wdata_15),
    .io_memStreams_scatters_0_wresp_ready(accel_io_memStreams_scatters_0_wresp_ready),
    .io_memStreams_scatters_0_wresp_valid(accel_io_memStreams_scatters_0_wresp_valid),
    .io_memStreams_scatters_0_wresp_bits(accel_io_memStreams_scatters_0_wresp_bits),
    .io_heap_0_req_valid(accel_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(accel_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(accel_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(accel_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(accel_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(accel_io_heap_0_resp_bits_sizeAddr),
    .io_argIns_0(accel_io_argIns_0),
    .io_argOuts_0_port_ready(accel_io_argOuts_0_port_ready),
    .io_argOuts_0_port_valid(accel_io_argOuts_0_port_valid),
    .io_argOuts_0_port_bits(accel_io_argOuts_0_port_bits),
    .io_argOuts_0_echo(accel_io_argOuts_0_echo),
    .io_argOuts_1_port_ready(accel_io_argOuts_1_port_ready),
    .io_argOuts_1_port_valid(accel_io_argOuts_1_port_valid),
    .io_argOuts_1_port_bits(accel_io_argOuts_1_port_bits),
    .io_argOuts_1_echo(accel_io_argOuts_1_echo),
    .io_argOuts_2_port_ready(accel_io_argOuts_2_port_ready),
    .io_argOuts_2_port_valid(accel_io_argOuts_2_port_valid),
    .io_argOuts_2_port_bits(accel_io_argOuts_2_port_bits),
    .io_argOuts_2_echo(accel_io_argOuts_2_echo),
    .io_argOuts_3_port_ready(accel_io_argOuts_3_port_ready),
    .io_argOuts_3_port_valid(accel_io_argOuts_3_port_valid),
    .io_argOuts_3_port_bits(accel_io_argOuts_3_port_bits),
    .io_argOuts_3_echo(accel_io_argOuts_3_echo),
    .io_argOuts_4_port_ready(accel_io_argOuts_4_port_ready),
    .io_argOuts_4_port_valid(accel_io_argOuts_4_port_valid),
    .io_argOuts_4_port_bits(accel_io_argOuts_4_port_bits),
    .io_argOuts_4_echo(accel_io_argOuts_4_echo),
    .io_argOuts_5_port_ready(accel_io_argOuts_5_port_ready),
    .io_argOuts_5_port_valid(accel_io_argOuts_5_port_valid),
    .io_argOuts_5_port_bits(accel_io_argOuts_5_port_bits),
    .io_argOuts_5_echo(accel_io_argOuts_5_echo),
    .io_argOuts_6_port_ready(accel_io_argOuts_6_port_ready),
    .io_argOuts_6_port_valid(accel_io_argOuts_6_port_valid),
    .io_argOuts_6_port_bits(accel_io_argOuts_6_port_bits),
    .io_argOuts_6_echo(accel_io_argOuts_6_echo),
    .io_argOuts_7_port_ready(accel_io_argOuts_7_port_ready),
    .io_argOuts_7_port_valid(accel_io_argOuts_7_port_valid),
    .io_argOuts_7_port_bits(accel_io_argOuts_7_port_bits),
    .io_argOuts_7_echo(accel_io_argOuts_7_echo),
    .io_argOuts_8_port_ready(accel_io_argOuts_8_port_ready),
    .io_argOuts_8_port_valid(accel_io_argOuts_8_port_valid),
    .io_argOuts_8_port_bits(accel_io_argOuts_8_port_bits),
    .io_argOuts_8_echo(accel_io_argOuts_8_echo),
    .io_argOuts_9_port_ready(accel_io_argOuts_9_port_ready),
    .io_argOuts_9_port_valid(accel_io_argOuts_9_port_valid),
    .io_argOuts_9_port_bits(accel_io_argOuts_9_port_bits),
    .io_argOuts_9_echo(accel_io_argOuts_9_echo),
    .io_argOuts_10_port_ready(accel_io_argOuts_10_port_ready),
    .io_argOuts_10_port_valid(accel_io_argOuts_10_port_valid),
    .io_argOuts_10_port_bits(accel_io_argOuts_10_port_bits),
    .io_argOuts_10_echo(accel_io_argOuts_10_echo),
    .io_argOuts_11_port_ready(accel_io_argOuts_11_port_ready),
    .io_argOuts_11_port_valid(accel_io_argOuts_11_port_valid),
    .io_argOuts_11_port_bits(accel_io_argOuts_11_port_bits),
    .io_argOuts_11_echo(accel_io_argOuts_11_echo),
    .io_argOuts_12_port_ready(accel_io_argOuts_12_port_ready),
    .io_argOuts_12_port_valid(accel_io_argOuts_12_port_valid),
    .io_argOuts_12_port_bits(accel_io_argOuts_12_port_bits),
    .io_argOuts_12_echo(accel_io_argOuts_12_echo),
    .io_argOuts_13_port_ready(accel_io_argOuts_13_port_ready),
    .io_argOuts_13_port_valid(accel_io_argOuts_13_port_valid),
    .io_argOuts_13_port_bits(accel_io_argOuts_13_port_bits),
    .io_argOuts_13_echo(accel_io_argOuts_13_echo),
    .io_argOuts_14_port_ready(accel_io_argOuts_14_port_ready),
    .io_argOuts_14_port_valid(accel_io_argOuts_14_port_valid),
    .io_argOuts_14_port_bits(accel_io_argOuts_14_port_bits),
    .io_argOuts_14_echo(accel_io_argOuts_14_echo),
    .io_argOuts_15_port_ready(accel_io_argOuts_15_port_ready),
    .io_argOuts_15_port_valid(accel_io_argOuts_15_port_valid),
    .io_argOuts_15_port_bits(accel_io_argOuts_15_port_bits),
    .io_argOuts_15_echo(accel_io_argOuts_15_echo)
  );
  FringeZynq FringeZynq ( // @[KCU1500.scala 21:24:@64727.4]
    .clock(FringeZynq_clock),
    .reset(FringeZynq_reset),
    .io_S_AXI_AWADDR(FringeZynq_io_S_AXI_AWADDR),
    .io_S_AXI_AWPROT(FringeZynq_io_S_AXI_AWPROT),
    .io_S_AXI_AWVALID(FringeZynq_io_S_AXI_AWVALID),
    .io_S_AXI_AWREADY(FringeZynq_io_S_AXI_AWREADY),
    .io_S_AXI_ARADDR(FringeZynq_io_S_AXI_ARADDR),
    .io_S_AXI_ARPROT(FringeZynq_io_S_AXI_ARPROT),
    .io_S_AXI_ARVALID(FringeZynq_io_S_AXI_ARVALID),
    .io_S_AXI_ARREADY(FringeZynq_io_S_AXI_ARREADY),
    .io_S_AXI_WDATA(FringeZynq_io_S_AXI_WDATA),
    .io_S_AXI_WSTRB(FringeZynq_io_S_AXI_WSTRB),
    .io_S_AXI_WVALID(FringeZynq_io_S_AXI_WVALID),
    .io_S_AXI_WREADY(FringeZynq_io_S_AXI_WREADY),
    .io_S_AXI_RDATA(FringeZynq_io_S_AXI_RDATA),
    .io_S_AXI_RRESP(FringeZynq_io_S_AXI_RRESP),
    .io_S_AXI_RVALID(FringeZynq_io_S_AXI_RVALID),
    .io_S_AXI_RREADY(FringeZynq_io_S_AXI_RREADY),
    .io_S_AXI_BRESP(FringeZynq_io_S_AXI_BRESP),
    .io_S_AXI_BVALID(FringeZynq_io_S_AXI_BVALID),
    .io_S_AXI_BREADY(FringeZynq_io_S_AXI_BREADY),
    .io_M_AXI_0_AWID(FringeZynq_io_M_AXI_0_AWID),
    .io_M_AXI_0_AWADDR(FringeZynq_io_M_AXI_0_AWADDR),
    .io_M_AXI_0_AWLEN(FringeZynq_io_M_AXI_0_AWLEN),
    .io_M_AXI_0_ARID(FringeZynq_io_M_AXI_0_ARID),
    .io_M_AXI_0_ARADDR(FringeZynq_io_M_AXI_0_ARADDR),
    .io_M_AXI_0_ARLEN(FringeZynq_io_M_AXI_0_ARLEN),
    .io_M_AXI_0_ARVALID(FringeZynq_io_M_AXI_0_ARVALID),
    .io_M_AXI_0_ARREADY(FringeZynq_io_M_AXI_0_ARREADY),
    .io_M_AXI_0_WLAST(FringeZynq_io_M_AXI_0_WLAST),
    .io_M_AXI_0_WREADY(FringeZynq_io_M_AXI_0_WREADY),
    .io_M_AXI_0_RID(FringeZynq_io_M_AXI_0_RID),
    .io_M_AXI_0_RDATA(FringeZynq_io_M_AXI_0_RDATA),
    .io_M_AXI_0_RVALID(FringeZynq_io_M_AXI_0_RVALID),
    .io_M_AXI_0_RREADY(FringeZynq_io_M_AXI_0_RREADY),
    .io_M_AXI_0_BID(FringeZynq_io_M_AXI_0_BID),
    .io_M_AXI_0_BVALID(FringeZynq_io_M_AXI_0_BVALID),
    .io_M_AXI_0_BREADY(FringeZynq_io_M_AXI_0_BREADY),
    .io_enable(FringeZynq_io_enable),
    .io_done(FringeZynq_io_done),
    .io_reset(FringeZynq_io_reset),
    .io_argIns_0(FringeZynq_io_argIns_0),
    .io_argOuts_0_valid(FringeZynq_io_argOuts_0_valid),
    .io_argOuts_0_bits(FringeZynq_io_argOuts_0_bits),
    .io_argOuts_1_valid(FringeZynq_io_argOuts_1_valid),
    .io_argOuts_1_bits(FringeZynq_io_argOuts_1_bits),
    .io_argOuts_2_valid(FringeZynq_io_argOuts_2_valid),
    .io_argOuts_2_bits(FringeZynq_io_argOuts_2_bits),
    .io_argOuts_3_valid(FringeZynq_io_argOuts_3_valid),
    .io_argOuts_3_bits(FringeZynq_io_argOuts_3_bits),
    .io_argOuts_4_valid(FringeZynq_io_argOuts_4_valid),
    .io_argOuts_4_bits(FringeZynq_io_argOuts_4_bits),
    .io_argOuts_5_valid(FringeZynq_io_argOuts_5_valid),
    .io_argOuts_5_bits(FringeZynq_io_argOuts_5_bits),
    .io_argOuts_6_valid(FringeZynq_io_argOuts_6_valid),
    .io_argOuts_6_bits(FringeZynq_io_argOuts_6_bits),
    .io_argOuts_7_valid(FringeZynq_io_argOuts_7_valid),
    .io_argOuts_7_bits(FringeZynq_io_argOuts_7_bits),
    .io_argOuts_8_valid(FringeZynq_io_argOuts_8_valid),
    .io_argOuts_8_bits(FringeZynq_io_argOuts_8_bits),
    .io_argOuts_9_valid(FringeZynq_io_argOuts_9_valid),
    .io_argOuts_9_bits(FringeZynq_io_argOuts_9_bits),
    .io_argOuts_10_valid(FringeZynq_io_argOuts_10_valid),
    .io_argOuts_10_bits(FringeZynq_io_argOuts_10_bits),
    .io_argOuts_11_valid(FringeZynq_io_argOuts_11_valid),
    .io_argOuts_11_bits(FringeZynq_io_argOuts_11_bits),
    .io_argOuts_12_valid(FringeZynq_io_argOuts_12_valid),
    .io_argOuts_12_bits(FringeZynq_io_argOuts_12_bits),
    .io_argOuts_13_valid(FringeZynq_io_argOuts_13_valid),
    .io_argOuts_13_bits(FringeZynq_io_argOuts_13_bits),
    .io_argOuts_14_valid(FringeZynq_io_argOuts_14_valid),
    .io_argOuts_14_bits(FringeZynq_io_argOuts_14_bits),
    .io_argOuts_15_valid(FringeZynq_io_argOuts_15_valid),
    .io_argOuts_15_bits(FringeZynq_io_argOuts_15_bits),
    .io_memStreams_loads_0_cmd_ready(FringeZynq_io_memStreams_loads_0_cmd_ready),
    .io_memStreams_loads_0_cmd_valid(FringeZynq_io_memStreams_loads_0_cmd_valid),
    .io_memStreams_loads_0_cmd_bits_addr(FringeZynq_io_memStreams_loads_0_cmd_bits_addr),
    .io_memStreams_loads_0_cmd_bits_size(FringeZynq_io_memStreams_loads_0_cmd_bits_size),
    .io_memStreams_loads_0_data_ready(FringeZynq_io_memStreams_loads_0_data_ready),
    .io_memStreams_loads_0_data_valid(FringeZynq_io_memStreams_loads_0_data_valid),
    .io_memStreams_loads_0_data_bits_rdata_0(FringeZynq_io_memStreams_loads_0_data_bits_rdata_0),
    .io_memStreams_stores_0_cmd_valid(FringeZynq_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(FringeZynq_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(FringeZynq_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_valid(FringeZynq_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(FringeZynq_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wstrb(FringeZynq_io_memStreams_stores_0_data_bits_wstrb),
    .io_heap_0_req_valid(FringeZynq_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(FringeZynq_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(FringeZynq_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(FringeZynq_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(FringeZynq_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(FringeZynq_io_heap_0_resp_bits_sizeAddr)
  );
  assign io_rdata = 1'h0;
  assign io_S_AXI_AWREADY = FringeZynq_io_S_AXI_AWREADY; // @[KCU1500.scala 24:21:@64745.4]
  assign io_S_AXI_ARREADY = FringeZynq_io_S_AXI_ARREADY; // @[KCU1500.scala 24:21:@64741.4]
  assign io_S_AXI_WREADY = FringeZynq_io_S_AXI_WREADY; // @[KCU1500.scala 24:21:@64737.4]
  assign io_S_AXI_RDATA = FringeZynq_io_S_AXI_RDATA; // @[KCU1500.scala 24:21:@64736.4]
  assign io_S_AXI_RRESP = FringeZynq_io_S_AXI_RRESP; // @[KCU1500.scala 24:21:@64735.4]
  assign io_S_AXI_RVALID = FringeZynq_io_S_AXI_RVALID; // @[KCU1500.scala 24:21:@64734.4]
  assign io_S_AXI_BRESP = FringeZynq_io_S_AXI_BRESP; // @[KCU1500.scala 24:21:@64732.4]
  assign io_S_AXI_BVALID = FringeZynq_io_S_AXI_BVALID; // @[KCU1500.scala 24:21:@64731.4]
  assign io_M_AXI_0_AWID = FringeZynq_io_M_AXI_0_AWID; // @[KCU1500.scala 27:14:@64789.4]
  assign io_M_AXI_0_AWUSER = 4'h0; // @[KCU1500.scala 27:14:@64788.4]
  assign io_M_AXI_0_AWADDR = FringeZynq_io_M_AXI_0_AWADDR; // @[KCU1500.scala 27:14:@64787.4]
  assign io_M_AXI_0_AWLEN = FringeZynq_io_M_AXI_0_AWLEN; // @[KCU1500.scala 27:14:@64786.4]
  assign io_M_AXI_0_AWSIZE = 3'h6; // @[KCU1500.scala 27:14:@64785.4]
  assign io_M_AXI_0_AWBURST = 2'h1; // @[KCU1500.scala 27:14:@64784.4]
  assign io_M_AXI_0_AWLOCK = 1'h0; // @[KCU1500.scala 27:14:@64783.4]
  assign io_M_AXI_0_AWCACHE = 4'h3; // @[KCU1500.scala 27:14:@64782.4]
  assign io_M_AXI_0_AWPROT = 3'h0; // @[KCU1500.scala 27:14:@64781.4]
  assign io_M_AXI_0_AWQOS = 4'h0; // @[KCU1500.scala 27:14:@64780.4]
  assign io_M_AXI_0_AWVALID = 1'h0; // @[KCU1500.scala 27:14:@64779.4]
  assign io_M_AXI_0_ARID = FringeZynq_io_M_AXI_0_ARID; // @[KCU1500.scala 27:14:@64777.4]
  assign io_M_AXI_0_ARUSER = 4'h0; // @[KCU1500.scala 27:14:@64776.4]
  assign io_M_AXI_0_ARADDR = FringeZynq_io_M_AXI_0_ARADDR; // @[KCU1500.scala 27:14:@64775.4]
  assign io_M_AXI_0_ARLEN = FringeZynq_io_M_AXI_0_ARLEN; // @[KCU1500.scala 27:14:@64774.4]
  assign io_M_AXI_0_ARSIZE = 3'h6; // @[KCU1500.scala 27:14:@64773.4]
  assign io_M_AXI_0_ARBURST = 2'h1; // @[KCU1500.scala 27:14:@64772.4]
  assign io_M_AXI_0_ARLOCK = 1'h0; // @[KCU1500.scala 27:14:@64771.4]
  assign io_M_AXI_0_ARCACHE = 4'h3; // @[KCU1500.scala 27:14:@64770.4]
  assign io_M_AXI_0_ARPROT = 3'h0; // @[KCU1500.scala 27:14:@64769.4]
  assign io_M_AXI_0_ARQOS = 4'h0; // @[KCU1500.scala 27:14:@64768.4]
  assign io_M_AXI_0_ARVALID = FringeZynq_io_M_AXI_0_ARVALID; // @[KCU1500.scala 27:14:@64767.4]
  assign io_M_AXI_0_WDATA = 512'h0; // @[KCU1500.scala 27:14:@64765.4]
  assign io_M_AXI_0_WSTRB = 64'h0; // @[KCU1500.scala 27:14:@64764.4]
  assign io_M_AXI_0_WLAST = FringeZynq_io_M_AXI_0_WLAST; // @[KCU1500.scala 27:14:@64763.4]
  assign io_M_AXI_0_WVALID = 1'h0; // @[KCU1500.scala 27:14:@64762.4]
  assign io_M_AXI_0_RREADY = FringeZynq_io_M_AXI_0_RREADY; // @[KCU1500.scala 27:14:@64754.4]
  assign io_M_AXI_0_BREADY = FringeZynq_io_M_AXI_0_BREADY; // @[KCU1500.scala 27:14:@64749.4]
  assign accel_clock = clock; // @[:@64545.4]
  assign accel_reset = FringeZynq_io_reset; // @[:@64546.4 KCU1500.scala 57:17:@65121.4]
  assign accel_io_enable = FringeZynq_io_enable; // @[KCU1500.scala 54:21:@65117.4]
  assign accel_io_reset = 1'h0;
  assign accel_io_memStreams_loads_0_cmd_ready = FringeZynq_io_memStreams_loads_0_cmd_ready; // @[KCU1500.scala 52:26:@65110.4]
  assign accel_io_memStreams_loads_0_data_valid = FringeZynq_io_memStreams_loads_0_data_valid; // @[KCU1500.scala 52:26:@65105.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_0 = FringeZynq_io_memStreams_loads_0_data_bits_rdata_0; // @[KCU1500.scala 52:26:@65104.4]
  assign accel_io_memStreams_stores_0_cmd_ready = 1'h0; // @[KCU1500.scala 52:26:@65103.4]
  assign accel_io_memStreams_stores_0_data_ready = 1'h0; // @[KCU1500.scala 52:26:@65099.4]
  assign accel_io_memStreams_stores_0_wresp_valid = 1'h0; // @[KCU1500.scala 52:26:@65079.4]
  assign accel_io_memStreams_stores_0_wresp_bits = 1'h0; // @[KCU1500.scala 52:26:@65078.4]
  assign accel_io_memStreams_gathers_0_cmd_ready = 1'h0; // @[KCU1500.scala 52:26:@65077.4]
  assign accel_io_memStreams_gathers_0_data_valid = 1'h0; // @[KCU1500.scala 52:26:@65058.4]
  assign accel_io_memStreams_gathers_0_data_bits_0 = 32'h0; // @[KCU1500.scala 52:26:@65042.4]
  assign accel_io_memStreams_gathers_0_data_bits_1 = 32'h0; // @[KCU1500.scala 52:26:@65043.4]
  assign accel_io_memStreams_gathers_0_data_bits_2 = 32'h0; // @[KCU1500.scala 52:26:@65044.4]
  assign accel_io_memStreams_gathers_0_data_bits_3 = 32'h0; // @[KCU1500.scala 52:26:@65045.4]
  assign accel_io_memStreams_gathers_0_data_bits_4 = 32'h0; // @[KCU1500.scala 52:26:@65046.4]
  assign accel_io_memStreams_gathers_0_data_bits_5 = 32'h0; // @[KCU1500.scala 52:26:@65047.4]
  assign accel_io_memStreams_gathers_0_data_bits_6 = 32'h0; // @[KCU1500.scala 52:26:@65048.4]
  assign accel_io_memStreams_gathers_0_data_bits_7 = 32'h0; // @[KCU1500.scala 52:26:@65049.4]
  assign accel_io_memStreams_gathers_0_data_bits_8 = 32'h0; // @[KCU1500.scala 52:26:@65050.4]
  assign accel_io_memStreams_gathers_0_data_bits_9 = 32'h0; // @[KCU1500.scala 52:26:@65051.4]
  assign accel_io_memStreams_gathers_0_data_bits_10 = 32'h0; // @[KCU1500.scala 52:26:@65052.4]
  assign accel_io_memStreams_gathers_0_data_bits_11 = 32'h0; // @[KCU1500.scala 52:26:@65053.4]
  assign accel_io_memStreams_gathers_0_data_bits_12 = 32'h0; // @[KCU1500.scala 52:26:@65054.4]
  assign accel_io_memStreams_gathers_0_data_bits_13 = 32'h0; // @[KCU1500.scala 52:26:@65055.4]
  assign accel_io_memStreams_gathers_0_data_bits_14 = 32'h0; // @[KCU1500.scala 52:26:@65056.4]
  assign accel_io_memStreams_gathers_0_data_bits_15 = 32'h0; // @[KCU1500.scala 52:26:@65057.4]
  assign accel_io_memStreams_scatters_0_cmd_ready = 1'h0; // @[KCU1500.scala 52:26:@65041.4]
  assign accel_io_memStreams_scatters_0_wresp_valid = 1'h0; // @[KCU1500.scala 52:26:@65006.4]
  assign accel_io_memStreams_scatters_0_wresp_bits = 1'h0; // @[KCU1500.scala 52:26:@65005.4]
  assign accel_io_heap_0_resp_valid = FringeZynq_io_heap_0_resp_valid; // @[KCU1500.scala 53:20:@65113.4]
  assign accel_io_heap_0_resp_bits_allocDealloc = FringeZynq_io_heap_0_resp_bits_allocDealloc; // @[KCU1500.scala 53:20:@65112.4]
  assign accel_io_heap_0_resp_bits_sizeAddr = FringeZynq_io_heap_0_resp_bits_sizeAddr; // @[KCU1500.scala 53:20:@65111.4]
  assign accel_io_argIns_0 = FringeZynq_io_argIns_0; // @[KCU1500.scala 37:21:@64955.4]
  assign accel_io_argOuts_0_port_ready = 1'h0;
  assign accel_io_argOuts_0_echo = 64'h0; // @[KCU1500.scala 43:24:@64988.4]
  assign accel_io_argOuts_1_port_ready = 1'h0;
  assign accel_io_argOuts_1_echo = 64'h0; // @[KCU1500.scala 43:24:@64989.4]
  assign accel_io_argOuts_2_port_ready = 1'h0;
  assign accel_io_argOuts_2_echo = 64'h0; // @[KCU1500.scala 43:24:@64990.4]
  assign accel_io_argOuts_3_port_ready = 1'h0;
  assign accel_io_argOuts_3_echo = 64'h0; // @[KCU1500.scala 43:24:@64991.4]
  assign accel_io_argOuts_4_port_ready = 1'h0;
  assign accel_io_argOuts_4_echo = 64'h0; // @[KCU1500.scala 43:24:@64992.4]
  assign accel_io_argOuts_5_port_ready = 1'h0;
  assign accel_io_argOuts_5_echo = 64'h0; // @[KCU1500.scala 43:24:@64993.4]
  assign accel_io_argOuts_6_port_ready = 1'h0;
  assign accel_io_argOuts_6_echo = 64'h0; // @[KCU1500.scala 43:24:@64994.4]
  assign accel_io_argOuts_7_port_ready = 1'h0;
  assign accel_io_argOuts_7_echo = 64'h0; // @[KCU1500.scala 43:24:@64995.4]
  assign accel_io_argOuts_8_port_ready = 1'h0;
  assign accel_io_argOuts_8_echo = 64'h0; // @[KCU1500.scala 43:24:@64996.4]
  assign accel_io_argOuts_9_port_ready = 1'h0;
  assign accel_io_argOuts_9_echo = 64'h0; // @[KCU1500.scala 43:24:@64997.4]
  assign accel_io_argOuts_10_port_ready = 1'h0;
  assign accel_io_argOuts_10_echo = 64'h0; // @[KCU1500.scala 43:24:@64998.4]
  assign accel_io_argOuts_11_port_ready = 1'h0;
  assign accel_io_argOuts_11_echo = 64'h0; // @[KCU1500.scala 43:24:@64999.4]
  assign accel_io_argOuts_12_port_ready = 1'h0;
  assign accel_io_argOuts_12_echo = 64'h0; // @[KCU1500.scala 43:24:@65000.4]
  assign accel_io_argOuts_13_port_ready = 1'h0;
  assign accel_io_argOuts_13_echo = 64'h0; // @[KCU1500.scala 43:24:@65001.4]
  assign accel_io_argOuts_14_port_ready = 1'h0;
  assign accel_io_argOuts_14_echo = 64'h0; // @[KCU1500.scala 43:24:@65002.4]
  assign accel_io_argOuts_15_port_ready = 1'h0;
  assign accel_io_argOuts_15_echo = 64'h0; // @[KCU1500.scala 43:24:@65003.4]
  assign FringeZynq_clock = clock; // @[:@64728.4]
  assign FringeZynq_reset = reset; // @[:@64729.4 KCU1500.scala 56:18:@65120.4]
  assign FringeZynq_io_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[KCU1500.scala 24:21:@64748.4]
  assign FringeZynq_io_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[KCU1500.scala 24:21:@64747.4]
  assign FringeZynq_io_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[KCU1500.scala 24:21:@64746.4]
  assign FringeZynq_io_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[KCU1500.scala 24:21:@64744.4]
  assign FringeZynq_io_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[KCU1500.scala 24:21:@64743.4]
  assign FringeZynq_io_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[KCU1500.scala 24:21:@64742.4]
  assign FringeZynq_io_S_AXI_WDATA = io_S_AXI_WDATA; // @[KCU1500.scala 24:21:@64740.4]
  assign FringeZynq_io_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[KCU1500.scala 24:21:@64739.4]
  assign FringeZynq_io_S_AXI_WVALID = io_S_AXI_WVALID; // @[KCU1500.scala 24:21:@64738.4]
  assign FringeZynq_io_S_AXI_RREADY = io_S_AXI_RREADY; // @[KCU1500.scala 24:21:@64733.4]
  assign FringeZynq_io_S_AXI_BREADY = io_S_AXI_BREADY; // @[KCU1500.scala 24:21:@64730.4]
  assign FringeZynq_io_M_AXI_0_ARREADY = io_M_AXI_0_ARREADY; // @[KCU1500.scala 27:14:@64766.4]
  assign FringeZynq_io_M_AXI_0_WREADY = io_M_AXI_0_WREADY; // @[KCU1500.scala 27:14:@64761.4]
  assign FringeZynq_io_M_AXI_0_RID = io_M_AXI_0_RID; // @[KCU1500.scala 27:14:@64760.4]
  assign FringeZynq_io_M_AXI_0_RDATA = io_M_AXI_0_RDATA; // @[KCU1500.scala 27:14:@64758.4]
  assign FringeZynq_io_M_AXI_0_RVALID = io_M_AXI_0_RVALID; // @[KCU1500.scala 27:14:@64755.4]
  assign FringeZynq_io_M_AXI_0_BID = io_M_AXI_0_BID; // @[KCU1500.scala 27:14:@64753.4]
  assign FringeZynq_io_M_AXI_0_BVALID = io_M_AXI_0_BVALID; // @[KCU1500.scala 27:14:@64750.4]
  assign FringeZynq_io_done = accel_io_done; // @[KCU1500.scala 55:20:@65118.4]
  assign FringeZynq_io_argOuts_0_valid = accel_io_argOuts_0_port_valid; // @[KCU1500.scala 40:26:@64957.4]
  assign FringeZynq_io_argOuts_0_bits = accel_io_argOuts_0_port_bits; // @[KCU1500.scala 39:25:@64956.4]
  assign FringeZynq_io_argOuts_1_valid = accel_io_argOuts_1_port_valid; // @[KCU1500.scala 40:26:@64959.4]
  assign FringeZynq_io_argOuts_1_bits = accel_io_argOuts_1_port_bits; // @[KCU1500.scala 39:25:@64958.4]
  assign FringeZynq_io_argOuts_2_valid = accel_io_argOuts_2_port_valid; // @[KCU1500.scala 40:26:@64961.4]
  assign FringeZynq_io_argOuts_2_bits = accel_io_argOuts_2_port_bits; // @[KCU1500.scala 39:25:@64960.4]
  assign FringeZynq_io_argOuts_3_valid = accel_io_argOuts_3_port_valid; // @[KCU1500.scala 40:26:@64963.4]
  assign FringeZynq_io_argOuts_3_bits = accel_io_argOuts_3_port_bits; // @[KCU1500.scala 39:25:@64962.4]
  assign FringeZynq_io_argOuts_4_valid = accel_io_argOuts_4_port_valid; // @[KCU1500.scala 40:26:@64965.4]
  assign FringeZynq_io_argOuts_4_bits = accel_io_argOuts_4_port_bits; // @[KCU1500.scala 39:25:@64964.4]
  assign FringeZynq_io_argOuts_5_valid = accel_io_argOuts_5_port_valid; // @[KCU1500.scala 40:26:@64967.4]
  assign FringeZynq_io_argOuts_5_bits = accel_io_argOuts_5_port_bits; // @[KCU1500.scala 39:25:@64966.4]
  assign FringeZynq_io_argOuts_6_valid = accel_io_argOuts_6_port_valid; // @[KCU1500.scala 40:26:@64969.4]
  assign FringeZynq_io_argOuts_6_bits = accel_io_argOuts_6_port_bits; // @[KCU1500.scala 39:25:@64968.4]
  assign FringeZynq_io_argOuts_7_valid = accel_io_argOuts_7_port_valid; // @[KCU1500.scala 40:26:@64971.4]
  assign FringeZynq_io_argOuts_7_bits = accel_io_argOuts_7_port_bits; // @[KCU1500.scala 39:25:@64970.4]
  assign FringeZynq_io_argOuts_8_valid = accel_io_argOuts_8_port_valid; // @[KCU1500.scala 40:26:@64973.4]
  assign FringeZynq_io_argOuts_8_bits = accel_io_argOuts_8_port_bits; // @[KCU1500.scala 39:25:@64972.4]
  assign FringeZynq_io_argOuts_9_valid = accel_io_argOuts_9_port_valid; // @[KCU1500.scala 40:26:@64975.4]
  assign FringeZynq_io_argOuts_9_bits = accel_io_argOuts_9_port_bits; // @[KCU1500.scala 39:25:@64974.4]
  assign FringeZynq_io_argOuts_10_valid = accel_io_argOuts_10_port_valid; // @[KCU1500.scala 40:26:@64977.4]
  assign FringeZynq_io_argOuts_10_bits = accel_io_argOuts_10_port_bits; // @[KCU1500.scala 39:25:@64976.4]
  assign FringeZynq_io_argOuts_11_valid = accel_io_argOuts_11_port_valid; // @[KCU1500.scala 40:26:@64979.4]
  assign FringeZynq_io_argOuts_11_bits = accel_io_argOuts_11_port_bits; // @[KCU1500.scala 39:25:@64978.4]
  assign FringeZynq_io_argOuts_12_valid = accel_io_argOuts_12_port_valid; // @[KCU1500.scala 40:26:@64981.4]
  assign FringeZynq_io_argOuts_12_bits = accel_io_argOuts_12_port_bits; // @[KCU1500.scala 39:25:@64980.4]
  assign FringeZynq_io_argOuts_13_valid = accel_io_argOuts_13_port_valid; // @[KCU1500.scala 40:26:@64983.4]
  assign FringeZynq_io_argOuts_13_bits = accel_io_argOuts_13_port_bits; // @[KCU1500.scala 39:25:@64982.4]
  assign FringeZynq_io_argOuts_14_valid = accel_io_argOuts_14_port_valid; // @[KCU1500.scala 40:26:@64985.4]
  assign FringeZynq_io_argOuts_14_bits = accel_io_argOuts_14_port_bits; // @[KCU1500.scala 39:25:@64984.4]
  assign FringeZynq_io_argOuts_15_valid = accel_io_argOuts_15_port_valid; // @[KCU1500.scala 40:26:@64987.4]
  assign FringeZynq_io_argOuts_15_bits = accel_io_argOuts_15_port_bits; // @[KCU1500.scala 39:25:@64986.4]
  assign FringeZynq_io_memStreams_loads_0_cmd_valid = accel_io_memStreams_loads_0_cmd_valid; // @[KCU1500.scala 52:26:@65109.4]
  assign FringeZynq_io_memStreams_loads_0_cmd_bits_addr = accel_io_memStreams_loads_0_cmd_bits_addr; // @[KCU1500.scala 52:26:@65108.4]
  assign FringeZynq_io_memStreams_loads_0_cmd_bits_size = accel_io_memStreams_loads_0_cmd_bits_size; // @[KCU1500.scala 52:26:@65107.4]
  assign FringeZynq_io_memStreams_loads_0_data_ready = accel_io_memStreams_loads_0_data_ready; // @[KCU1500.scala 52:26:@65106.4]
  assign FringeZynq_io_memStreams_stores_0_cmd_valid = accel_io_memStreams_stores_0_cmd_valid; // @[KCU1500.scala 52:26:@65102.4]
  assign FringeZynq_io_memStreams_stores_0_cmd_bits_addr = accel_io_memStreams_stores_0_cmd_bits_addr; // @[KCU1500.scala 52:26:@65101.4]
  assign FringeZynq_io_memStreams_stores_0_cmd_bits_size = accel_io_memStreams_stores_0_cmd_bits_size; // @[KCU1500.scala 52:26:@65100.4]
  assign FringeZynq_io_memStreams_stores_0_data_valid = accel_io_memStreams_stores_0_data_valid; // @[KCU1500.scala 52:26:@65098.4]
  assign FringeZynq_io_memStreams_stores_0_data_bits_wdata_0 = accel_io_memStreams_stores_0_data_bits_wdata_0; // @[KCU1500.scala 52:26:@65082.4]
  assign FringeZynq_io_memStreams_stores_0_data_bits_wstrb = accel_io_memStreams_stores_0_data_bits_wstrb; // @[KCU1500.scala 52:26:@65081.4]
  assign FringeZynq_io_heap_0_req_valid = accel_io_heap_0_req_valid; // @[KCU1500.scala 53:20:@65116.4]
  assign FringeZynq_io_heap_0_req_bits_allocDealloc = accel_io_heap_0_req_bits_allocDealloc; // @[KCU1500.scala 53:20:@65115.4]
  assign FringeZynq_io_heap_0_req_bits_sizeAddr = accel_io_heap_0_req_bits_sizeAddr; // @[KCU1500.scala 53:20:@65114.4]
endmodule
module SRAMVerilogAWS
#(
    parameter WORDS = 1024,
    parameter AWIDTH = 10,
    parameter DWIDTH = 32)
(
    input clk,
    input [AWIDTH-1:0] raddr,
    input [AWIDTH-1:0] waddr,
    input raddrEn,
    input waddrEn,
    input wen,
    input [DWIDTH-1:0] wdata,
    input backpressure,
    output reg [DWIDTH-1:0] rdata
);

    reg [DWIDTH-1:0] mem [0:WORDS-1];

    always @(posedge clk) begin
      if (wen) mem[waddr] <= wdata;
      if (backpressure) rdata <= mem[raddr];
    end

endmodule
