module FF( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  output [31:0] io_rPort_0_output_0, // @[:@6.4]
  input  [31:0] io_wPort_0_data_0, // @[:@6.4]
  input         io_wPort_0_reset, // @[:@6.4]
  input         io_wPort_0_en_0 // @[:@6.4]
);
  reg [31:0] ff; // @[MemPrimitives.scala 173:19:@21.4]
  reg [31:0] _RAND_0;
  wire [31:0] _T_68; // @[MemPrimitives.scala 177:32:@23.4]
  wire [31:0] _T_69; // @[MemPrimitives.scala 177:12:@24.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 177:32:@23.4]
  assign _T_69 = io_wPort_0_reset ? 32'h0 : _T_68; // @[MemPrimitives.scala 177:12:@24.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 178:34:@26.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 32'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 32'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SRFF( // @[:@28.2]
  input   clock, // @[:@29.4]
  input   reset, // @[:@30.4]
  input   io_input_set, // @[:@31.4]
  input   io_input_reset, // @[:@31.4]
  input   io_input_asyn_reset, // @[:@31.4]
  output  io_output // @[:@31.4]
);
  reg  _T_15; // @[SRFF.scala 20:21:@33.4]
  reg [31:0] _RAND_0;
  wire  _T_19; // @[SRFF.scala 21:74:@34.4]
  wire  _T_20; // @[SRFF.scala 21:48:@35.4]
  wire  _T_21; // @[SRFF.scala 21:14:@36.4]
  assign _T_19 = io_input_reset ? 1'h0 : _T_15; // @[SRFF.scala 21:74:@34.4]
  assign _T_20 = io_input_set ? 1'h1 : _T_19; // @[SRFF.scala 21:48:@35.4]
  assign _T_21 = io_input_asyn_reset ? 1'h0 : _T_20; // @[SRFF.scala 21:14:@36.4]
  assign io_output = io_input_asyn_reset ? 1'h0 : _T_15; // @[SRFF.scala 22:15:@39.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_15 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_15 <= 1'h0;
    end else begin
      if (io_input_asyn_reset) begin
        _T_15 <= 1'h0;
      end else begin
        if (io_input_set) begin
          _T_15 <= 1'h1;
        end else begin
          if (io_input_reset) begin
            _T_15 <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module SingleCounter( // @[:@41.2]
  input   clock, // @[:@42.4]
  input   reset, // @[:@43.4]
  input   io_input_reset, // @[:@44.4]
  output  io_output_done // @[:@44.4]
);
  wire  bases_0_clock; // @[Counter.scala 253:53:@57.4]
  wire  bases_0_reset; // @[Counter.scala 253:53:@57.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 253:53:@57.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 253:53:@57.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 253:53:@57.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 253:53:@57.4]
  wire  SRFF_clock; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_reset; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_input_set; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_output; // @[Counter.scala 255:22:@73.4]
  wire [31:0] _T_48; // @[Counter.scala 279:52:@101.4]
  wire [32:0] _T_50; // @[Counter.scala 283:33:@102.4]
  wire [31:0] _T_51; // @[Counter.scala 283:33:@103.4]
  wire [31:0] _T_52; // @[Counter.scala 283:33:@104.4]
  wire  _T_57; // @[Counter.scala 285:18:@106.4]
  wire [31:0] _T_68; // @[Counter.scala 291:115:@114.4]
  wire [31:0] _T_71; // @[Counter.scala 291:152:@117.4]
  wire [31:0] _T_72; // @[Counter.scala 291:74:@118.4]
  FF bases_0 ( // @[Counter.scala 253:53:@57.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 255:22:@73.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 279:52:@101.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@102.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@103.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 283:33:@104.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh0); // @[Counter.scala 285:18:@106.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 291:115:@114.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 291:152:@117.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 291:74:@118.4]
  assign io_output_done = $signed(_T_52) >= $signed(32'sh0); // @[Counter.scala 325:20:@127.4]
  assign bases_0_clock = clock; // @[:@58.4]
  assign bases_0_reset = reset; // @[:@59.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 291:31:@120.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 273:27:@99.4]
  assign bases_0_io_wPort_0_en_0 = 1'h1; // @[Counter.scala 276:29:@100.4]
  assign SRFF_clock = clock; // @[:@74.4]
  assign SRFF_reset = reset; // @[:@75.4]
  assign SRFF_io_input_set = io_input_reset == 1'h0; // @[Counter.scala 256:23:@78.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 257:25:@80.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 258:30:@81.4]
endmodule
module RetimeWrapper( // @[:@144.2]
  input   clock, // @[:@145.4]
  input   reset, // @[:@146.4]
  input   io_flow, // @[:@147.4]
  input   io_in, // @[:@147.4]
  output  io_out // @[:@147.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@149.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@149.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@162.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@161.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@160.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@159.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@158.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@156.4]
endmodule
module RootController_sm( // @[:@351.2]
  input   clock, // @[:@352.4]
  input   reset, // @[:@353.4]
  input   io_enable, // @[:@354.4]
  output  io_done, // @[:@354.4]
  input   io_rst, // @[:@354.4]
  input   io_ctrDone, // @[:@354.4]
  output  io_ctrInc, // @[:@354.4]
  input   io_doneIn_0, // @[:@354.4]
  input   io_doneIn_1, // @[:@354.4]
  output  io_enableOut_0, // @[:@354.4]
  output  io_enableOut_1, // @[:@354.4]
  output  io_childAck_0, // @[:@354.4]
  output  io_childAck_1 // @[:@354.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@357.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@357.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@357.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@357.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@357.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@357.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@360.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@360.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@360.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@360.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@360.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@360.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@363.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@363.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@363.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@363.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@363.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@363.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@366.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@366.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@366.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@366.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@366.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@366.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@395.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@395.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@395.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@395.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@395.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@395.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@398.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@398.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@398.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@398.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@398.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@398.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@427.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@427.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@427.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@427.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@427.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@523.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@523.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@523.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@523.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@523.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@540.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@540.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@540.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@540.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@540.4]
  wire  allDone; // @[Controllers.scala 80:47:@369.4]
  wire  _T_77; // @[Controllers.scala 81:26:@370.4]
  wire  finished; // @[Controllers.scala 81:37:@371.4]
  wire  synchronize; // @[package.scala 96:25:@432.4 package.scala 96:25:@433.4]
  wire  _T_144; // @[Controllers.scala 128:33:@441.4]
  wire  _T_146; // @[Controllers.scala 128:54:@442.4]
  wire  _T_147; // @[Controllers.scala 128:52:@443.4]
  wire  _T_148; // @[Controllers.scala 128:66:@444.4]
  wire  _T_150; // @[Controllers.scala 128:98:@446.4]
  wire  _T_151; // @[Controllers.scala 128:96:@447.4]
  wire  _T_153; // @[Controllers.scala 128:123:@448.4]
  wire  _T_155; // @[Controllers.scala 129:48:@451.4]
  wire  _T_160; // @[Controllers.scala 130:52:@456.4]
  wire  _T_161; // @[Controllers.scala 130:50:@457.4]
  wire  _T_169; // @[Controllers.scala 130:129:@463.4]
  wire  _T_172; // @[Controllers.scala 131:45:@466.4]
  wire  _T_175; // @[Controllers.scala 135:80:@470.4]
  wire  _T_176; // @[Controllers.scala 135:78:@471.4]
  wire  _T_178; // @[Controllers.scala 135:105:@472.4]
  wire  _T_179; // @[Controllers.scala 135:103:@473.4]
  wire  _T_180; // @[Controllers.scala 135:119:@474.4]
  wire  _T_182; // @[Controllers.scala 135:51:@476.4]
  wire  _T_205; // @[Controllers.scala 213:68:@501.4]
  wire  _T_207; // @[Controllers.scala 213:90:@503.4]
  wire  _T_209; // @[Controllers.scala 213:132:@505.4]
  wire  _T_210; // @[Controllers.scala 213:130:@506.4]
  wire  _T_211; // @[Controllers.scala 213:156:@507.4]
  wire  _T_213; // @[Controllers.scala 213:68:@510.4]
  wire  _T_215; // @[Controllers.scala 213:90:@512.4]
  wire  _T_222; // @[package.scala 100:49:@518.4]
  reg  _T_225; // @[package.scala 48:56:@519.4]
  reg [31:0] _RAND_0;
  reg  _T_239; // @[package.scala 48:56:@537.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@357.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@360.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@363.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@366.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@395.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@398.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@427.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@523.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@540.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  assign allDone = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@369.4]
  assign _T_77 = allDone | io_done; // @[Controllers.scala 81:26:@370.4]
  assign finished = _T_77 | done_1_io_input_set; // @[Controllers.scala 81:37:@371.4]
  assign synchronize = RetimeWrapper_io_out; // @[package.scala 96:25:@432.4 package.scala 96:25:@433.4]
  assign _T_144 = done_0_io_output == 1'h0; // @[Controllers.scala 128:33:@441.4]
  assign _T_146 = io_ctrDone == 1'h0; // @[Controllers.scala 128:54:@442.4]
  assign _T_147 = _T_144 & _T_146; // @[Controllers.scala 128:52:@443.4]
  assign _T_148 = _T_147 & io_enable; // @[Controllers.scala 128:66:@444.4]
  assign _T_150 = ~ iterDone_0_io_output; // @[Controllers.scala 128:98:@446.4]
  assign _T_151 = _T_148 & _T_150; // @[Controllers.scala 128:96:@447.4]
  assign _T_153 = io_doneIn_0 == 1'h0; // @[Controllers.scala 128:123:@448.4]
  assign _T_155 = io_doneIn_0 | io_rst; // @[Controllers.scala 129:48:@451.4]
  assign _T_160 = synchronize == 1'h0; // @[Controllers.scala 130:52:@456.4]
  assign _T_161 = io_doneIn_0 & _T_160; // @[Controllers.scala 130:50:@457.4]
  assign _T_169 = finished == 1'h0; // @[Controllers.scala 130:129:@463.4]
  assign _T_172 = io_rst == 1'h0; // @[Controllers.scala 131:45:@466.4]
  assign _T_175 = ~ iterDone_1_io_output; // @[Controllers.scala 135:80:@470.4]
  assign _T_176 = iterDone_0_io_output & _T_175; // @[Controllers.scala 135:78:@471.4]
  assign _T_178 = io_doneIn_1 == 1'h0; // @[Controllers.scala 135:105:@472.4]
  assign _T_179 = _T_176 & _T_178; // @[Controllers.scala 135:103:@473.4]
  assign _T_180 = _T_179 & io_enable; // @[Controllers.scala 135:119:@474.4]
  assign _T_182 = io_doneIn_0 | _T_180; // @[Controllers.scala 135:51:@476.4]
  assign _T_205 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@501.4]
  assign _T_207 = _T_205 & _T_150; // @[Controllers.scala 213:90:@503.4]
  assign _T_209 = ~ allDone; // @[Controllers.scala 213:132:@505.4]
  assign _T_210 = _T_207 & _T_209; // @[Controllers.scala 213:130:@506.4]
  assign _T_211 = ~ io_ctrDone; // @[Controllers.scala 213:156:@507.4]
  assign _T_213 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@510.4]
  assign _T_215 = _T_213 & _T_175; // @[Controllers.scala 213:90:@512.4]
  assign _T_222 = allDone == 1'h0; // @[package.scala 100:49:@518.4]
  assign io_done = RetimeWrapper_2_io_out; // @[Controllers.scala 245:13:@547.4]
  assign io_ctrInc = io_doneIn_1; // @[Controllers.scala 122:17:@426.4]
  assign io_enableOut_0 = _T_210 & _T_211; // @[Controllers.scala 213:55:@509.4]
  assign io_enableOut_1 = _T_215 & _T_209; // @[Controllers.scala 213:55:@517.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@498.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@500.4]
  assign active_0_clock = clock; // @[:@358.4]
  assign active_0_reset = reset; // @[:@359.4]
  assign active_0_io_input_set = _T_151 & _T_153; // @[Controllers.scala 128:30:@450.4]
  assign active_0_io_input_reset = _T_155 | allDone; // @[Controllers.scala 129:32:@455.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@372.4]
  assign active_1_clock = clock; // @[:@361.4]
  assign active_1_reset = reset; // @[:@362.4]
  assign active_1_io_input_set = _T_182 & _T_160; // @[Controllers.scala 135:32:@479.4]
  assign active_1_io_input_reset = io_doneIn_1 | io_rst; // @[Controllers.scala 136:34:@483.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@373.4]
  assign done_0_clock = clock; // @[:@364.4]
  assign done_0_reset = reset; // @[:@365.4]
  assign done_0_io_input_set = io_ctrDone & _T_172; // @[Controllers.scala 131:28:@469.4]
  assign done_0_io_input_reset = io_rst | allDone; // @[Controllers.scala 86:33:@384.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@374.4]
  assign done_1_clock = clock; // @[:@367.4]
  assign done_1_reset = reset; // @[:@368.4]
  assign done_1_io_input_set = io_ctrDone & _T_172; // @[Controllers.scala 138:30:@496.4]
  assign done_1_io_input_reset = io_rst | allDone; // @[Controllers.scala 86:33:@393.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@375.4]
  assign iterDone_0_clock = clock; // @[:@396.4]
  assign iterDone_0_reset = reset; // @[:@397.4]
  assign iterDone_0_io_input_set = _T_161 & _T_169; // @[Controllers.scala 130:32:@465.4]
  assign iterDone_0_io_input_reset = synchronize | io_rst; // @[Controllers.scala 92:37:@411.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@401.4]
  assign iterDone_1_clock = clock; // @[:@399.4]
  assign iterDone_1_reset = reset; // @[:@400.4]
  assign iterDone_1_io_input_set = io_doneIn_1 & _T_160; // @[Controllers.scala 137:34:@492.4]
  assign iterDone_1_io_input_reset = synchronize | io_rst; // @[Controllers.scala 92:37:@420.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@402.4]
  assign RetimeWrapper_clock = clock; // @[:@428.4]
  assign RetimeWrapper_reset = reset; // @[:@429.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@431.4]
  assign RetimeWrapper_io_in = io_doneIn_1; // @[package.scala 94:16:@430.4]
  assign RetimeWrapper_1_clock = clock; // @[:@524.4]
  assign RetimeWrapper_1_reset = reset; // @[:@525.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@527.4]
  assign RetimeWrapper_1_io_in = allDone & _T_225; // @[package.scala 94:16:@526.4]
  assign RetimeWrapper_2_clock = clock; // @[:@541.4]
  assign RetimeWrapper_2_reset = reset; // @[:@542.4]
  assign RetimeWrapper_2_io_flow = io_enable; // @[package.scala 95:18:@544.4]
  assign RetimeWrapper_2_io_in = allDone & _T_239; // @[package.scala 94:16:@543.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_225 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_239 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_225 <= 1'h0;
    end else begin
      _T_225 <= _T_222;
    end
    if (reset) begin
      _T_239 <= 1'h0;
    end else begin
      _T_239 <= _T_222;
    end
  end
endmodule
module SRAM( // @[:@613.2]
  input         clock, // @[:@614.4]
  input         reset, // @[:@615.4]
  input  [8:0]  io_raddr, // @[:@616.4]
  input         io_wen, // @[:@616.4]
  input  [8:0]  io_waddr, // @[:@616.4]
  input  [31:0] io_wdata, // @[:@616.4]
  output [31:0] io_rdata, // @[:@616.4]
  input         io_backpressure // @[:@616.4]
);
  wire [31:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 124:30:@618.4]
  wire [31:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 124:30:@618.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 124:30:@618.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 124:30:@618.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 124:30:@618.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 124:30:@618.4]
  wire [8:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 124:30:@618.4]
  wire [8:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 124:30:@618.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 124:30:@618.4]
  wire  _T_19; // @[SRAM.scala 137:49:@636.4]
  wire  _T_20; // @[SRAM.scala 137:37:@637.4]
  reg  _T_23; // @[SRAM.scala 137:29:@638.4]
  reg [31:0] _RAND_0;
  reg [31:0] _T_26; // @[SRAM.scala 138:29:@640.4]
  reg [31:0] _RAND_1;
  SRAMVerilogAWS #(.DWIDTH(32), .WORDS(384), .AWIDTH(9)) SRAMVerilogAWS ( // @[SRAM.scala 124:30:@618.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_19 = io_raddr == io_waddr; // @[SRAM.scala 137:49:@636.4]
  assign _T_20 = io_wen & _T_19; // @[SRAM.scala 137:37:@637.4]
  assign io_rdata = _T_23 ? _T_26 : SRAMVerilogAWS_rdata; // @[SRAM.scala 139:16:@645.4]
  assign SRAMVerilogAWS_wdata = io_wdata; // @[SRAM.scala 130:20:@632.4]
  assign SRAMVerilogAWS_backpressure = io_backpressure; // @[SRAM.scala 131:27:@633.4]
  assign SRAMVerilogAWS_wen = io_wen; // @[SRAM.scala 128:18:@630.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 133:22:@635.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 132:22:@634.4]
  assign SRAMVerilogAWS_waddr = io_waddr; // @[SRAM.scala 129:20:@631.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 127:20:@629.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 126:18:@628.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_23 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_26 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_23 <= 1'h0;
    end else begin
      _T_23 <= _T_20;
    end
    if (reset) begin
      _T_26 <= 32'h0;
    end else begin
      _T_26 <= io_wdata;
    end
  end
endmodule
module RetimeWrapper_5( // @[:@659.2]
  input        clock, // @[:@660.4]
  input        reset, // @[:@661.4]
  input        io_flow, // @[:@662.4]
  input  [8:0] io_in, // @[:@662.4]
  output [8:0] io_out // @[:@662.4]
);
  wire [8:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@664.4]
  wire [8:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@664.4]
  wire [8:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@664.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@664.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@664.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@664.4]
  RetimeShiftRegister #(.WIDTH(9), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@664.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@677.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@676.4]
  assign sr_init = 9'h0; // @[RetimeShiftRegister.scala 19:16:@675.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@674.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@673.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@671.4]
endmodule
module Mem1D( // @[:@679.2]
  input         clock, // @[:@680.4]
  input         reset, // @[:@681.4]
  input  [8:0]  io_r_ofs_0, // @[:@682.4]
  input         io_r_backpressure, // @[:@682.4]
  input  [8:0]  io_w_ofs_0, // @[:@682.4]
  input  [31:0] io_w_data_0, // @[:@682.4]
  input         io_w_en_0, // @[:@682.4]
  output [31:0] io_output // @[:@682.4]
);
  wire  SRAM_clock; // @[MemPrimitives.scala 567:21:@686.4]
  wire  SRAM_reset; // @[MemPrimitives.scala 567:21:@686.4]
  wire [8:0] SRAM_io_raddr; // @[MemPrimitives.scala 567:21:@686.4]
  wire  SRAM_io_wen; // @[MemPrimitives.scala 567:21:@686.4]
  wire [8:0] SRAM_io_waddr; // @[MemPrimitives.scala 567:21:@686.4]
  wire [31:0] SRAM_io_wdata; // @[MemPrimitives.scala 567:21:@686.4]
  wire [31:0] SRAM_io_rdata; // @[MemPrimitives.scala 567:21:@686.4]
  wire  SRAM_io_backpressure; // @[MemPrimitives.scala 567:21:@686.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@689.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@689.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@689.4]
  wire [8:0] RetimeWrapper_io_in; // @[package.scala 93:22:@689.4]
  wire [8:0] RetimeWrapper_io_out; // @[package.scala 93:22:@689.4]
  wire  wInBound; // @[MemPrimitives.scala 554:32:@684.4]
  SRAM SRAM ( // @[MemPrimitives.scala 567:21:@686.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata(SRAM_io_wdata),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  RetimeWrapper_5 RetimeWrapper ( // @[package.scala 93:22:@689.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign wInBound = io_w_ofs_0 <= 9'h180; // @[MemPrimitives.scala 554:32:@684.4]
  assign io_output = SRAM_io_rdata; // @[MemPrimitives.scala 574:17:@702.4]
  assign SRAM_clock = clock; // @[:@687.4]
  assign SRAM_reset = reset; // @[:@688.4]
  assign SRAM_io_raddr = RetimeWrapper_io_out; // @[MemPrimitives.scala 568:37:@696.4]
  assign SRAM_io_wen = io_w_en_0 & wInBound; // @[MemPrimitives.scala 571:22:@699.4]
  assign SRAM_io_waddr = io_w_ofs_0; // @[MemPrimitives.scala 570:22:@697.4]
  assign SRAM_io_wdata = io_w_data_0; // @[MemPrimitives.scala 572:22:@700.4]
  assign SRAM_io_backpressure = io_r_backpressure; // @[MemPrimitives.scala 573:30:@701.4]
  assign RetimeWrapper_clock = clock; // @[:@690.4]
  assign RetimeWrapper_reset = reset; // @[:@691.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@693.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@692.4]
endmodule
module StickySelects( // @[:@704.2]
  input   io_ins_0, // @[:@707.4]
  output  io_outs_0 // @[:@707.4]
);
  assign io_outs_0 = io_ins_0; // @[StickySelects.scala 12:26:@709.4]
endmodule
module x43_mem_0( // @[:@711.2]
  input         clock, // @[:@712.4]
  input         reset, // @[:@713.4]
  input         io_rPort_0_en_0, // @[:@714.4]
  output [31:0] io_rPort_0_output_0, // @[:@714.4]
  input  [8:0]  io_wPort_0_ofs_0, // @[:@714.4]
  input  [31:0] io_wPort_0_data_0, // @[:@714.4]
  input         io_wPort_0_en_0 // @[:@714.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@729.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@729.4]
  wire [8:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@729.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@729.4]
  wire [8:0] Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@729.4]
  wire [31:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@729.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@729.4]
  wire [31:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@729.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 121:29:@755.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 121:29:@755.4]
  wire [41:0] _T_70; // @[Cat.scala 30:58:@747.4]
  wire  _T_76; // @[MemPrimitives.scala 123:41:@759.4]
  wire [10:0] _T_78; // @[Cat.scala 30:58:@761.4]
  Mem1D Mem1D ( // @[MemPrimitives.scala 64:21:@729.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  StickySelects StickySelects ( // @[MemPrimitives.scala 121:29:@755.4]
    .io_ins_0(StickySelects_io_ins_0),
    .io_outs_0(StickySelects_io_outs_0)
  );
  assign _T_70 = {io_wPort_0_en_0,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@747.4]
  assign _T_76 = StickySelects_io_outs_0; // @[MemPrimitives.scala 123:41:@759.4]
  assign _T_78 = {_T_76,1'h1,9'h17f}; // @[Cat.scala 30:58:@761.4]
  assign io_rPort_0_output_0 = Mem1D_io_output; // @[MemPrimitives.scala 148:13:@769.4]
  assign Mem1D_clock = clock; // @[:@730.4]
  assign Mem1D_reset = reset; // @[:@731.4]
  assign Mem1D_io_r_ofs_0 = _T_78[8:0]; // @[MemPrimitives.scala 127:28:@765.4]
  assign Mem1D_io_r_backpressure = _T_78[9]; // @[MemPrimitives.scala 128:32:@766.4]
  assign Mem1D_io_w_ofs_0 = _T_70[8:0]; // @[MemPrimitives.scala 94:28:@751.4]
  assign Mem1D_io_w_data_0 = _T_70[40:9]; // @[MemPrimitives.scala 95:29:@752.4]
  assign Mem1D_io_w_en_0 = _T_70[41]; // @[MemPrimitives.scala 96:27:@753.4]
  assign StickySelects_io_ins_0 = io_rPort_0_en_0; // @[MemPrimitives.scala 122:60:@758.4]
endmodule
module SingleCounter_1( // @[:@809.2]
  input         clock, // @[:@810.4]
  input         reset, // @[:@811.4]
  input         io_input_reset, // @[:@812.4]
  input         io_input_enable, // @[:@812.4]
  output [31:0] io_output_count_0, // @[:@812.4]
  output        io_output_oobs_0, // @[:@812.4]
  output        io_output_done // @[:@812.4]
);
  wire  bases_0_clock; // @[Counter.scala 253:53:@825.4]
  wire  bases_0_reset; // @[Counter.scala 253:53:@825.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 253:53:@825.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 253:53:@825.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 253:53:@825.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 253:53:@825.4]
  wire  SRFF_clock; // @[Counter.scala 255:22:@841.4]
  wire  SRFF_reset; // @[Counter.scala 255:22:@841.4]
  wire  SRFF_io_input_set; // @[Counter.scala 255:22:@841.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 255:22:@841.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 255:22:@841.4]
  wire  SRFF_io_output; // @[Counter.scala 255:22:@841.4]
  wire  _T_36; // @[Counter.scala 256:45:@844.4]
  wire [31:0] _T_48; // @[Counter.scala 279:52:@869.4]
  wire [32:0] _T_50; // @[Counter.scala 283:33:@870.4]
  wire [31:0] _T_51; // @[Counter.scala 283:33:@871.4]
  wire [31:0] _T_52; // @[Counter.scala 283:33:@872.4]
  wire  _T_57; // @[Counter.scala 285:18:@874.4]
  wire [31:0] _T_68; // @[Counter.scala 291:115:@882.4]
  wire [31:0] _T_71; // @[Counter.scala 291:152:@885.4]
  wire [31:0] _T_72; // @[Counter.scala 291:74:@886.4]
  wire  _T_75; // @[Counter.scala 314:102:@890.4]
  wire  _T_77; // @[Counter.scala 314:130:@891.4]
  FF bases_0 ( // @[Counter.scala 253:53:@825.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 255:22:@841.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 256:45:@844.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 279:52:@869.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@870.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@871.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 283:33:@872.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh180); // @[Counter.scala 285:18:@874.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 291:115:@882.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 291:152:@885.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 291:74:@886.4]
  assign _T_75 = $signed(_T_48) < $signed(32'sh0); // @[Counter.scala 314:102:@890.4]
  assign _T_77 = $signed(_T_48) >= $signed(32'sh180); // @[Counter.scala 314:130:@891.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 296:28:@889.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 314:60:@893.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 325:20:@895.4]
  assign bases_0_clock = clock; // @[:@826.4]
  assign bases_0_reset = reset; // @[:@827.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 291:31:@888.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 273:27:@867.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 276:29:@868.4]
  assign SRFF_clock = clock; // @[:@842.4]
  assign SRFF_reset = reset; // @[:@843.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 256:23:@846.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 257:25:@848.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 258:30:@849.4]
endmodule
module x45_ctrchain( // @[:@900.2]
  input         clock, // @[:@901.4]
  input         reset, // @[:@902.4]
  input         io_input_reset, // @[:@903.4]
  input         io_input_enable, // @[:@903.4]
  output [31:0] io_output_counts_0, // @[:@903.4]
  output        io_output_oobs_0, // @[:@903.4]
  output        io_output_done // @[:@903.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 505:46:@905.4]
  wire  ctrs_0_reset; // @[Counter.scala 505:46:@905.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 505:46:@905.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 505:46:@905.4]
  wire [31:0] ctrs_0_io_output_count_0; // @[Counter.scala 505:46:@905.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 505:46:@905.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 505:46:@905.4]
  reg  wasDone; // @[Counter.scala 534:24:@914.4]
  reg [31:0] _RAND_0;
  wire  _T_45; // @[Counter.scala 538:69:@920.4]
  wire  _T_47; // @[Counter.scala 538:80:@921.4]
  reg  doneLatch; // @[Counter.scala 542:26:@926.4]
  reg [31:0] _RAND_1;
  wire  _T_54; // @[Counter.scala 543:48:@927.4]
  wire  _T_55; // @[Counter.scala 543:19:@928.4]
  SingleCounter_1 ctrs_0 ( // @[Counter.scala 505:46:@905.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done)
  );
  assign _T_45 = io_input_enable & ctrs_0_io_output_done; // @[Counter.scala 538:69:@920.4]
  assign _T_47 = wasDone == 1'h0; // @[Counter.scala 538:80:@921.4]
  assign _T_54 = ctrs_0_io_output_done ? 1'h1 : doneLatch; // @[Counter.scala 543:48:@927.4]
  assign _T_55 = io_input_reset ? 1'h0 : _T_54; // @[Counter.scala 543:19:@928.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 549:32:@930.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 550:30:@932.4]
  assign io_output_done = _T_45 & _T_47; // @[Counter.scala 538:18:@923.4]
  assign ctrs_0_clock = clock; // @[:@906.4]
  assign ctrs_0_reset = reset; // @[:@907.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 512:24:@911.4]
  assign ctrs_0_io_input_enable = io_input_enable; // @[Counter.scala 516:33:@912.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= ctrs_0_io_output_done;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (ctrs_0_io_output_done) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module x53_inr_Foreach_sm( // @[:@1024.2]
  input   clock, // @[:@1025.4]
  input   reset, // @[:@1026.4]
  input   io_enable, // @[:@1027.4]
  output  io_done, // @[:@1027.4]
  input   io_ctrDone, // @[:@1027.4]
  output  io_datapathEn, // @[:@1027.4]
  output  io_ctrInc, // @[:@1027.4]
  output  io_ctrRst, // @[:@1027.4]
  input   io_parentAck, // @[:@1027.4]
  input   io_break // @[:@1027.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@1029.4]
  wire  active_reset; // @[Controllers.scala 261:22:@1029.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@1029.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@1029.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@1029.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@1029.4]
  wire  done_clock; // @[Controllers.scala 262:20:@1032.4]
  wire  done_reset; // @[Controllers.scala 262:20:@1032.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@1032.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@1032.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@1032.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@1032.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@1086.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@1086.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@1086.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@1086.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@1086.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@1094.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@1094.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@1094.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@1094.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@1094.4]
  wire  _T_80; // @[Controllers.scala 264:48:@1037.4]
  wire  _T_81; // @[Controllers.scala 264:46:@1038.4]
  wire  _T_82; // @[Controllers.scala 264:62:@1039.4]
  wire  _T_100; // @[package.scala 100:49:@1057.4]
  reg  _T_103; // @[package.scala 48:56:@1058.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 100:49:@1066.4]
  reg  _T_111; // @[package.scala 48:56:@1067.4]
  reg [31:0] _RAND_1;
  wire  _T_112; // @[package.scala 100:41:@1069.4]
  wire  _T_116; // @[Controllers.scala 283:41:@1074.4]
  reg  _T_125; // @[package.scala 48:56:@1082.4]
  reg [31:0] _RAND_2;
  SRFF active ( // @[Controllers.scala 261:22:@1029.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@1032.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@1086.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@1094.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@1037.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@1038.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@1039.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@1057.4]
  assign _T_108 = done_io_output == 1'h0; // @[package.scala 100:49:@1066.4]
  assign _T_112 = done_io_output & _T_111; // @[package.scala 100:41:@1069.4]
  assign _T_116 = active_io_output & _T_82; // @[Controllers.scala 283:41:@1074.4]
  assign io_done = done_io_output & _T_125; // @[Controllers.scala 287:13:@1085.4]
  assign io_datapathEn = _T_116 & io_enable; // @[Controllers.scala 283:21:@1077.4]
  assign io_ctrInc = active_io_output & io_enable; // @[Controllers.scala 284:17:@1080.4]
  assign io_ctrRst = _T_112 | io_parentAck; // @[Controllers.scala 274:13:@1072.4]
  assign active_clock = clock; // @[:@1030.4]
  assign active_reset = reset; // @[:@1031.4]
  assign active_io_input_set = _T_81 & _T_82; // @[Controllers.scala 264:23:@1042.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@1046.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@1047.4]
  assign done_clock = clock; // @[:@1033.4]
  assign done_reset = reset; // @[:@1034.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@1062.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@1055.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@1056.4]
  assign RetimeWrapper_clock = clock; // @[:@1087.4]
  assign RetimeWrapper_reset = reset; // @[:@1088.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@1090.4]
  assign RetimeWrapper_io_in = 1'h0; // @[package.scala 94:16:@1089.4]
  assign RetimeWrapper_1_clock = clock; // @[:@1095.4]
  assign RetimeWrapper_1_reset = reset; // @[:@1096.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@1098.4]
  assign RetimeWrapper_1_io_in = io_ctrDone; // @[package.scala 94:16:@1097.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_111 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_125 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_111 <= 1'h0;
    end else begin
      _T_111 <= _T_108;
    end
    if (reset) begin
      _T_125 <= 1'h0;
    end else begin
      _T_125 <= _T_108;
    end
  end
endmodule
module fix2fixBox( // @[:@1219.2]
  input  [31:0] io_a, // @[:@1222.4]
  output [31:0] io_b // @[:@1222.4]
);
  assign io_b = io_a; // @[Converter.scala 95:38:@1232.4]
endmodule
module _( // @[:@1234.2]
  input  [31:0] io_b, // @[:@1237.4]
  output [31:0] io_result // @[:@1237.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@1242.4]
  wire [31:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@1242.4]
  fix2fixBox fix2fixBox ( // @[BigIPZynq.scala 219:30:@1242.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 706:17:@1250.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@1245.4]
endmodule
module fix2fixBox_1( // @[:@1252.2]
  input  [31:0] io_a, // @[:@1255.4]
  output [32:0] io_b // @[:@1255.4]
);
  wire  _T_20; // @[implicits.scala 69:16:@1262.4]
  assign _T_20 = io_a[31]; // @[implicits.scala 69:16:@1262.4]
  assign io_b = {_T_20,io_a}; // @[Converter.scala 95:38:@1267.4]
endmodule
module __1( // @[:@1269.2]
  input  [31:0] io_b, // @[:@1272.4]
  output [32:0] io_result // @[:@1272.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@1277.4]
  wire [32:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@1277.4]
  fix2fixBox_1 fix2fixBox ( // @[BigIPZynq.scala 219:30:@1277.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 706:17:@1285.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@1280.4]
endmodule
module fix2fixBox_3( // @[:@1322.2]
  input  [32:0] io_a, // @[:@1325.4]
  output [31:0] io_b // @[:@1325.4]
);
  assign io_b = io_a[31:0]; // @[Converter.scala 95:38:@1335.4]
endmodule
module x49_sum( // @[:@1337.2]
  input  [31:0] io_a, // @[:@1340.4]
  input  [31:0] io_b, // @[:@1340.4]
  output [31:0] io_result // @[:@1340.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@1348.4]
  wire [32:0] __io_result; // @[Math.scala 709:24:@1348.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@1355.4]
  wire [32:0] __1_io_result; // @[Math.scala 709:24:@1355.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@1373.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@1373.4]
  wire [32:0] a_upcast_number; // @[Math.scala 712:22:@1353.4 Math.scala 713:14:@1354.4]
  wire [32:0] b_upcast_number; // @[Math.scala 712:22:@1360.4 Math.scala 713:14:@1361.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@1362.4]
  __1 _ ( // @[Math.scala 709:24:@1348.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __1 __1 ( // @[Math.scala 709:24:@1355.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_3 fix2fixBox ( // @[Math.scala 141:30:@1373.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@1353.4 Math.scala 713:14:@1354.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@1360.4 Math.scala 713:14:@1361.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@1362.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@1381.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@1351.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@1358.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@1376.4]
endmodule
module x53_inr_Foreach_kernelx53_inr_Foreach_concrete1( // @[:@1383.2]
  input  [63:0] io_in_x38_x, // @[:@1386.4]
  output [8:0]  io_in_x43_mem_0_wPort_0_ofs_0, // @[:@1386.4]
  output [31:0] io_in_x43_mem_0_wPort_0_data_0, // @[:@1386.4]
  output        io_in_x43_mem_0_wPort_0_en_0, // @[:@1386.4]
  input         io_sigsIn_datapathEn, // @[:@1386.4]
  input         io_sigsIn_break, // @[:@1386.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@1386.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@1386.4]
  input         io_rr // @[:@1386.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@1413.4]
  wire [31:0] __io_result; // @[Math.scala 709:24:@1413.4]
  wire [31:0] x49_sum_1_io_a; // @[Math.scala 150:24:@1425.4]
  wire [31:0] x49_sum_1_io_b; // @[Math.scala 150:24:@1425.4]
  wire [31:0] x49_sum_1_io_result; // @[Math.scala 150:24:@1425.4]
  wire  b47; // @[sm_x53_inr_Foreach.scala 61:17:@1421.4]
  wire  _T_261; // @[sm_x53_inr_Foreach.scala 70:92:@1436.4]
  wire  _T_265; // @[implicits.scala 55:10:@1439.4]
  wire  _T_266; // @[sm_x53_inr_Foreach.scala 70:109:@1440.4]
  wire  _T_268; // @[sm_x53_inr_Foreach.scala 70:196:@1442.4]
  wire [31:0] b46_number; // @[Math.scala 712:22:@1418.4 Math.scala 713:14:@1419.4]
  _ _ ( // @[Math.scala 709:24:@1413.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  x49_sum x49_sum_1 ( // @[Math.scala 150:24:@1425.4]
    .io_a(x49_sum_1_io_a),
    .io_b(x49_sum_1_io_b),
    .io_result(x49_sum_1_io_result)
  );
  assign b47 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x53_inr_Foreach.scala 61:17:@1421.4]
  assign _T_261 = ~ io_sigsIn_break; // @[sm_x53_inr_Foreach.scala 70:92:@1436.4]
  assign _T_265 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 55:10:@1439.4]
  assign _T_266 = _T_261 & _T_265; // @[sm_x53_inr_Foreach.scala 70:109:@1440.4]
  assign _T_268 = _T_266 & _T_261; // @[sm_x53_inr_Foreach.scala 70:196:@1442.4]
  assign b46_number = __io_result; // @[Math.scala 712:22:@1418.4 Math.scala 713:14:@1419.4]
  assign io_in_x43_mem_0_wPort_0_ofs_0 = b46_number[8:0]; // @[MemInterfaceType.scala 89:54:@1446.4]
  assign io_in_x43_mem_0_wPort_0_data_0 = x49_sum_1_io_result; // @[MemInterfaceType.scala 90:56:@1447.4]
  assign io_in_x43_mem_0_wPort_0_en_0 = _T_268 & b47; // @[MemInterfaceType.scala 93:57:@1449.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 710:17:@1416.4]
  assign x49_sum_1_io_a = io_in_x38_x[31:0]; // @[Math.scala 151:17:@1428.4]
  assign x49_sum_1_io_b = __io_result; // @[Math.scala 152:17:@1429.4]
endmodule
module x57_inr_UnitPipe_kernelx57_inr_UnitPipe_concrete1( // @[:@1704.2]
  output        io_in_x43_mem_0_rPort_0_en_0, // @[:@1707.4]
  input  [31:0] io_in_x43_mem_0_rPort_0_output_0, // @[:@1707.4]
  output        io_in_x39_y_port_0_valid, // @[:@1707.4]
  output [63:0] io_in_x39_y_port_0_bits, // @[:@1707.4]
  input         io_sigsIn_datapathEn, // @[:@1707.4]
  input         io_sigsIn_break, // @[:@1707.4]
  input         io_rr // @[:@1707.4]
);
  wire  _T_277; // @[sm_x57_inr_UnitPipe.scala 65:120:@1739.4]
  wire  _T_281; // @[implicits.scala 55:10:@1742.4]
  wire  _T_286; // @[FixedPoint.scala 50:25:@1752.4]
  wire [31:0] _T_290; // @[Bitwise.scala 72:12:@1754.4]
  assign _T_277 = ~ io_sigsIn_break; // @[sm_x57_inr_UnitPipe.scala 65:120:@1739.4]
  assign _T_281 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 55:10:@1742.4]
  assign _T_286 = io_in_x43_mem_0_rPort_0_output_0[31]; // @[FixedPoint.scala 50:25:@1752.4]
  assign _T_290 = _T_286 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12:@1754.4]
  assign io_in_x43_mem_0_rPort_0_en_0 = _T_277 & _T_281; // @[MemInterfaceType.scala 110:79:@1748.4]
  assign io_in_x39_y_port_0_valid = io_sigsIn_datapathEn; // @[MemInterfaceType.scala 311:132:@1759.4]
  assign io_in_x39_y_port_0_bits = {_T_290,io_in_x43_mem_0_rPort_0_output_0}; // @[MemInterfaceType.scala 311:109:@1758.4]
endmodule
module RootController_kernelRootController_concrete1( // @[:@1761.2]
  input         clock, // @[:@1762.4]
  input         reset, // @[:@1763.4]
  input  [63:0] io_in_x38_x, // @[:@1764.4]
  output        io_in_x39_y_port_0_valid, // @[:@1764.4]
  output [63:0] io_in_x39_y_port_0_bits, // @[:@1764.4]
  input         io_sigsIn_smEnableOuts_0, // @[:@1764.4]
  input         io_sigsIn_smEnableOuts_1, // @[:@1764.4]
  input         io_sigsIn_smChildAcks_0, // @[:@1764.4]
  input         io_sigsIn_smChildAcks_1, // @[:@1764.4]
  output        io_sigsOut_smDoneIn_0, // @[:@1764.4]
  output        io_sigsOut_smDoneIn_1, // @[:@1764.4]
  input         io_rr // @[:@1764.4]
);
  wire  x43_mem_0_clock; // @[m_x43_mem_0.scala 26:17:@1780.4]
  wire  x43_mem_0_reset; // @[m_x43_mem_0.scala 26:17:@1780.4]
  wire  x43_mem_0_io_rPort_0_en_0; // @[m_x43_mem_0.scala 26:17:@1780.4]
  wire [31:0] x43_mem_0_io_rPort_0_output_0; // @[m_x43_mem_0.scala 26:17:@1780.4]
  wire [8:0] x43_mem_0_io_wPort_0_ofs_0; // @[m_x43_mem_0.scala 26:17:@1780.4]
  wire [31:0] x43_mem_0_io_wPort_0_data_0; // @[m_x43_mem_0.scala 26:17:@1780.4]
  wire  x43_mem_0_io_wPort_0_en_0; // @[m_x43_mem_0.scala 26:17:@1780.4]
  wire  x45_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@1797.4]
  wire  x45_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@1797.4]
  wire  x45_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@1797.4]
  wire  x45_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@1797.4]
  wire [31:0] x45_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@1797.4]
  wire  x45_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@1797.4]
  wire  x45_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@1797.4]
  wire  x53_inr_Foreach_sm_clock; // @[sm_x53_inr_Foreach.scala 32:18:@1849.4]
  wire  x53_inr_Foreach_sm_reset; // @[sm_x53_inr_Foreach.scala 32:18:@1849.4]
  wire  x53_inr_Foreach_sm_io_enable; // @[sm_x53_inr_Foreach.scala 32:18:@1849.4]
  wire  x53_inr_Foreach_sm_io_done; // @[sm_x53_inr_Foreach.scala 32:18:@1849.4]
  wire  x53_inr_Foreach_sm_io_ctrDone; // @[sm_x53_inr_Foreach.scala 32:18:@1849.4]
  wire  x53_inr_Foreach_sm_io_datapathEn; // @[sm_x53_inr_Foreach.scala 32:18:@1849.4]
  wire  x53_inr_Foreach_sm_io_ctrInc; // @[sm_x53_inr_Foreach.scala 32:18:@1849.4]
  wire  x53_inr_Foreach_sm_io_ctrRst; // @[sm_x53_inr_Foreach.scala 32:18:@1849.4]
  wire  x53_inr_Foreach_sm_io_parentAck; // @[sm_x53_inr_Foreach.scala 32:18:@1849.4]
  wire  x53_inr_Foreach_sm_io_break; // @[sm_x53_inr_Foreach.scala 32:18:@1849.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@1877.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@1877.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@1877.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@1877.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@1877.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@1917.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@1917.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@1917.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@1917.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@1917.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@1925.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@1925.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@1925.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@1925.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@1925.4]
  wire [63:0] x53_inr_Foreach_kernelx53_inr_Foreach_concrete1_io_in_x38_x; // @[sm_x53_inr_Foreach.scala 72:24:@1956.4]
  wire [8:0] x53_inr_Foreach_kernelx53_inr_Foreach_concrete1_io_in_x43_mem_0_wPort_0_ofs_0; // @[sm_x53_inr_Foreach.scala 72:24:@1956.4]
  wire [31:0] x53_inr_Foreach_kernelx53_inr_Foreach_concrete1_io_in_x43_mem_0_wPort_0_data_0; // @[sm_x53_inr_Foreach.scala 72:24:@1956.4]
  wire  x53_inr_Foreach_kernelx53_inr_Foreach_concrete1_io_in_x43_mem_0_wPort_0_en_0; // @[sm_x53_inr_Foreach.scala 72:24:@1956.4]
  wire  x53_inr_Foreach_kernelx53_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x53_inr_Foreach.scala 72:24:@1956.4]
  wire  x53_inr_Foreach_kernelx53_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x53_inr_Foreach.scala 72:24:@1956.4]
  wire [31:0] x53_inr_Foreach_kernelx53_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x53_inr_Foreach.scala 72:24:@1956.4]
  wire  x53_inr_Foreach_kernelx53_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x53_inr_Foreach.scala 72:24:@1956.4]
  wire  x53_inr_Foreach_kernelx53_inr_Foreach_concrete1_io_rr; // @[sm_x53_inr_Foreach.scala 72:24:@1956.4]
  wire  x57_inr_UnitPipe_sm_clock; // @[sm_x57_inr_UnitPipe.scala 32:18:@2069.4]
  wire  x57_inr_UnitPipe_sm_reset; // @[sm_x57_inr_UnitPipe.scala 32:18:@2069.4]
  wire  x57_inr_UnitPipe_sm_io_enable; // @[sm_x57_inr_UnitPipe.scala 32:18:@2069.4]
  wire  x57_inr_UnitPipe_sm_io_done; // @[sm_x57_inr_UnitPipe.scala 32:18:@2069.4]
  wire  x57_inr_UnitPipe_sm_io_ctrDone; // @[sm_x57_inr_UnitPipe.scala 32:18:@2069.4]
  wire  x57_inr_UnitPipe_sm_io_datapathEn; // @[sm_x57_inr_UnitPipe.scala 32:18:@2069.4]
  wire  x57_inr_UnitPipe_sm_io_ctrInc; // @[sm_x57_inr_UnitPipe.scala 32:18:@2069.4]
  wire  x57_inr_UnitPipe_sm_io_ctrRst; // @[sm_x57_inr_UnitPipe.scala 32:18:@2069.4]
  wire  x57_inr_UnitPipe_sm_io_parentAck; // @[sm_x57_inr_UnitPipe.scala 32:18:@2069.4]
  wire  x57_inr_UnitPipe_sm_io_break; // @[sm_x57_inr_UnitPipe.scala 32:18:@2069.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@2126.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@2126.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@2126.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@2126.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@2126.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@2134.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@2134.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@2134.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@2134.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@2134.4]
  wire  x57_inr_UnitPipe_kernelx57_inr_UnitPipe_concrete1_io_in_x43_mem_0_rPort_0_en_0; // @[sm_x57_inr_UnitPipe.scala 70:24:@2160.4]
  wire [31:0] x57_inr_UnitPipe_kernelx57_inr_UnitPipe_concrete1_io_in_x43_mem_0_rPort_0_output_0; // @[sm_x57_inr_UnitPipe.scala 70:24:@2160.4]
  wire  x57_inr_UnitPipe_kernelx57_inr_UnitPipe_concrete1_io_in_x39_y_port_0_valid; // @[sm_x57_inr_UnitPipe.scala 70:24:@2160.4]
  wire [63:0] x57_inr_UnitPipe_kernelx57_inr_UnitPipe_concrete1_io_in_x39_y_port_0_bits; // @[sm_x57_inr_UnitPipe.scala 70:24:@2160.4]
  wire  x57_inr_UnitPipe_kernelx57_inr_UnitPipe_concrete1_io_sigsIn_datapathEn; // @[sm_x57_inr_UnitPipe.scala 70:24:@2160.4]
  wire  x57_inr_UnitPipe_kernelx57_inr_UnitPipe_concrete1_io_sigsIn_break; // @[sm_x57_inr_UnitPipe.scala 70:24:@2160.4]
  wire  x57_inr_UnitPipe_kernelx57_inr_UnitPipe_concrete1_io_rr; // @[sm_x57_inr_UnitPipe.scala 70:24:@2160.4]
  wire  _T_200; // @[package.scala 96:25:@1882.4 package.scala 96:25:@1883.4]
  wire  _T_215; // @[package.scala 96:25:@1922.4 package.scala 96:25:@1923.4]
  wire  _T_221; // @[package.scala 96:25:@1930.4 package.scala 96:25:@1931.4]
  wire  _T_224; // @[SpatialBlocks.scala 110:93:@1933.4]
  wire  _T_226; // @[SpatialBlocks.scala 128:36:@1942.4]
  wire  _T_227; // @[SpatialBlocks.scala 128:78:@1943.4]
  wire  _T_292; // @[package.scala 100:49:@2097.4]
  reg  _T_295; // @[package.scala 48:56:@2098.4]
  reg [31:0] _RAND_0;
  wire  _T_309; // @[package.scala 96:25:@2131.4 package.scala 96:25:@2132.4]
  wire  _T_315; // @[package.scala 96:25:@2139.4 package.scala 96:25:@2140.4]
  wire  _T_318; // @[SpatialBlocks.scala 110:93:@2142.4]
  x43_mem_0 x43_mem_0 ( // @[m_x43_mem_0.scala 26:17:@1780.4]
    .clock(x43_mem_0_clock),
    .reset(x43_mem_0_reset),
    .io_rPort_0_en_0(x43_mem_0_io_rPort_0_en_0),
    .io_rPort_0_output_0(x43_mem_0_io_rPort_0_output_0),
    .io_wPort_0_ofs_0(x43_mem_0_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x43_mem_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x43_mem_0_io_wPort_0_en_0)
  );
  x45_ctrchain x45_ctrchain ( // @[SpatialBlocks.scala 37:22:@1797.4]
    .clock(x45_ctrchain_clock),
    .reset(x45_ctrchain_reset),
    .io_input_reset(x45_ctrchain_io_input_reset),
    .io_input_enable(x45_ctrchain_io_input_enable),
    .io_output_counts_0(x45_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x45_ctrchain_io_output_oobs_0),
    .io_output_done(x45_ctrchain_io_output_done)
  );
  x53_inr_Foreach_sm x53_inr_Foreach_sm ( // @[sm_x53_inr_Foreach.scala 32:18:@1849.4]
    .clock(x53_inr_Foreach_sm_clock),
    .reset(x53_inr_Foreach_sm_reset),
    .io_enable(x53_inr_Foreach_sm_io_enable),
    .io_done(x53_inr_Foreach_sm_io_done),
    .io_ctrDone(x53_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x53_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x53_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x53_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x53_inr_Foreach_sm_io_parentAck),
    .io_break(x53_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@1877.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@1917.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@1925.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x53_inr_Foreach_kernelx53_inr_Foreach_concrete1 x53_inr_Foreach_kernelx53_inr_Foreach_concrete1 ( // @[sm_x53_inr_Foreach.scala 72:24:@1956.4]
    .io_in_x38_x(x53_inr_Foreach_kernelx53_inr_Foreach_concrete1_io_in_x38_x),
    .io_in_x43_mem_0_wPort_0_ofs_0(x53_inr_Foreach_kernelx53_inr_Foreach_concrete1_io_in_x43_mem_0_wPort_0_ofs_0),
    .io_in_x43_mem_0_wPort_0_data_0(x53_inr_Foreach_kernelx53_inr_Foreach_concrete1_io_in_x43_mem_0_wPort_0_data_0),
    .io_in_x43_mem_0_wPort_0_en_0(x53_inr_Foreach_kernelx53_inr_Foreach_concrete1_io_in_x43_mem_0_wPort_0_en_0),
    .io_sigsIn_datapathEn(x53_inr_Foreach_kernelx53_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x53_inr_Foreach_kernelx53_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_0(x53_inr_Foreach_kernelx53_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x53_inr_Foreach_kernelx53_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_rr(x53_inr_Foreach_kernelx53_inr_Foreach_concrete1_io_rr)
  );
  x53_inr_Foreach_sm x57_inr_UnitPipe_sm ( // @[sm_x57_inr_UnitPipe.scala 32:18:@2069.4]
    .clock(x57_inr_UnitPipe_sm_clock),
    .reset(x57_inr_UnitPipe_sm_reset),
    .io_enable(x57_inr_UnitPipe_sm_io_enable),
    .io_done(x57_inr_UnitPipe_sm_io_done),
    .io_ctrDone(x57_inr_UnitPipe_sm_io_ctrDone),
    .io_datapathEn(x57_inr_UnitPipe_sm_io_datapathEn),
    .io_ctrInc(x57_inr_UnitPipe_sm_io_ctrInc),
    .io_ctrRst(x57_inr_UnitPipe_sm_io_ctrRst),
    .io_parentAck(x57_inr_UnitPipe_sm_io_parentAck),
    .io_break(x57_inr_UnitPipe_sm_io_break)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@2126.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@2134.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  x57_inr_UnitPipe_kernelx57_inr_UnitPipe_concrete1 x57_inr_UnitPipe_kernelx57_inr_UnitPipe_concrete1 ( // @[sm_x57_inr_UnitPipe.scala 70:24:@2160.4]
    .io_in_x43_mem_0_rPort_0_en_0(x57_inr_UnitPipe_kernelx57_inr_UnitPipe_concrete1_io_in_x43_mem_0_rPort_0_en_0),
    .io_in_x43_mem_0_rPort_0_output_0(x57_inr_UnitPipe_kernelx57_inr_UnitPipe_concrete1_io_in_x43_mem_0_rPort_0_output_0),
    .io_in_x39_y_port_0_valid(x57_inr_UnitPipe_kernelx57_inr_UnitPipe_concrete1_io_in_x39_y_port_0_valid),
    .io_in_x39_y_port_0_bits(x57_inr_UnitPipe_kernelx57_inr_UnitPipe_concrete1_io_in_x39_y_port_0_bits),
    .io_sigsIn_datapathEn(x57_inr_UnitPipe_kernelx57_inr_UnitPipe_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x57_inr_UnitPipe_kernelx57_inr_UnitPipe_concrete1_io_sigsIn_break),
    .io_rr(x57_inr_UnitPipe_kernelx57_inr_UnitPipe_concrete1_io_rr)
  );
  assign _T_200 = RetimeWrapper_io_out; // @[package.scala 96:25:@1882.4 package.scala 96:25:@1883.4]
  assign _T_215 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@1922.4 package.scala 96:25:@1923.4]
  assign _T_221 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@1930.4 package.scala 96:25:@1931.4]
  assign _T_224 = ~ _T_221; // @[SpatialBlocks.scala 110:93:@1933.4]
  assign _T_226 = x53_inr_Foreach_sm_io_datapathEn; // @[SpatialBlocks.scala 128:36:@1942.4]
  assign _T_227 = ~ x53_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 128:78:@1943.4]
  assign _T_292 = x57_inr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@2097.4]
  assign _T_309 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@2131.4 package.scala 96:25:@2132.4]
  assign _T_315 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@2139.4 package.scala 96:25:@2140.4]
  assign _T_318 = ~ _T_315; // @[SpatialBlocks.scala 110:93:@2142.4]
  assign io_in_x39_y_port_0_valid = x57_inr_UnitPipe_kernelx57_inr_UnitPipe_concrete1_io_in_x39_y_port_0_valid; // @[MemInterfaceType.scala 317:38:@2213.4]
  assign io_in_x39_y_port_0_bits = x57_inr_UnitPipe_kernelx57_inr_UnitPipe_concrete1_io_in_x39_y_port_0_bits; // @[MemInterfaceType.scala 317:38:@2212.4]
  assign io_sigsOut_smDoneIn_0 = x53_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 127:53:@1940.4]
  assign io_sigsOut_smDoneIn_1 = x57_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 127:53:@2149.4]
  assign x43_mem_0_clock = clock; // @[:@1781.4]
  assign x43_mem_0_reset = reset; // @[:@1782.4]
  assign x43_mem_0_io_rPort_0_en_0 = x57_inr_UnitPipe_kernelx57_inr_UnitPipe_concrete1_io_in_x43_mem_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@2209.4]
  assign x43_mem_0_io_wPort_0_ofs_0 = x53_inr_Foreach_kernelx53_inr_Foreach_concrete1_io_in_x43_mem_0_wPort_0_ofs_0; // @[MemInterfaceType.scala 67:44:@2006.4]
  assign x43_mem_0_io_wPort_0_data_0 = x53_inr_Foreach_kernelx53_inr_Foreach_concrete1_io_in_x43_mem_0_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@2005.4]
  assign x43_mem_0_io_wPort_0_en_0 = x53_inr_Foreach_kernelx53_inr_Foreach_concrete1_io_in_x43_mem_0_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@2001.4]
  assign x45_ctrchain_clock = clock; // @[:@1798.4]
  assign x45_ctrchain_reset = reset; // @[:@1799.4]
  assign x45_ctrchain_io_input_reset = x53_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 130:103:@1955.4]
  assign x45_ctrchain_io_input_enable = x53_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 104:75:@1910.4 SpatialBlocks.scala 130:45:@1954.4]
  assign x53_inr_Foreach_sm_clock = clock; // @[:@1850.4]
  assign x53_inr_Foreach_sm_reset = reset; // @[:@1851.4]
  assign x53_inr_Foreach_sm_io_enable = _T_215 & _T_224; // @[SpatialBlocks.scala 112:18:@1937.4]
  assign x53_inr_Foreach_sm_io_ctrDone = io_rr ? _T_200 : 1'h0; // @[sm_RootController.scala 67:37:@1885.4]
  assign x53_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 114:21:@1939.4]
  assign x53_inr_Foreach_sm_io_break = 1'h0; // @[sm_RootController.scala 71:35:@1891.4]
  assign RetimeWrapper_clock = clock; // @[:@1878.4]
  assign RetimeWrapper_reset = reset; // @[:@1879.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@1881.4]
  assign RetimeWrapper_io_in = x45_ctrchain_io_output_done; // @[package.scala 94:16:@1880.4]
  assign RetimeWrapper_1_clock = clock; // @[:@1918.4]
  assign RetimeWrapper_1_reset = reset; // @[:@1919.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@1921.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@1920.4]
  assign RetimeWrapper_2_clock = clock; // @[:@1926.4]
  assign RetimeWrapper_2_reset = reset; // @[:@1927.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@1929.4]
  assign RetimeWrapper_2_io_in = x53_inr_Foreach_sm_io_done; // @[package.scala 94:16:@1928.4]
  assign x53_inr_Foreach_kernelx53_inr_Foreach_concrete1_io_in_x38_x = io_in_x38_x; // @[sm_x53_inr_Foreach.scala 48:24:@2000.4]
  assign x53_inr_Foreach_kernelx53_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_226 & _T_227; // @[sm_x53_inr_Foreach.scala 76:22:@2020.4]
  assign x53_inr_Foreach_kernelx53_inr_Foreach_concrete1_io_sigsIn_break = x53_inr_Foreach_sm_io_break; // @[sm_x53_inr_Foreach.scala 76:22:@2018.4]
  assign x53_inr_Foreach_kernelx53_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = x45_ctrchain_io_output_counts_0; // @[sm_x53_inr_Foreach.scala 76:22:@2013.4]
  assign x53_inr_Foreach_kernelx53_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x45_ctrchain_io_output_oobs_0; // @[sm_x53_inr_Foreach.scala 76:22:@2012.4]
  assign x53_inr_Foreach_kernelx53_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x53_inr_Foreach.scala 75:18:@2008.4]
  assign x57_inr_UnitPipe_sm_clock = clock; // @[:@2070.4]
  assign x57_inr_UnitPipe_sm_reset = reset; // @[:@2071.4]
  assign x57_inr_UnitPipe_sm_io_enable = _T_309 & _T_318; // @[SpatialBlocks.scala 112:18:@2146.4]
  assign x57_inr_UnitPipe_sm_io_ctrDone = x57_inr_UnitPipe_sm_io_ctrInc & _T_295; // @[sm_RootController.scala 76:38:@2101.4]
  assign x57_inr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 114:21:@2148.4]
  assign x57_inr_UnitPipe_sm_io_break = 1'h0; // @[sm_RootController.scala 80:36:@2107.4]
  assign RetimeWrapper_3_clock = clock; // @[:@2127.4]
  assign RetimeWrapper_3_reset = reset; // @[:@2128.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@2130.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@2129.4]
  assign RetimeWrapper_4_clock = clock; // @[:@2135.4]
  assign RetimeWrapper_4_reset = reset; // @[:@2136.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@2138.4]
  assign RetimeWrapper_4_io_in = x57_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@2137.4]
  assign x57_inr_UnitPipe_kernelx57_inr_UnitPipe_concrete1_io_in_x43_mem_0_rPort_0_output_0 = x43_mem_0_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@2207.4]
  assign x57_inr_UnitPipe_kernelx57_inr_UnitPipe_concrete1_io_sigsIn_datapathEn = x57_inr_UnitPipe_sm_io_datapathEn; // @[sm_x57_inr_UnitPipe.scala 74:22:@2229.4]
  assign x57_inr_UnitPipe_kernelx57_inr_UnitPipe_concrete1_io_sigsIn_break = x57_inr_UnitPipe_sm_io_break; // @[sm_x57_inr_UnitPipe.scala 74:22:@2227.4]
  assign x57_inr_UnitPipe_kernelx57_inr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x57_inr_UnitPipe.scala 73:18:@2217.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_295 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_295 <= 1'h0;
    end else begin
      _T_295 <= _T_292;
    end
  end
endmodule
module AccelTop( // @[:@2244.2]
  input         clock, // @[:@2245.4]
  input         reset, // @[:@2246.4]
  input         io_enable, // @[:@2247.4]
  output        io_done, // @[:@2247.4]
  input         io_reset, // @[:@2247.4]
  input         io_memStreams_loads_0_cmd_ready, // @[:@2247.4]
  output        io_memStreams_loads_0_cmd_valid, // @[:@2247.4]
  output [63:0] io_memStreams_loads_0_cmd_bits_addr, // @[:@2247.4]
  output [31:0] io_memStreams_loads_0_cmd_bits_size, // @[:@2247.4]
  output        io_memStreams_loads_0_data_ready, // @[:@2247.4]
  input         io_memStreams_loads_0_data_valid, // @[:@2247.4]
  input  [31:0] io_memStreams_loads_0_data_bits_rdata_0, // @[:@2247.4]
  input  [31:0] io_memStreams_loads_0_data_bits_rdata_1, // @[:@2247.4]
  input  [31:0] io_memStreams_loads_0_data_bits_rdata_2, // @[:@2247.4]
  input  [31:0] io_memStreams_loads_0_data_bits_rdata_3, // @[:@2247.4]
  input  [31:0] io_memStreams_loads_0_data_bits_rdata_4, // @[:@2247.4]
  input  [31:0] io_memStreams_loads_0_data_bits_rdata_5, // @[:@2247.4]
  input  [31:0] io_memStreams_loads_0_data_bits_rdata_6, // @[:@2247.4]
  input  [31:0] io_memStreams_loads_0_data_bits_rdata_7, // @[:@2247.4]
  input  [31:0] io_memStreams_loads_0_data_bits_rdata_8, // @[:@2247.4]
  input  [31:0] io_memStreams_loads_0_data_bits_rdata_9, // @[:@2247.4]
  input  [31:0] io_memStreams_loads_0_data_bits_rdata_10, // @[:@2247.4]
  input  [31:0] io_memStreams_loads_0_data_bits_rdata_11, // @[:@2247.4]
  input  [31:0] io_memStreams_loads_0_data_bits_rdata_12, // @[:@2247.4]
  input  [31:0] io_memStreams_loads_0_data_bits_rdata_13, // @[:@2247.4]
  input  [31:0] io_memStreams_loads_0_data_bits_rdata_14, // @[:@2247.4]
  input  [31:0] io_memStreams_loads_0_data_bits_rdata_15, // @[:@2247.4]
  input         io_memStreams_stores_0_cmd_ready, // @[:@2247.4]
  output        io_memStreams_stores_0_cmd_valid, // @[:@2247.4]
  output [63:0] io_memStreams_stores_0_cmd_bits_addr, // @[:@2247.4]
  output [31:0] io_memStreams_stores_0_cmd_bits_size, // @[:@2247.4]
  input         io_memStreams_stores_0_data_ready, // @[:@2247.4]
  output        io_memStreams_stores_0_data_valid, // @[:@2247.4]
  output [31:0] io_memStreams_stores_0_data_bits_wdata_0, // @[:@2247.4]
  output [31:0] io_memStreams_stores_0_data_bits_wdata_1, // @[:@2247.4]
  output [31:0] io_memStreams_stores_0_data_bits_wdata_2, // @[:@2247.4]
  output [31:0] io_memStreams_stores_0_data_bits_wdata_3, // @[:@2247.4]
  output [31:0] io_memStreams_stores_0_data_bits_wdata_4, // @[:@2247.4]
  output [31:0] io_memStreams_stores_0_data_bits_wdata_5, // @[:@2247.4]
  output [31:0] io_memStreams_stores_0_data_bits_wdata_6, // @[:@2247.4]
  output [31:0] io_memStreams_stores_0_data_bits_wdata_7, // @[:@2247.4]
  output [31:0] io_memStreams_stores_0_data_bits_wdata_8, // @[:@2247.4]
  output [31:0] io_memStreams_stores_0_data_bits_wdata_9, // @[:@2247.4]
  output [31:0] io_memStreams_stores_0_data_bits_wdata_10, // @[:@2247.4]
  output [31:0] io_memStreams_stores_0_data_bits_wdata_11, // @[:@2247.4]
  output [31:0] io_memStreams_stores_0_data_bits_wdata_12, // @[:@2247.4]
  output [31:0] io_memStreams_stores_0_data_bits_wdata_13, // @[:@2247.4]
  output [31:0] io_memStreams_stores_0_data_bits_wdata_14, // @[:@2247.4]
  output [31:0] io_memStreams_stores_0_data_bits_wdata_15, // @[:@2247.4]
  output [15:0] io_memStreams_stores_0_data_bits_wstrb, // @[:@2247.4]
  output        io_memStreams_stores_0_wresp_ready, // @[:@2247.4]
  input         io_memStreams_stores_0_wresp_valid, // @[:@2247.4]
  input         io_memStreams_stores_0_wresp_bits, // @[:@2247.4]
  input         io_memStreams_gathers_0_cmd_ready, // @[:@2247.4]
  output        io_memStreams_gathers_0_cmd_valid, // @[:@2247.4]
  output [63:0] io_memStreams_gathers_0_cmd_bits_addr_0, // @[:@2247.4]
  output [63:0] io_memStreams_gathers_0_cmd_bits_addr_1, // @[:@2247.4]
  output [63:0] io_memStreams_gathers_0_cmd_bits_addr_2, // @[:@2247.4]
  output [63:0] io_memStreams_gathers_0_cmd_bits_addr_3, // @[:@2247.4]
  output [63:0] io_memStreams_gathers_0_cmd_bits_addr_4, // @[:@2247.4]
  output [63:0] io_memStreams_gathers_0_cmd_bits_addr_5, // @[:@2247.4]
  output [63:0] io_memStreams_gathers_0_cmd_bits_addr_6, // @[:@2247.4]
  output [63:0] io_memStreams_gathers_0_cmd_bits_addr_7, // @[:@2247.4]
  output [63:0] io_memStreams_gathers_0_cmd_bits_addr_8, // @[:@2247.4]
  output [63:0] io_memStreams_gathers_0_cmd_bits_addr_9, // @[:@2247.4]
  output [63:0] io_memStreams_gathers_0_cmd_bits_addr_10, // @[:@2247.4]
  output [63:0] io_memStreams_gathers_0_cmd_bits_addr_11, // @[:@2247.4]
  output [63:0] io_memStreams_gathers_0_cmd_bits_addr_12, // @[:@2247.4]
  output [63:0] io_memStreams_gathers_0_cmd_bits_addr_13, // @[:@2247.4]
  output [63:0] io_memStreams_gathers_0_cmd_bits_addr_14, // @[:@2247.4]
  output [63:0] io_memStreams_gathers_0_cmd_bits_addr_15, // @[:@2247.4]
  output        io_memStreams_gathers_0_data_ready, // @[:@2247.4]
  input         io_memStreams_gathers_0_data_valid, // @[:@2247.4]
  input  [31:0] io_memStreams_gathers_0_data_bits_0, // @[:@2247.4]
  input  [31:0] io_memStreams_gathers_0_data_bits_1, // @[:@2247.4]
  input  [31:0] io_memStreams_gathers_0_data_bits_2, // @[:@2247.4]
  input  [31:0] io_memStreams_gathers_0_data_bits_3, // @[:@2247.4]
  input  [31:0] io_memStreams_gathers_0_data_bits_4, // @[:@2247.4]
  input  [31:0] io_memStreams_gathers_0_data_bits_5, // @[:@2247.4]
  input  [31:0] io_memStreams_gathers_0_data_bits_6, // @[:@2247.4]
  input  [31:0] io_memStreams_gathers_0_data_bits_7, // @[:@2247.4]
  input  [31:0] io_memStreams_gathers_0_data_bits_8, // @[:@2247.4]
  input  [31:0] io_memStreams_gathers_0_data_bits_9, // @[:@2247.4]
  input  [31:0] io_memStreams_gathers_0_data_bits_10, // @[:@2247.4]
  input  [31:0] io_memStreams_gathers_0_data_bits_11, // @[:@2247.4]
  input  [31:0] io_memStreams_gathers_0_data_bits_12, // @[:@2247.4]
  input  [31:0] io_memStreams_gathers_0_data_bits_13, // @[:@2247.4]
  input  [31:0] io_memStreams_gathers_0_data_bits_14, // @[:@2247.4]
  input  [31:0] io_memStreams_gathers_0_data_bits_15, // @[:@2247.4]
  input         io_memStreams_scatters_0_cmd_ready, // @[:@2247.4]
  output        io_memStreams_scatters_0_cmd_valid, // @[:@2247.4]
  output [63:0] io_memStreams_scatters_0_cmd_bits_addr_addr_0, // @[:@2247.4]
  output [63:0] io_memStreams_scatters_0_cmd_bits_addr_addr_1, // @[:@2247.4]
  output [63:0] io_memStreams_scatters_0_cmd_bits_addr_addr_2, // @[:@2247.4]
  output [63:0] io_memStreams_scatters_0_cmd_bits_addr_addr_3, // @[:@2247.4]
  output [63:0] io_memStreams_scatters_0_cmd_bits_addr_addr_4, // @[:@2247.4]
  output [63:0] io_memStreams_scatters_0_cmd_bits_addr_addr_5, // @[:@2247.4]
  output [63:0] io_memStreams_scatters_0_cmd_bits_addr_addr_6, // @[:@2247.4]
  output [63:0] io_memStreams_scatters_0_cmd_bits_addr_addr_7, // @[:@2247.4]
  output [63:0] io_memStreams_scatters_0_cmd_bits_addr_addr_8, // @[:@2247.4]
  output [63:0] io_memStreams_scatters_0_cmd_bits_addr_addr_9, // @[:@2247.4]
  output [63:0] io_memStreams_scatters_0_cmd_bits_addr_addr_10, // @[:@2247.4]
  output [63:0] io_memStreams_scatters_0_cmd_bits_addr_addr_11, // @[:@2247.4]
  output [63:0] io_memStreams_scatters_0_cmd_bits_addr_addr_12, // @[:@2247.4]
  output [63:0] io_memStreams_scatters_0_cmd_bits_addr_addr_13, // @[:@2247.4]
  output [63:0] io_memStreams_scatters_0_cmd_bits_addr_addr_14, // @[:@2247.4]
  output [63:0] io_memStreams_scatters_0_cmd_bits_addr_addr_15, // @[:@2247.4]
  output [31:0] io_memStreams_scatters_0_cmd_bits_wdata_0, // @[:@2247.4]
  output [31:0] io_memStreams_scatters_0_cmd_bits_wdata_1, // @[:@2247.4]
  output [31:0] io_memStreams_scatters_0_cmd_bits_wdata_2, // @[:@2247.4]
  output [31:0] io_memStreams_scatters_0_cmd_bits_wdata_3, // @[:@2247.4]
  output [31:0] io_memStreams_scatters_0_cmd_bits_wdata_4, // @[:@2247.4]
  output [31:0] io_memStreams_scatters_0_cmd_bits_wdata_5, // @[:@2247.4]
  output [31:0] io_memStreams_scatters_0_cmd_bits_wdata_6, // @[:@2247.4]
  output [31:0] io_memStreams_scatters_0_cmd_bits_wdata_7, // @[:@2247.4]
  output [31:0] io_memStreams_scatters_0_cmd_bits_wdata_8, // @[:@2247.4]
  output [31:0] io_memStreams_scatters_0_cmd_bits_wdata_9, // @[:@2247.4]
  output [31:0] io_memStreams_scatters_0_cmd_bits_wdata_10, // @[:@2247.4]
  output [31:0] io_memStreams_scatters_0_cmd_bits_wdata_11, // @[:@2247.4]
  output [31:0] io_memStreams_scatters_0_cmd_bits_wdata_12, // @[:@2247.4]
  output [31:0] io_memStreams_scatters_0_cmd_bits_wdata_13, // @[:@2247.4]
  output [31:0] io_memStreams_scatters_0_cmd_bits_wdata_14, // @[:@2247.4]
  output [31:0] io_memStreams_scatters_0_cmd_bits_wdata_15, // @[:@2247.4]
  output        io_memStreams_scatters_0_wresp_ready, // @[:@2247.4]
  input         io_memStreams_scatters_0_wresp_valid, // @[:@2247.4]
  input         io_memStreams_scatters_0_wresp_bits, // @[:@2247.4]
  output        io_heap_0_req_valid, // @[:@2247.4]
  output        io_heap_0_req_bits_allocDealloc, // @[:@2247.4]
  output [63:0] io_heap_0_req_bits_sizeAddr, // @[:@2247.4]
  input         io_heap_0_resp_valid, // @[:@2247.4]
  input         io_heap_0_resp_bits_allocDealloc, // @[:@2247.4]
  input  [63:0] io_heap_0_resp_bits_sizeAddr, // @[:@2247.4]
  input  [63:0] io_argIns_0, // @[:@2247.4]
  input         io_argOuts_0_port_ready, // @[:@2247.4]
  output        io_argOuts_0_port_valid, // @[:@2247.4]
  output [63:0] io_argOuts_0_port_bits, // @[:@2247.4]
  input  [63:0] io_argOuts_0_echo // @[:@2247.4]
);
  wire  SingleCounter_clock; // @[Main.scala 32:32:@2395.4]
  wire  SingleCounter_reset; // @[Main.scala 32:32:@2395.4]
  wire  SingleCounter_io_input_reset; // @[Main.scala 32:32:@2395.4]
  wire  SingleCounter_io_output_done; // @[Main.scala 32:32:@2395.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@2413.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@2413.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@2413.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@2413.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@2413.4]
  wire  SRFF_clock; // @[Main.scala 36:28:@2422.4]
  wire  SRFF_reset; // @[Main.scala 36:28:@2422.4]
  wire  SRFF_io_input_set; // @[Main.scala 36:28:@2422.4]
  wire  SRFF_io_input_reset; // @[Main.scala 36:28:@2422.4]
  wire  SRFF_io_input_asyn_reset; // @[Main.scala 36:28:@2422.4]
  wire  SRFF_io_output; // @[Main.scala 36:28:@2422.4]
  wire  RootController_sm_clock; // @[sm_RootController.scala 32:18:@2465.4]
  wire  RootController_sm_reset; // @[sm_RootController.scala 32:18:@2465.4]
  wire  RootController_sm_io_enable; // @[sm_RootController.scala 32:18:@2465.4]
  wire  RootController_sm_io_done; // @[sm_RootController.scala 32:18:@2465.4]
  wire  RootController_sm_io_rst; // @[sm_RootController.scala 32:18:@2465.4]
  wire  RootController_sm_io_ctrDone; // @[sm_RootController.scala 32:18:@2465.4]
  wire  RootController_sm_io_ctrInc; // @[sm_RootController.scala 32:18:@2465.4]
  wire  RootController_sm_io_doneIn_0; // @[sm_RootController.scala 32:18:@2465.4]
  wire  RootController_sm_io_doneIn_1; // @[sm_RootController.scala 32:18:@2465.4]
  wire  RootController_sm_io_enableOut_0; // @[sm_RootController.scala 32:18:@2465.4]
  wire  RootController_sm_io_enableOut_1; // @[sm_RootController.scala 32:18:@2465.4]
  wire  RootController_sm_io_childAck_0; // @[sm_RootController.scala 32:18:@2465.4]
  wire  RootController_sm_io_childAck_1; // @[sm_RootController.scala 32:18:@2465.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@2502.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@2502.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@2502.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@2502.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@2502.4]
  wire  RootController_kernelRootController_concrete1_clock; // @[sm_RootController.scala 85:24:@2566.4]
  wire  RootController_kernelRootController_concrete1_reset; // @[sm_RootController.scala 85:24:@2566.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x38_x; // @[sm_RootController.scala 85:24:@2566.4]
  wire  RootController_kernelRootController_concrete1_io_in_x39_y_port_0_valid; // @[sm_RootController.scala 85:24:@2566.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x39_y_port_0_bits; // @[sm_RootController.scala 85:24:@2566.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_RootController.scala 85:24:@2566.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_RootController.scala 85:24:@2566.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0; // @[sm_RootController.scala 85:24:@2566.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_1; // @[sm_RootController.scala 85:24:@2566.4]
  wire  RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[sm_RootController.scala 85:24:@2566.4]
  wire  RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_1; // @[sm_RootController.scala 85:24:@2566.4]
  wire  RootController_kernelRootController_concrete1_io_rr; // @[sm_RootController.scala 85:24:@2566.4]
  wire  _T_555; // @[package.scala 96:25:@2418.4 package.scala 96:25:@2419.4]
  wire  _T_620; // @[Main.scala 38:44:@2498.4]
  wire  _T_621; // @[Main.scala 38:53:@2499.4]
  wire  _T_633; // @[package.scala 100:49:@2519.4]
  reg  _T_636; // @[package.scala 48:56:@2520.4]
  reg [31:0] _RAND_0;
  SingleCounter SingleCounter ( // @[Main.scala 32:32:@2395.4]
    .clock(SingleCounter_clock),
    .reset(SingleCounter_reset),
    .io_input_reset(SingleCounter_io_input_reset),
    .io_output_done(SingleCounter_io_output_done)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@2413.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  SRFF SRFF ( // @[Main.scala 36:28:@2422.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  RootController_sm RootController_sm ( // @[sm_RootController.scala 32:18:@2465.4]
    .clock(RootController_sm_clock),
    .reset(RootController_sm_reset),
    .io_enable(RootController_sm_io_enable),
    .io_done(RootController_sm_io_done),
    .io_rst(RootController_sm_io_rst),
    .io_ctrDone(RootController_sm_io_ctrDone),
    .io_ctrInc(RootController_sm_io_ctrInc),
    .io_doneIn_0(RootController_sm_io_doneIn_0),
    .io_doneIn_1(RootController_sm_io_doneIn_1),
    .io_enableOut_0(RootController_sm_io_enableOut_0),
    .io_enableOut_1(RootController_sm_io_enableOut_1),
    .io_childAck_0(RootController_sm_io_childAck_0),
    .io_childAck_1(RootController_sm_io_childAck_1)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@2502.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RootController_kernelRootController_concrete1 RootController_kernelRootController_concrete1 ( // @[sm_RootController.scala 85:24:@2566.4]
    .clock(RootController_kernelRootController_concrete1_clock),
    .reset(RootController_kernelRootController_concrete1_reset),
    .io_in_x38_x(RootController_kernelRootController_concrete1_io_in_x38_x),
    .io_in_x39_y_port_0_valid(RootController_kernelRootController_concrete1_io_in_x39_y_port_0_valid),
    .io_in_x39_y_port_0_bits(RootController_kernelRootController_concrete1_io_in_x39_y_port_0_bits),
    .io_sigsIn_smEnableOuts_0(RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smChildAcks_0(RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsOut_smDoneIn_0(RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_1),
    .io_rr(RootController_kernelRootController_concrete1_io_rr)
  );
  assign _T_555 = RetimeWrapper_io_out; // @[package.scala 96:25:@2418.4 package.scala 96:25:@2419.4]
  assign _T_620 = io_enable & _T_555; // @[Main.scala 38:44:@2498.4]
  assign _T_621 = ~ SRFF_io_output; // @[Main.scala 38:53:@2499.4]
  assign _T_633 = RootController_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@2519.4]
  assign io_done = SRFF_io_output; // @[Main.scala 45:17:@2518.4]
  assign io_memStreams_loads_0_cmd_valid = 1'h0;
  assign io_memStreams_loads_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_loads_0_cmd_bits_size = 32'h0;
  assign io_memStreams_loads_0_data_ready = 1'h0;
  assign io_memStreams_stores_0_cmd_valid = 1'h0;
  assign io_memStreams_stores_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_stores_0_cmd_bits_size = 32'h0;
  assign io_memStreams_stores_0_data_valid = 1'h0;
  assign io_memStreams_stores_0_data_bits_wdata_0 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_1 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_2 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_3 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_4 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_5 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_6 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_7 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_8 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_9 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_10 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_11 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_12 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_13 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_14 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_15 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wstrb = 16'h0;
  assign io_memStreams_stores_0_wresp_ready = 1'h0;
  assign io_memStreams_gathers_0_cmd_valid = 1'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_0 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_1 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_2 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_3 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_4 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_5 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_6 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_7 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_8 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_9 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_10 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_11 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_12 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_13 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_14 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_15 = 64'h0;
  assign io_memStreams_gathers_0_data_ready = 1'h0;
  assign io_memStreams_scatters_0_cmd_valid = 1'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_0 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_1 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_2 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_3 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_4 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_5 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_6 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_7 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_8 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_9 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_10 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_11 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_12 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_13 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_14 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_15 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_0 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_1 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_2 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_3 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_4 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_5 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_6 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_7 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_8 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_9 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_10 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_11 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_12 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_13 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_14 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_15 = 32'h0;
  assign io_memStreams_scatters_0_wresp_ready = 1'h0;
  assign io_heap_0_req_valid = 1'h0;
  assign io_heap_0_req_bits_allocDealloc = 1'h0;
  assign io_heap_0_req_bits_sizeAddr = 64'h0;
  assign io_argOuts_0_port_valid = RootController_kernelRootController_concrete1_io_in_x39_y_port_0_valid; // @[Main.scala 28:57:@2391.4]
  assign io_argOuts_0_port_bits = RootController_kernelRootController_concrete1_io_in_x39_y_port_0_bits; // @[Main.scala 29:56:@2392.4]
  assign SingleCounter_clock = clock; // @[:@2396.4]
  assign SingleCounter_reset = reset; // @[:@2397.4]
  assign SingleCounter_io_input_reset = reset; // @[Main.scala 33:79:@2411.4]
  assign RetimeWrapper_clock = clock; // @[:@2414.4]
  assign RetimeWrapper_reset = reset; // @[:@2415.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@2417.4]
  assign RetimeWrapper_io_in = SingleCounter_io_output_done; // @[package.scala 94:16:@2416.4]
  assign SRFF_clock = clock; // @[:@2423.4]
  assign SRFF_reset = reset; // @[:@2424.4]
  assign SRFF_io_input_set = RootController_sm_io_done; // @[Main.scala 54:29:@2643.4]
  assign SRFF_io_input_reset = RetimeWrapper_1_io_out; // @[Main.scala 43:31:@2516.4]
  assign SRFF_io_input_asyn_reset = RetimeWrapper_1_io_out; // @[Main.scala 44:36:@2517.4]
  assign RootController_sm_clock = clock; // @[:@2466.4]
  assign RootController_sm_reset = reset; // @[:@2467.4]
  assign RootController_sm_io_enable = _T_620 & _T_621; // @[Main.scala 42:33:@2515.4 SpatialBlocks.scala 112:18:@2554.4]
  assign RootController_sm_io_rst = RetimeWrapper_1_io_out; // @[SpatialBlocks.scala 106:15:@2548.4]
  assign RootController_sm_io_ctrDone = RootController_sm_io_ctrInc & _T_636; // @[Main.scala 46:34:@2523.4]
  assign RootController_sm_io_doneIn_0 = RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 102:67:@2543.4]
  assign RootController_sm_io_doneIn_1 = RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 102:67:@2544.4]
  assign RetimeWrapper_1_clock = clock; // @[:@2503.4]
  assign RetimeWrapper_1_reset = reset; // @[:@2504.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@2506.4]
  assign RetimeWrapper_1_io_in = reset | io_reset; // @[package.scala 94:16:@2505.4]
  assign RootController_kernelRootController_concrete1_clock = clock; // @[:@2567.4]
  assign RootController_kernelRootController_concrete1_reset = reset; // @[:@2568.4]
  assign RootController_kernelRootController_concrete1_io_in_x38_x = io_argIns_0; // @[sm_RootController.scala 48:24:@2606.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0 = RootController_sm_io_enableOut_0; // @[sm_RootController.scala 89:22:@2622.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_1 = RootController_sm_io_enableOut_1; // @[sm_RootController.scala 89:22:@2623.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0 = RootController_sm_io_childAck_0; // @[sm_RootController.scala 89:22:@2618.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_1 = RootController_sm_io_childAck_1; // @[sm_RootController.scala 89:22:@2619.4]
  assign RootController_kernelRootController_concrete1_io_rr = RetimeWrapper_io_out; // @[sm_RootController.scala 88:18:@2612.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_636 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_636 <= 1'h0;
    end else begin
      _T_636 <= _T_633;
    end
  end
endmodule
module DRAMHeap( // @[:@3550.2]
  input         io_accel_0_req_valid, // @[:@3553.4]
  input         io_accel_0_req_bits_allocDealloc, // @[:@3553.4]
  input  [63:0] io_accel_0_req_bits_sizeAddr, // @[:@3553.4]
  output        io_accel_0_resp_valid, // @[:@3553.4]
  output        io_accel_0_resp_bits_allocDealloc, // @[:@3553.4]
  output [63:0] io_accel_0_resp_bits_sizeAddr, // @[:@3553.4]
  output        io_host_0_req_valid, // @[:@3553.4]
  output        io_host_0_req_bits_allocDealloc, // @[:@3553.4]
  output [63:0] io_host_0_req_bits_sizeAddr, // @[:@3553.4]
  input         io_host_0_resp_valid, // @[:@3553.4]
  input         io_host_0_resp_bits_allocDealloc, // @[:@3553.4]
  input  [63:0] io_host_0_resp_bits_sizeAddr // @[:@3553.4]
);
  assign io_accel_0_resp_valid = io_host_0_resp_valid; // @[DRAMHeap.scala 24:18:@3560.4]
  assign io_accel_0_resp_bits_allocDealloc = io_host_0_resp_bits_allocDealloc; // @[DRAMHeap.scala 25:17:@3562.4]
  assign io_accel_0_resp_bits_sizeAddr = io_host_0_resp_bits_sizeAddr; // @[DRAMHeap.scala 25:17:@3561.4]
  assign io_host_0_req_valid = io_accel_0_req_valid; // @[DRAMHeap.scala 21:18:@3557.4]
  assign io_host_0_req_bits_allocDealloc = io_accel_0_req_bits_allocDealloc; // @[DRAMHeap.scala 21:18:@3556.4]
  assign io_host_0_req_bits_sizeAddr = io_accel_0_req_bits_sizeAddr; // @[DRAMHeap.scala 21:18:@3555.4]
endmodule
module RetimeWrapper_15( // @[:@3576.2]
  input         clock, // @[:@3577.4]
  input         reset, // @[:@3578.4]
  input         io_flow, // @[:@3579.4]
  input  [63:0] io_in, // @[:@3579.4]
  output [63:0] io_out // @[:@3579.4]
);
  wire [63:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@3581.4]
  wire [63:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@3581.4]
  wire [63:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@3581.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3581.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3581.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3581.4]
  RetimeShiftRegister #(.WIDTH(64), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@3581.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3594.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3593.4]
  assign sr_init = 64'h0; // @[RetimeShiftRegister.scala 19:16:@3592.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3591.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3590.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3588.4]
endmodule
module FringeFF( // @[:@3596.2]
  input         clock, // @[:@3597.4]
  input         reset, // @[:@3598.4]
  input  [63:0] io_in, // @[:@3599.4]
  input         io_reset, // @[:@3599.4]
  output [63:0] io_out, // @[:@3599.4]
  input         io_enable // @[:@3599.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3602.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3602.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3602.4]
  wire [63:0] RetimeWrapper_io_in; // @[package.scala 93:22:@3602.4]
  wire [63:0] RetimeWrapper_io_out; // @[package.scala 93:22:@3602.4]
  wire [63:0] _T_18; // @[package.scala 96:25:@3607.4 package.scala 96:25:@3608.4]
  wire [63:0] _GEN_0; // @[FringeFF.scala 21:27:@3613.6]
  RetimeWrapper_15 RetimeWrapper ( // @[package.scala 93:22:@3602.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@3607.4 package.scala 96:25:@3608.4]
  assign _GEN_0 = io_reset ? 64'h0 : _T_18; // @[FringeFF.scala 21:27:@3613.6]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@3619.4]
  assign RetimeWrapper_clock = clock; // @[:@3603.4]
  assign RetimeWrapper_reset = reset; // @[:@3604.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@3606.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _GEN_0; // @[package.scala 94:16:@3605.4]
endmodule
module MuxN( // @[:@32235.2]
  input  [63:0] io_ins_0, // @[:@32238.4]
  input  [63:0] io_ins_1, // @[:@32238.4]
  input  [63:0] io_ins_2, // @[:@32238.4]
  input  [63:0] io_ins_3, // @[:@32238.4]
  input  [63:0] io_ins_4, // @[:@32238.4]
  input  [63:0] io_ins_5, // @[:@32238.4]
  input  [63:0] io_ins_6, // @[:@32238.4]
  input  [63:0] io_ins_7, // @[:@32238.4]
  input  [63:0] io_ins_8, // @[:@32238.4]
  input  [63:0] io_ins_9, // @[:@32238.4]
  input  [63:0] io_ins_10, // @[:@32238.4]
  input  [63:0] io_ins_11, // @[:@32238.4]
  input  [63:0] io_ins_12, // @[:@32238.4]
  input  [63:0] io_ins_13, // @[:@32238.4]
  input  [63:0] io_ins_14, // @[:@32238.4]
  input  [63:0] io_ins_15, // @[:@32238.4]
  input  [63:0] io_ins_16, // @[:@32238.4]
  input  [63:0] io_ins_17, // @[:@32238.4]
  input  [63:0] io_ins_18, // @[:@32238.4]
  input  [63:0] io_ins_19, // @[:@32238.4]
  input  [63:0] io_ins_20, // @[:@32238.4]
  input  [63:0] io_ins_21, // @[:@32238.4]
  input  [63:0] io_ins_22, // @[:@32238.4]
  input  [63:0] io_ins_23, // @[:@32238.4]
  input  [63:0] io_ins_24, // @[:@32238.4]
  input  [63:0] io_ins_25, // @[:@32238.4]
  input  [63:0] io_ins_26, // @[:@32238.4]
  input  [63:0] io_ins_27, // @[:@32238.4]
  input  [63:0] io_ins_28, // @[:@32238.4]
  input  [63:0] io_ins_29, // @[:@32238.4]
  input  [63:0] io_ins_30, // @[:@32238.4]
  input  [63:0] io_ins_31, // @[:@32238.4]
  input  [63:0] io_ins_32, // @[:@32238.4]
  input  [63:0] io_ins_33, // @[:@32238.4]
  input  [63:0] io_ins_34, // @[:@32238.4]
  input  [63:0] io_ins_35, // @[:@32238.4]
  input  [63:0] io_ins_36, // @[:@32238.4]
  input  [63:0] io_ins_37, // @[:@32238.4]
  input  [63:0] io_ins_38, // @[:@32238.4]
  input  [63:0] io_ins_39, // @[:@32238.4]
  input  [63:0] io_ins_40, // @[:@32238.4]
  input  [63:0] io_ins_41, // @[:@32238.4]
  input  [63:0] io_ins_42, // @[:@32238.4]
  input  [63:0] io_ins_43, // @[:@32238.4]
  input  [63:0] io_ins_44, // @[:@32238.4]
  input  [63:0] io_ins_45, // @[:@32238.4]
  input  [63:0] io_ins_46, // @[:@32238.4]
  input  [63:0] io_ins_47, // @[:@32238.4]
  input  [63:0] io_ins_48, // @[:@32238.4]
  input  [63:0] io_ins_49, // @[:@32238.4]
  input  [63:0] io_ins_50, // @[:@32238.4]
  input  [63:0] io_ins_51, // @[:@32238.4]
  input  [63:0] io_ins_52, // @[:@32238.4]
  input  [63:0] io_ins_53, // @[:@32238.4]
  input  [63:0] io_ins_54, // @[:@32238.4]
  input  [63:0] io_ins_55, // @[:@32238.4]
  input  [63:0] io_ins_56, // @[:@32238.4]
  input  [63:0] io_ins_57, // @[:@32238.4]
  input  [63:0] io_ins_58, // @[:@32238.4]
  input  [63:0] io_ins_59, // @[:@32238.4]
  input  [63:0] io_ins_60, // @[:@32238.4]
  input  [63:0] io_ins_61, // @[:@32238.4]
  input  [63:0] io_ins_62, // @[:@32238.4]
  input  [63:0] io_ins_63, // @[:@32238.4]
  input  [63:0] io_ins_64, // @[:@32238.4]
  input  [63:0] io_ins_65, // @[:@32238.4]
  input  [63:0] io_ins_66, // @[:@32238.4]
  input  [63:0] io_ins_67, // @[:@32238.4]
  input  [63:0] io_ins_68, // @[:@32238.4]
  input  [63:0] io_ins_69, // @[:@32238.4]
  input  [63:0] io_ins_70, // @[:@32238.4]
  input  [63:0] io_ins_71, // @[:@32238.4]
  input  [63:0] io_ins_72, // @[:@32238.4]
  input  [63:0] io_ins_73, // @[:@32238.4]
  input  [63:0] io_ins_74, // @[:@32238.4]
  input  [63:0] io_ins_75, // @[:@32238.4]
  input  [63:0] io_ins_76, // @[:@32238.4]
  input  [63:0] io_ins_77, // @[:@32238.4]
  input  [63:0] io_ins_78, // @[:@32238.4]
  input  [63:0] io_ins_79, // @[:@32238.4]
  input  [63:0] io_ins_80, // @[:@32238.4]
  input  [63:0] io_ins_81, // @[:@32238.4]
  input  [63:0] io_ins_82, // @[:@32238.4]
  input  [63:0] io_ins_83, // @[:@32238.4]
  input  [63:0] io_ins_84, // @[:@32238.4]
  input  [63:0] io_ins_85, // @[:@32238.4]
  input  [63:0] io_ins_86, // @[:@32238.4]
  input  [63:0] io_ins_87, // @[:@32238.4]
  input  [63:0] io_ins_88, // @[:@32238.4]
  input  [63:0] io_ins_89, // @[:@32238.4]
  input  [63:0] io_ins_90, // @[:@32238.4]
  input  [63:0] io_ins_91, // @[:@32238.4]
  input  [63:0] io_ins_92, // @[:@32238.4]
  input  [63:0] io_ins_93, // @[:@32238.4]
  input  [63:0] io_ins_94, // @[:@32238.4]
  input  [63:0] io_ins_95, // @[:@32238.4]
  input  [63:0] io_ins_96, // @[:@32238.4]
  input  [63:0] io_ins_97, // @[:@32238.4]
  input  [63:0] io_ins_98, // @[:@32238.4]
  input  [63:0] io_ins_99, // @[:@32238.4]
  input  [63:0] io_ins_100, // @[:@32238.4]
  input  [63:0] io_ins_101, // @[:@32238.4]
  input  [63:0] io_ins_102, // @[:@32238.4]
  input  [63:0] io_ins_103, // @[:@32238.4]
  input  [63:0] io_ins_104, // @[:@32238.4]
  input  [63:0] io_ins_105, // @[:@32238.4]
  input  [63:0] io_ins_106, // @[:@32238.4]
  input  [63:0] io_ins_107, // @[:@32238.4]
  input  [63:0] io_ins_108, // @[:@32238.4]
  input  [63:0] io_ins_109, // @[:@32238.4]
  input  [63:0] io_ins_110, // @[:@32238.4]
  input  [63:0] io_ins_111, // @[:@32238.4]
  input  [63:0] io_ins_112, // @[:@32238.4]
  input  [63:0] io_ins_113, // @[:@32238.4]
  input  [63:0] io_ins_114, // @[:@32238.4]
  input  [63:0] io_ins_115, // @[:@32238.4]
  input  [63:0] io_ins_116, // @[:@32238.4]
  input  [63:0] io_ins_117, // @[:@32238.4]
  input  [63:0] io_ins_118, // @[:@32238.4]
  input  [63:0] io_ins_119, // @[:@32238.4]
  input  [63:0] io_ins_120, // @[:@32238.4]
  input  [63:0] io_ins_121, // @[:@32238.4]
  input  [63:0] io_ins_122, // @[:@32238.4]
  input  [63:0] io_ins_123, // @[:@32238.4]
  input  [63:0] io_ins_124, // @[:@32238.4]
  input  [63:0] io_ins_125, // @[:@32238.4]
  input  [63:0] io_ins_126, // @[:@32238.4]
  input  [63:0] io_ins_127, // @[:@32238.4]
  input  [63:0] io_ins_128, // @[:@32238.4]
  input  [63:0] io_ins_129, // @[:@32238.4]
  input  [63:0] io_ins_130, // @[:@32238.4]
  input  [63:0] io_ins_131, // @[:@32238.4]
  input  [63:0] io_ins_132, // @[:@32238.4]
  input  [63:0] io_ins_133, // @[:@32238.4]
  input  [63:0] io_ins_134, // @[:@32238.4]
  input  [63:0] io_ins_135, // @[:@32238.4]
  input  [63:0] io_ins_136, // @[:@32238.4]
  input  [63:0] io_ins_137, // @[:@32238.4]
  input  [63:0] io_ins_138, // @[:@32238.4]
  input  [63:0] io_ins_139, // @[:@32238.4]
  input  [63:0] io_ins_140, // @[:@32238.4]
  input  [63:0] io_ins_141, // @[:@32238.4]
  input  [63:0] io_ins_142, // @[:@32238.4]
  input  [63:0] io_ins_143, // @[:@32238.4]
  input  [63:0] io_ins_144, // @[:@32238.4]
  input  [63:0] io_ins_145, // @[:@32238.4]
  input  [63:0] io_ins_146, // @[:@32238.4]
  input  [63:0] io_ins_147, // @[:@32238.4]
  input  [63:0] io_ins_148, // @[:@32238.4]
  input  [63:0] io_ins_149, // @[:@32238.4]
  input  [63:0] io_ins_150, // @[:@32238.4]
  input  [63:0] io_ins_151, // @[:@32238.4]
  input  [63:0] io_ins_152, // @[:@32238.4]
  input  [63:0] io_ins_153, // @[:@32238.4]
  input  [63:0] io_ins_154, // @[:@32238.4]
  input  [63:0] io_ins_155, // @[:@32238.4]
  input  [63:0] io_ins_156, // @[:@32238.4]
  input  [63:0] io_ins_157, // @[:@32238.4]
  input  [63:0] io_ins_158, // @[:@32238.4]
  input  [63:0] io_ins_159, // @[:@32238.4]
  input  [63:0] io_ins_160, // @[:@32238.4]
  input  [63:0] io_ins_161, // @[:@32238.4]
  input  [63:0] io_ins_162, // @[:@32238.4]
  input  [63:0] io_ins_163, // @[:@32238.4]
  input  [63:0] io_ins_164, // @[:@32238.4]
  input  [63:0] io_ins_165, // @[:@32238.4]
  input  [63:0] io_ins_166, // @[:@32238.4]
  input  [63:0] io_ins_167, // @[:@32238.4]
  input  [63:0] io_ins_168, // @[:@32238.4]
  input  [63:0] io_ins_169, // @[:@32238.4]
  input  [63:0] io_ins_170, // @[:@32238.4]
  input  [63:0] io_ins_171, // @[:@32238.4]
  input  [63:0] io_ins_172, // @[:@32238.4]
  input  [63:0] io_ins_173, // @[:@32238.4]
  input  [63:0] io_ins_174, // @[:@32238.4]
  input  [63:0] io_ins_175, // @[:@32238.4]
  input  [63:0] io_ins_176, // @[:@32238.4]
  input  [63:0] io_ins_177, // @[:@32238.4]
  input  [63:0] io_ins_178, // @[:@32238.4]
  input  [63:0] io_ins_179, // @[:@32238.4]
  input  [63:0] io_ins_180, // @[:@32238.4]
  input  [63:0] io_ins_181, // @[:@32238.4]
  input  [63:0] io_ins_182, // @[:@32238.4]
  input  [63:0] io_ins_183, // @[:@32238.4]
  input  [63:0] io_ins_184, // @[:@32238.4]
  input  [63:0] io_ins_185, // @[:@32238.4]
  input  [63:0] io_ins_186, // @[:@32238.4]
  input  [63:0] io_ins_187, // @[:@32238.4]
  input  [63:0] io_ins_188, // @[:@32238.4]
  input  [63:0] io_ins_189, // @[:@32238.4]
  input  [63:0] io_ins_190, // @[:@32238.4]
  input  [63:0] io_ins_191, // @[:@32238.4]
  input  [63:0] io_ins_192, // @[:@32238.4]
  input  [63:0] io_ins_193, // @[:@32238.4]
  input  [63:0] io_ins_194, // @[:@32238.4]
  input  [63:0] io_ins_195, // @[:@32238.4]
  input  [63:0] io_ins_196, // @[:@32238.4]
  input  [63:0] io_ins_197, // @[:@32238.4]
  input  [63:0] io_ins_198, // @[:@32238.4]
  input  [63:0] io_ins_199, // @[:@32238.4]
  input  [63:0] io_ins_200, // @[:@32238.4]
  input  [63:0] io_ins_201, // @[:@32238.4]
  input  [63:0] io_ins_202, // @[:@32238.4]
  input  [63:0] io_ins_203, // @[:@32238.4]
  input  [63:0] io_ins_204, // @[:@32238.4]
  input  [63:0] io_ins_205, // @[:@32238.4]
  input  [63:0] io_ins_206, // @[:@32238.4]
  input  [63:0] io_ins_207, // @[:@32238.4]
  input  [63:0] io_ins_208, // @[:@32238.4]
  input  [63:0] io_ins_209, // @[:@32238.4]
  input  [63:0] io_ins_210, // @[:@32238.4]
  input  [63:0] io_ins_211, // @[:@32238.4]
  input  [63:0] io_ins_212, // @[:@32238.4]
  input  [63:0] io_ins_213, // @[:@32238.4]
  input  [63:0] io_ins_214, // @[:@32238.4]
  input  [63:0] io_ins_215, // @[:@32238.4]
  input  [63:0] io_ins_216, // @[:@32238.4]
  input  [63:0] io_ins_217, // @[:@32238.4]
  input  [63:0] io_ins_218, // @[:@32238.4]
  input  [63:0] io_ins_219, // @[:@32238.4]
  input  [63:0] io_ins_220, // @[:@32238.4]
  input  [63:0] io_ins_221, // @[:@32238.4]
  input  [63:0] io_ins_222, // @[:@32238.4]
  input  [63:0] io_ins_223, // @[:@32238.4]
  input  [63:0] io_ins_224, // @[:@32238.4]
  input  [63:0] io_ins_225, // @[:@32238.4]
  input  [63:0] io_ins_226, // @[:@32238.4]
  input  [63:0] io_ins_227, // @[:@32238.4]
  input  [63:0] io_ins_228, // @[:@32238.4]
  input  [63:0] io_ins_229, // @[:@32238.4]
  input  [63:0] io_ins_230, // @[:@32238.4]
  input  [63:0] io_ins_231, // @[:@32238.4]
  input  [63:0] io_ins_232, // @[:@32238.4]
  input  [63:0] io_ins_233, // @[:@32238.4]
  input  [63:0] io_ins_234, // @[:@32238.4]
  input  [63:0] io_ins_235, // @[:@32238.4]
  input  [63:0] io_ins_236, // @[:@32238.4]
  input  [63:0] io_ins_237, // @[:@32238.4]
  input  [63:0] io_ins_238, // @[:@32238.4]
  input  [63:0] io_ins_239, // @[:@32238.4]
  input  [63:0] io_ins_240, // @[:@32238.4]
  input  [63:0] io_ins_241, // @[:@32238.4]
  input  [63:0] io_ins_242, // @[:@32238.4]
  input  [63:0] io_ins_243, // @[:@32238.4]
  input  [63:0] io_ins_244, // @[:@32238.4]
  input  [63:0] io_ins_245, // @[:@32238.4]
  input  [63:0] io_ins_246, // @[:@32238.4]
  input  [63:0] io_ins_247, // @[:@32238.4]
  input  [63:0] io_ins_248, // @[:@32238.4]
  input  [63:0] io_ins_249, // @[:@32238.4]
  input  [63:0] io_ins_250, // @[:@32238.4]
  input  [63:0] io_ins_251, // @[:@32238.4]
  input  [63:0] io_ins_252, // @[:@32238.4]
  input  [63:0] io_ins_253, // @[:@32238.4]
  input  [63:0] io_ins_254, // @[:@32238.4]
  input  [63:0] io_ins_255, // @[:@32238.4]
  input  [63:0] io_ins_256, // @[:@32238.4]
  input  [63:0] io_ins_257, // @[:@32238.4]
  input  [63:0] io_ins_258, // @[:@32238.4]
  input  [63:0] io_ins_259, // @[:@32238.4]
  input  [63:0] io_ins_260, // @[:@32238.4]
  input  [63:0] io_ins_261, // @[:@32238.4]
  input  [63:0] io_ins_262, // @[:@32238.4]
  input  [63:0] io_ins_263, // @[:@32238.4]
  input  [63:0] io_ins_264, // @[:@32238.4]
  input  [63:0] io_ins_265, // @[:@32238.4]
  input  [63:0] io_ins_266, // @[:@32238.4]
  input  [63:0] io_ins_267, // @[:@32238.4]
  input  [63:0] io_ins_268, // @[:@32238.4]
  input  [63:0] io_ins_269, // @[:@32238.4]
  input  [63:0] io_ins_270, // @[:@32238.4]
  input  [63:0] io_ins_271, // @[:@32238.4]
  input  [63:0] io_ins_272, // @[:@32238.4]
  input  [63:0] io_ins_273, // @[:@32238.4]
  input  [63:0] io_ins_274, // @[:@32238.4]
  input  [63:0] io_ins_275, // @[:@32238.4]
  input  [63:0] io_ins_276, // @[:@32238.4]
  input  [63:0] io_ins_277, // @[:@32238.4]
  input  [63:0] io_ins_278, // @[:@32238.4]
  input  [63:0] io_ins_279, // @[:@32238.4]
  input  [63:0] io_ins_280, // @[:@32238.4]
  input  [63:0] io_ins_281, // @[:@32238.4]
  input  [63:0] io_ins_282, // @[:@32238.4]
  input  [63:0] io_ins_283, // @[:@32238.4]
  input  [63:0] io_ins_284, // @[:@32238.4]
  input  [63:0] io_ins_285, // @[:@32238.4]
  input  [63:0] io_ins_286, // @[:@32238.4]
  input  [63:0] io_ins_287, // @[:@32238.4]
  input  [63:0] io_ins_288, // @[:@32238.4]
  input  [63:0] io_ins_289, // @[:@32238.4]
  input  [63:0] io_ins_290, // @[:@32238.4]
  input  [63:0] io_ins_291, // @[:@32238.4]
  input  [63:0] io_ins_292, // @[:@32238.4]
  input  [63:0] io_ins_293, // @[:@32238.4]
  input  [63:0] io_ins_294, // @[:@32238.4]
  input  [63:0] io_ins_295, // @[:@32238.4]
  input  [63:0] io_ins_296, // @[:@32238.4]
  input  [63:0] io_ins_297, // @[:@32238.4]
  input  [63:0] io_ins_298, // @[:@32238.4]
  input  [63:0] io_ins_299, // @[:@32238.4]
  input  [63:0] io_ins_300, // @[:@32238.4]
  input  [63:0] io_ins_301, // @[:@32238.4]
  input  [63:0] io_ins_302, // @[:@32238.4]
  input  [63:0] io_ins_303, // @[:@32238.4]
  input  [63:0] io_ins_304, // @[:@32238.4]
  input  [63:0] io_ins_305, // @[:@32238.4]
  input  [63:0] io_ins_306, // @[:@32238.4]
  input  [63:0] io_ins_307, // @[:@32238.4]
  input  [63:0] io_ins_308, // @[:@32238.4]
  input  [63:0] io_ins_309, // @[:@32238.4]
  input  [63:0] io_ins_310, // @[:@32238.4]
  input  [63:0] io_ins_311, // @[:@32238.4]
  input  [63:0] io_ins_312, // @[:@32238.4]
  input  [63:0] io_ins_313, // @[:@32238.4]
  input  [63:0] io_ins_314, // @[:@32238.4]
  input  [63:0] io_ins_315, // @[:@32238.4]
  input  [63:0] io_ins_316, // @[:@32238.4]
  input  [63:0] io_ins_317, // @[:@32238.4]
  input  [63:0] io_ins_318, // @[:@32238.4]
  input  [63:0] io_ins_319, // @[:@32238.4]
  input  [63:0] io_ins_320, // @[:@32238.4]
  input  [63:0] io_ins_321, // @[:@32238.4]
  input  [63:0] io_ins_322, // @[:@32238.4]
  input  [63:0] io_ins_323, // @[:@32238.4]
  input  [63:0] io_ins_324, // @[:@32238.4]
  input  [63:0] io_ins_325, // @[:@32238.4]
  input  [63:0] io_ins_326, // @[:@32238.4]
  input  [63:0] io_ins_327, // @[:@32238.4]
  input  [63:0] io_ins_328, // @[:@32238.4]
  input  [63:0] io_ins_329, // @[:@32238.4]
  input  [63:0] io_ins_330, // @[:@32238.4]
  input  [63:0] io_ins_331, // @[:@32238.4]
  input  [63:0] io_ins_332, // @[:@32238.4]
  input  [63:0] io_ins_333, // @[:@32238.4]
  input  [63:0] io_ins_334, // @[:@32238.4]
  input  [63:0] io_ins_335, // @[:@32238.4]
  input  [63:0] io_ins_336, // @[:@32238.4]
  input  [63:0] io_ins_337, // @[:@32238.4]
  input  [63:0] io_ins_338, // @[:@32238.4]
  input  [63:0] io_ins_339, // @[:@32238.4]
  input  [63:0] io_ins_340, // @[:@32238.4]
  input  [63:0] io_ins_341, // @[:@32238.4]
  input  [63:0] io_ins_342, // @[:@32238.4]
  input  [63:0] io_ins_343, // @[:@32238.4]
  input  [63:0] io_ins_344, // @[:@32238.4]
  input  [63:0] io_ins_345, // @[:@32238.4]
  input  [63:0] io_ins_346, // @[:@32238.4]
  input  [63:0] io_ins_347, // @[:@32238.4]
  input  [63:0] io_ins_348, // @[:@32238.4]
  input  [63:0] io_ins_349, // @[:@32238.4]
  input  [63:0] io_ins_350, // @[:@32238.4]
  input  [63:0] io_ins_351, // @[:@32238.4]
  input  [63:0] io_ins_352, // @[:@32238.4]
  input  [63:0] io_ins_353, // @[:@32238.4]
  input  [63:0] io_ins_354, // @[:@32238.4]
  input  [63:0] io_ins_355, // @[:@32238.4]
  input  [63:0] io_ins_356, // @[:@32238.4]
  input  [63:0] io_ins_357, // @[:@32238.4]
  input  [63:0] io_ins_358, // @[:@32238.4]
  input  [63:0] io_ins_359, // @[:@32238.4]
  input  [63:0] io_ins_360, // @[:@32238.4]
  input  [63:0] io_ins_361, // @[:@32238.4]
  input  [63:0] io_ins_362, // @[:@32238.4]
  input  [63:0] io_ins_363, // @[:@32238.4]
  input  [63:0] io_ins_364, // @[:@32238.4]
  input  [63:0] io_ins_365, // @[:@32238.4]
  input  [63:0] io_ins_366, // @[:@32238.4]
  input  [63:0] io_ins_367, // @[:@32238.4]
  input  [63:0] io_ins_368, // @[:@32238.4]
  input  [63:0] io_ins_369, // @[:@32238.4]
  input  [63:0] io_ins_370, // @[:@32238.4]
  input  [63:0] io_ins_371, // @[:@32238.4]
  input  [63:0] io_ins_372, // @[:@32238.4]
  input  [63:0] io_ins_373, // @[:@32238.4]
  input  [63:0] io_ins_374, // @[:@32238.4]
  input  [63:0] io_ins_375, // @[:@32238.4]
  input  [63:0] io_ins_376, // @[:@32238.4]
  input  [63:0] io_ins_377, // @[:@32238.4]
  input  [63:0] io_ins_378, // @[:@32238.4]
  input  [63:0] io_ins_379, // @[:@32238.4]
  input  [63:0] io_ins_380, // @[:@32238.4]
  input  [63:0] io_ins_381, // @[:@32238.4]
  input  [63:0] io_ins_382, // @[:@32238.4]
  input  [63:0] io_ins_383, // @[:@32238.4]
  input  [63:0] io_ins_384, // @[:@32238.4]
  input  [63:0] io_ins_385, // @[:@32238.4]
  input  [63:0] io_ins_386, // @[:@32238.4]
  input  [63:0] io_ins_387, // @[:@32238.4]
  input  [63:0] io_ins_388, // @[:@32238.4]
  input  [63:0] io_ins_389, // @[:@32238.4]
  input  [63:0] io_ins_390, // @[:@32238.4]
  input  [63:0] io_ins_391, // @[:@32238.4]
  input  [63:0] io_ins_392, // @[:@32238.4]
  input  [63:0] io_ins_393, // @[:@32238.4]
  input  [63:0] io_ins_394, // @[:@32238.4]
  input  [63:0] io_ins_395, // @[:@32238.4]
  input  [63:0] io_ins_396, // @[:@32238.4]
  input  [63:0] io_ins_397, // @[:@32238.4]
  input  [63:0] io_ins_398, // @[:@32238.4]
  input  [63:0] io_ins_399, // @[:@32238.4]
  input  [63:0] io_ins_400, // @[:@32238.4]
  input  [63:0] io_ins_401, // @[:@32238.4]
  input  [63:0] io_ins_402, // @[:@32238.4]
  input  [63:0] io_ins_403, // @[:@32238.4]
  input  [63:0] io_ins_404, // @[:@32238.4]
  input  [63:0] io_ins_405, // @[:@32238.4]
  input  [63:0] io_ins_406, // @[:@32238.4]
  input  [63:0] io_ins_407, // @[:@32238.4]
  input  [63:0] io_ins_408, // @[:@32238.4]
  input  [63:0] io_ins_409, // @[:@32238.4]
  input  [63:0] io_ins_410, // @[:@32238.4]
  input  [63:0] io_ins_411, // @[:@32238.4]
  input  [63:0] io_ins_412, // @[:@32238.4]
  input  [63:0] io_ins_413, // @[:@32238.4]
  input  [63:0] io_ins_414, // @[:@32238.4]
  input  [63:0] io_ins_415, // @[:@32238.4]
  input  [63:0] io_ins_416, // @[:@32238.4]
  input  [63:0] io_ins_417, // @[:@32238.4]
  input  [63:0] io_ins_418, // @[:@32238.4]
  input  [63:0] io_ins_419, // @[:@32238.4]
  input  [63:0] io_ins_420, // @[:@32238.4]
  input  [63:0] io_ins_421, // @[:@32238.4]
  input  [63:0] io_ins_422, // @[:@32238.4]
  input  [63:0] io_ins_423, // @[:@32238.4]
  input  [63:0] io_ins_424, // @[:@32238.4]
  input  [63:0] io_ins_425, // @[:@32238.4]
  input  [63:0] io_ins_426, // @[:@32238.4]
  input  [63:0] io_ins_427, // @[:@32238.4]
  input  [63:0] io_ins_428, // @[:@32238.4]
  input  [63:0] io_ins_429, // @[:@32238.4]
  input  [63:0] io_ins_430, // @[:@32238.4]
  input  [63:0] io_ins_431, // @[:@32238.4]
  input  [63:0] io_ins_432, // @[:@32238.4]
  input  [63:0] io_ins_433, // @[:@32238.4]
  input  [63:0] io_ins_434, // @[:@32238.4]
  input  [63:0] io_ins_435, // @[:@32238.4]
  input  [63:0] io_ins_436, // @[:@32238.4]
  input  [63:0] io_ins_437, // @[:@32238.4]
  input  [63:0] io_ins_438, // @[:@32238.4]
  input  [63:0] io_ins_439, // @[:@32238.4]
  input  [63:0] io_ins_440, // @[:@32238.4]
  input  [63:0] io_ins_441, // @[:@32238.4]
  input  [63:0] io_ins_442, // @[:@32238.4]
  input  [63:0] io_ins_443, // @[:@32238.4]
  input  [63:0] io_ins_444, // @[:@32238.4]
  input  [63:0] io_ins_445, // @[:@32238.4]
  input  [63:0] io_ins_446, // @[:@32238.4]
  input  [63:0] io_ins_447, // @[:@32238.4]
  input  [63:0] io_ins_448, // @[:@32238.4]
  input  [63:0] io_ins_449, // @[:@32238.4]
  input  [63:0] io_ins_450, // @[:@32238.4]
  input  [63:0] io_ins_451, // @[:@32238.4]
  input  [63:0] io_ins_452, // @[:@32238.4]
  input  [63:0] io_ins_453, // @[:@32238.4]
  input  [63:0] io_ins_454, // @[:@32238.4]
  input  [63:0] io_ins_455, // @[:@32238.4]
  input  [63:0] io_ins_456, // @[:@32238.4]
  input  [63:0] io_ins_457, // @[:@32238.4]
  input  [63:0] io_ins_458, // @[:@32238.4]
  input  [63:0] io_ins_459, // @[:@32238.4]
  input  [63:0] io_ins_460, // @[:@32238.4]
  input  [63:0] io_ins_461, // @[:@32238.4]
  input  [63:0] io_ins_462, // @[:@32238.4]
  input  [63:0] io_ins_463, // @[:@32238.4]
  input  [63:0] io_ins_464, // @[:@32238.4]
  input  [63:0] io_ins_465, // @[:@32238.4]
  input  [63:0] io_ins_466, // @[:@32238.4]
  input  [63:0] io_ins_467, // @[:@32238.4]
  input  [63:0] io_ins_468, // @[:@32238.4]
  input  [63:0] io_ins_469, // @[:@32238.4]
  input  [63:0] io_ins_470, // @[:@32238.4]
  input  [63:0] io_ins_471, // @[:@32238.4]
  input  [63:0] io_ins_472, // @[:@32238.4]
  input  [63:0] io_ins_473, // @[:@32238.4]
  input  [63:0] io_ins_474, // @[:@32238.4]
  input  [63:0] io_ins_475, // @[:@32238.4]
  input  [63:0] io_ins_476, // @[:@32238.4]
  input  [63:0] io_ins_477, // @[:@32238.4]
  input  [63:0] io_ins_478, // @[:@32238.4]
  input  [63:0] io_ins_479, // @[:@32238.4]
  input  [63:0] io_ins_480, // @[:@32238.4]
  input  [63:0] io_ins_481, // @[:@32238.4]
  input  [63:0] io_ins_482, // @[:@32238.4]
  input  [63:0] io_ins_483, // @[:@32238.4]
  input  [63:0] io_ins_484, // @[:@32238.4]
  input  [63:0] io_ins_485, // @[:@32238.4]
  input  [63:0] io_ins_486, // @[:@32238.4]
  input  [63:0] io_ins_487, // @[:@32238.4]
  input  [63:0] io_ins_488, // @[:@32238.4]
  input  [63:0] io_ins_489, // @[:@32238.4]
  input  [63:0] io_ins_490, // @[:@32238.4]
  input  [63:0] io_ins_491, // @[:@32238.4]
  input  [63:0] io_ins_492, // @[:@32238.4]
  input  [63:0] io_ins_493, // @[:@32238.4]
  input  [63:0] io_ins_494, // @[:@32238.4]
  input  [63:0] io_ins_495, // @[:@32238.4]
  input  [63:0] io_ins_496, // @[:@32238.4]
  input  [63:0] io_ins_497, // @[:@32238.4]
  input  [63:0] io_ins_498, // @[:@32238.4]
  input  [63:0] io_ins_499, // @[:@32238.4]
  input  [63:0] io_ins_500, // @[:@32238.4]
  input  [63:0] io_ins_501, // @[:@32238.4]
  input  [63:0] io_ins_502, // @[:@32238.4]
  input  [8:0]  io_sel, // @[:@32238.4]
  output [63:0] io_out // @[:@32238.4]
);
  wire [63:0] _GEN_1; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_2; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_3; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_4; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_5; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_6; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_7; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_8; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_9; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_10; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_11; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_12; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_13; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_14; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_15; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_16; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_17; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_18; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_19; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_20; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_21; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_22; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_23; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_24; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_25; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_26; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_27; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_28; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_29; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_30; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_31; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_32; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_33; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_34; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_35; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_36; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_37; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_38; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_39; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_40; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_41; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_42; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_43; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_44; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_45; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_46; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_47; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_48; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_49; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_50; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_51; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_52; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_53; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_54; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_55; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_56; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_57; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_58; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_59; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_60; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_61; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_62; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_63; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_64; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_65; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_66; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_67; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_68; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_69; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_70; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_71; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_72; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_73; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_74; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_75; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_76; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_77; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_78; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_79; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_80; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_81; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_82; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_83; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_84; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_85; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_86; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_87; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_88; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_89; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_90; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_91; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_92; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_93; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_94; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_95; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_96; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_97; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_98; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_99; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_100; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_101; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_102; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_103; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_104; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_105; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_106; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_107; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_108; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_109; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_110; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_111; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_112; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_113; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_114; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_115; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_116; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_117; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_118; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_119; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_120; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_121; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_122; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_123; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_124; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_125; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_126; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_127; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_128; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_129; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_130; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_131; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_132; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_133; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_134; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_135; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_136; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_137; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_138; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_139; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_140; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_141; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_142; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_143; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_144; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_145; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_146; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_147; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_148; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_149; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_150; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_151; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_152; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_153; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_154; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_155; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_156; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_157; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_158; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_159; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_160; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_161; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_162; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_163; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_164; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_165; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_166; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_167; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_168; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_169; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_170; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_171; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_172; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_173; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_174; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_175; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_176; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_177; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_178; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_179; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_180; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_181; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_182; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_183; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_184; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_185; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_186; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_187; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_188; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_189; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_190; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_191; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_192; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_193; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_194; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_195; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_196; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_197; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_198; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_199; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_200; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_201; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_202; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_203; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_204; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_205; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_206; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_207; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_208; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_209; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_210; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_211; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_212; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_213; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_214; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_215; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_216; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_217; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_218; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_219; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_220; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_221; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_222; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_223; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_224; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_225; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_226; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_227; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_228; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_229; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_230; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_231; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_232; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_233; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_234; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_235; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_236; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_237; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_238; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_239; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_240; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_241; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_242; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_243; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_244; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_245; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_246; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_247; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_248; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_249; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_250; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_251; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_252; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_253; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_254; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_255; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_256; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_257; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_258; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_259; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_260; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_261; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_262; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_263; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_264; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_265; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_266; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_267; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_268; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_269; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_270; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_271; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_272; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_273; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_274; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_275; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_276; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_277; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_278; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_279; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_280; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_281; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_282; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_283; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_284; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_285; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_286; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_287; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_288; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_289; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_290; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_291; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_292; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_293; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_294; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_295; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_296; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_297; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_298; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_299; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_300; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_301; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_302; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_303; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_304; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_305; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_306; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_307; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_308; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_309; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_310; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_311; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_312; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_313; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_314; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_315; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_316; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_317; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_318; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_319; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_320; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_321; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_322; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_323; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_324; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_325; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_326; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_327; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_328; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_329; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_330; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_331; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_332; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_333; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_334; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_335; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_336; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_337; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_338; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_339; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_340; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_341; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_342; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_343; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_344; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_345; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_346; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_347; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_348; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_349; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_350; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_351; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_352; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_353; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_354; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_355; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_356; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_357; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_358; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_359; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_360; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_361; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_362; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_363; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_364; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_365; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_366; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_367; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_368; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_369; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_370; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_371; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_372; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_373; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_374; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_375; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_376; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_377; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_378; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_379; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_380; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_381; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_382; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_383; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_384; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_385; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_386; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_387; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_388; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_389; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_390; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_391; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_392; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_393; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_394; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_395; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_396; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_397; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_398; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_399; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_400; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_401; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_402; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_403; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_404; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_405; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_406; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_407; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_408; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_409; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_410; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_411; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_412; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_413; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_414; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_415; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_416; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_417; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_418; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_419; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_420; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_421; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_422; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_423; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_424; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_425; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_426; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_427; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_428; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_429; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_430; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_431; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_432; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_433; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_434; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_435; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_436; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_437; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_438; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_439; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_440; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_441; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_442; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_443; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_444; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_445; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_446; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_447; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_448; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_449; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_450; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_451; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_452; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_453; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_454; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_455; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_456; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_457; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_458; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_459; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_460; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_461; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_462; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_463; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_464; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_465; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_466; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_467; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_468; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_469; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_470; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_471; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_472; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_473; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_474; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_475; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_476; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_477; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_478; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_479; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_480; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_481; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_482; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_483; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_484; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_485; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_486; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_487; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_488; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_489; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_490; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_491; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_492; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_493; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_494; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_495; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_496; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_497; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_498; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_499; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_500; // @[MuxN.scala 16:10:@32240.4]
  wire [63:0] _GEN_501; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_1 = 9'h1 == io_sel ? io_ins_1 : io_ins_0; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_2 = 9'h2 == io_sel ? io_ins_2 : _GEN_1; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_3 = 9'h3 == io_sel ? io_ins_3 : _GEN_2; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_4 = 9'h4 == io_sel ? io_ins_4 : _GEN_3; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_5 = 9'h5 == io_sel ? io_ins_5 : _GEN_4; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_6 = 9'h6 == io_sel ? io_ins_6 : _GEN_5; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_7 = 9'h7 == io_sel ? io_ins_7 : _GEN_6; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_8 = 9'h8 == io_sel ? io_ins_8 : _GEN_7; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_9 = 9'h9 == io_sel ? io_ins_9 : _GEN_8; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_10 = 9'ha == io_sel ? io_ins_10 : _GEN_9; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_11 = 9'hb == io_sel ? io_ins_11 : _GEN_10; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_12 = 9'hc == io_sel ? io_ins_12 : _GEN_11; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_13 = 9'hd == io_sel ? io_ins_13 : _GEN_12; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_14 = 9'he == io_sel ? io_ins_14 : _GEN_13; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_15 = 9'hf == io_sel ? io_ins_15 : _GEN_14; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_16 = 9'h10 == io_sel ? io_ins_16 : _GEN_15; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_17 = 9'h11 == io_sel ? io_ins_17 : _GEN_16; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_18 = 9'h12 == io_sel ? io_ins_18 : _GEN_17; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_19 = 9'h13 == io_sel ? io_ins_19 : _GEN_18; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_20 = 9'h14 == io_sel ? io_ins_20 : _GEN_19; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_21 = 9'h15 == io_sel ? io_ins_21 : _GEN_20; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_22 = 9'h16 == io_sel ? io_ins_22 : _GEN_21; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_23 = 9'h17 == io_sel ? io_ins_23 : _GEN_22; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_24 = 9'h18 == io_sel ? io_ins_24 : _GEN_23; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_25 = 9'h19 == io_sel ? io_ins_25 : _GEN_24; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_26 = 9'h1a == io_sel ? io_ins_26 : _GEN_25; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_27 = 9'h1b == io_sel ? io_ins_27 : _GEN_26; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_28 = 9'h1c == io_sel ? io_ins_28 : _GEN_27; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_29 = 9'h1d == io_sel ? io_ins_29 : _GEN_28; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_30 = 9'h1e == io_sel ? io_ins_30 : _GEN_29; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_31 = 9'h1f == io_sel ? io_ins_31 : _GEN_30; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_32 = 9'h20 == io_sel ? io_ins_32 : _GEN_31; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_33 = 9'h21 == io_sel ? io_ins_33 : _GEN_32; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_34 = 9'h22 == io_sel ? io_ins_34 : _GEN_33; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_35 = 9'h23 == io_sel ? io_ins_35 : _GEN_34; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_36 = 9'h24 == io_sel ? io_ins_36 : _GEN_35; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_37 = 9'h25 == io_sel ? io_ins_37 : _GEN_36; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_38 = 9'h26 == io_sel ? io_ins_38 : _GEN_37; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_39 = 9'h27 == io_sel ? io_ins_39 : _GEN_38; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_40 = 9'h28 == io_sel ? io_ins_40 : _GEN_39; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_41 = 9'h29 == io_sel ? io_ins_41 : _GEN_40; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_42 = 9'h2a == io_sel ? io_ins_42 : _GEN_41; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_43 = 9'h2b == io_sel ? io_ins_43 : _GEN_42; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_44 = 9'h2c == io_sel ? io_ins_44 : _GEN_43; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_45 = 9'h2d == io_sel ? io_ins_45 : _GEN_44; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_46 = 9'h2e == io_sel ? io_ins_46 : _GEN_45; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_47 = 9'h2f == io_sel ? io_ins_47 : _GEN_46; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_48 = 9'h30 == io_sel ? io_ins_48 : _GEN_47; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_49 = 9'h31 == io_sel ? io_ins_49 : _GEN_48; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_50 = 9'h32 == io_sel ? io_ins_50 : _GEN_49; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_51 = 9'h33 == io_sel ? io_ins_51 : _GEN_50; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_52 = 9'h34 == io_sel ? io_ins_52 : _GEN_51; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_53 = 9'h35 == io_sel ? io_ins_53 : _GEN_52; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_54 = 9'h36 == io_sel ? io_ins_54 : _GEN_53; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_55 = 9'h37 == io_sel ? io_ins_55 : _GEN_54; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_56 = 9'h38 == io_sel ? io_ins_56 : _GEN_55; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_57 = 9'h39 == io_sel ? io_ins_57 : _GEN_56; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_58 = 9'h3a == io_sel ? io_ins_58 : _GEN_57; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_59 = 9'h3b == io_sel ? io_ins_59 : _GEN_58; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_60 = 9'h3c == io_sel ? io_ins_60 : _GEN_59; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_61 = 9'h3d == io_sel ? io_ins_61 : _GEN_60; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_62 = 9'h3e == io_sel ? io_ins_62 : _GEN_61; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_63 = 9'h3f == io_sel ? io_ins_63 : _GEN_62; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_64 = 9'h40 == io_sel ? io_ins_64 : _GEN_63; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_65 = 9'h41 == io_sel ? io_ins_65 : _GEN_64; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_66 = 9'h42 == io_sel ? io_ins_66 : _GEN_65; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_67 = 9'h43 == io_sel ? io_ins_67 : _GEN_66; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_68 = 9'h44 == io_sel ? io_ins_68 : _GEN_67; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_69 = 9'h45 == io_sel ? io_ins_69 : _GEN_68; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_70 = 9'h46 == io_sel ? io_ins_70 : _GEN_69; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_71 = 9'h47 == io_sel ? io_ins_71 : _GEN_70; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_72 = 9'h48 == io_sel ? io_ins_72 : _GEN_71; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_73 = 9'h49 == io_sel ? io_ins_73 : _GEN_72; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_74 = 9'h4a == io_sel ? io_ins_74 : _GEN_73; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_75 = 9'h4b == io_sel ? io_ins_75 : _GEN_74; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_76 = 9'h4c == io_sel ? io_ins_76 : _GEN_75; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_77 = 9'h4d == io_sel ? io_ins_77 : _GEN_76; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_78 = 9'h4e == io_sel ? io_ins_78 : _GEN_77; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_79 = 9'h4f == io_sel ? io_ins_79 : _GEN_78; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_80 = 9'h50 == io_sel ? io_ins_80 : _GEN_79; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_81 = 9'h51 == io_sel ? io_ins_81 : _GEN_80; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_82 = 9'h52 == io_sel ? io_ins_82 : _GEN_81; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_83 = 9'h53 == io_sel ? io_ins_83 : _GEN_82; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_84 = 9'h54 == io_sel ? io_ins_84 : _GEN_83; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_85 = 9'h55 == io_sel ? io_ins_85 : _GEN_84; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_86 = 9'h56 == io_sel ? io_ins_86 : _GEN_85; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_87 = 9'h57 == io_sel ? io_ins_87 : _GEN_86; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_88 = 9'h58 == io_sel ? io_ins_88 : _GEN_87; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_89 = 9'h59 == io_sel ? io_ins_89 : _GEN_88; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_90 = 9'h5a == io_sel ? io_ins_90 : _GEN_89; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_91 = 9'h5b == io_sel ? io_ins_91 : _GEN_90; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_92 = 9'h5c == io_sel ? io_ins_92 : _GEN_91; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_93 = 9'h5d == io_sel ? io_ins_93 : _GEN_92; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_94 = 9'h5e == io_sel ? io_ins_94 : _GEN_93; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_95 = 9'h5f == io_sel ? io_ins_95 : _GEN_94; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_96 = 9'h60 == io_sel ? io_ins_96 : _GEN_95; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_97 = 9'h61 == io_sel ? io_ins_97 : _GEN_96; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_98 = 9'h62 == io_sel ? io_ins_98 : _GEN_97; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_99 = 9'h63 == io_sel ? io_ins_99 : _GEN_98; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_100 = 9'h64 == io_sel ? io_ins_100 : _GEN_99; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_101 = 9'h65 == io_sel ? io_ins_101 : _GEN_100; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_102 = 9'h66 == io_sel ? io_ins_102 : _GEN_101; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_103 = 9'h67 == io_sel ? io_ins_103 : _GEN_102; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_104 = 9'h68 == io_sel ? io_ins_104 : _GEN_103; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_105 = 9'h69 == io_sel ? io_ins_105 : _GEN_104; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_106 = 9'h6a == io_sel ? io_ins_106 : _GEN_105; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_107 = 9'h6b == io_sel ? io_ins_107 : _GEN_106; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_108 = 9'h6c == io_sel ? io_ins_108 : _GEN_107; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_109 = 9'h6d == io_sel ? io_ins_109 : _GEN_108; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_110 = 9'h6e == io_sel ? io_ins_110 : _GEN_109; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_111 = 9'h6f == io_sel ? io_ins_111 : _GEN_110; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_112 = 9'h70 == io_sel ? io_ins_112 : _GEN_111; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_113 = 9'h71 == io_sel ? io_ins_113 : _GEN_112; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_114 = 9'h72 == io_sel ? io_ins_114 : _GEN_113; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_115 = 9'h73 == io_sel ? io_ins_115 : _GEN_114; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_116 = 9'h74 == io_sel ? io_ins_116 : _GEN_115; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_117 = 9'h75 == io_sel ? io_ins_117 : _GEN_116; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_118 = 9'h76 == io_sel ? io_ins_118 : _GEN_117; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_119 = 9'h77 == io_sel ? io_ins_119 : _GEN_118; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_120 = 9'h78 == io_sel ? io_ins_120 : _GEN_119; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_121 = 9'h79 == io_sel ? io_ins_121 : _GEN_120; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_122 = 9'h7a == io_sel ? io_ins_122 : _GEN_121; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_123 = 9'h7b == io_sel ? io_ins_123 : _GEN_122; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_124 = 9'h7c == io_sel ? io_ins_124 : _GEN_123; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_125 = 9'h7d == io_sel ? io_ins_125 : _GEN_124; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_126 = 9'h7e == io_sel ? io_ins_126 : _GEN_125; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_127 = 9'h7f == io_sel ? io_ins_127 : _GEN_126; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_128 = 9'h80 == io_sel ? io_ins_128 : _GEN_127; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_129 = 9'h81 == io_sel ? io_ins_129 : _GEN_128; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_130 = 9'h82 == io_sel ? io_ins_130 : _GEN_129; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_131 = 9'h83 == io_sel ? io_ins_131 : _GEN_130; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_132 = 9'h84 == io_sel ? io_ins_132 : _GEN_131; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_133 = 9'h85 == io_sel ? io_ins_133 : _GEN_132; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_134 = 9'h86 == io_sel ? io_ins_134 : _GEN_133; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_135 = 9'h87 == io_sel ? io_ins_135 : _GEN_134; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_136 = 9'h88 == io_sel ? io_ins_136 : _GEN_135; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_137 = 9'h89 == io_sel ? io_ins_137 : _GEN_136; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_138 = 9'h8a == io_sel ? io_ins_138 : _GEN_137; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_139 = 9'h8b == io_sel ? io_ins_139 : _GEN_138; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_140 = 9'h8c == io_sel ? io_ins_140 : _GEN_139; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_141 = 9'h8d == io_sel ? io_ins_141 : _GEN_140; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_142 = 9'h8e == io_sel ? io_ins_142 : _GEN_141; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_143 = 9'h8f == io_sel ? io_ins_143 : _GEN_142; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_144 = 9'h90 == io_sel ? io_ins_144 : _GEN_143; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_145 = 9'h91 == io_sel ? io_ins_145 : _GEN_144; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_146 = 9'h92 == io_sel ? io_ins_146 : _GEN_145; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_147 = 9'h93 == io_sel ? io_ins_147 : _GEN_146; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_148 = 9'h94 == io_sel ? io_ins_148 : _GEN_147; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_149 = 9'h95 == io_sel ? io_ins_149 : _GEN_148; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_150 = 9'h96 == io_sel ? io_ins_150 : _GEN_149; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_151 = 9'h97 == io_sel ? io_ins_151 : _GEN_150; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_152 = 9'h98 == io_sel ? io_ins_152 : _GEN_151; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_153 = 9'h99 == io_sel ? io_ins_153 : _GEN_152; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_154 = 9'h9a == io_sel ? io_ins_154 : _GEN_153; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_155 = 9'h9b == io_sel ? io_ins_155 : _GEN_154; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_156 = 9'h9c == io_sel ? io_ins_156 : _GEN_155; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_157 = 9'h9d == io_sel ? io_ins_157 : _GEN_156; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_158 = 9'h9e == io_sel ? io_ins_158 : _GEN_157; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_159 = 9'h9f == io_sel ? io_ins_159 : _GEN_158; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_160 = 9'ha0 == io_sel ? io_ins_160 : _GEN_159; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_161 = 9'ha1 == io_sel ? io_ins_161 : _GEN_160; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_162 = 9'ha2 == io_sel ? io_ins_162 : _GEN_161; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_163 = 9'ha3 == io_sel ? io_ins_163 : _GEN_162; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_164 = 9'ha4 == io_sel ? io_ins_164 : _GEN_163; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_165 = 9'ha5 == io_sel ? io_ins_165 : _GEN_164; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_166 = 9'ha6 == io_sel ? io_ins_166 : _GEN_165; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_167 = 9'ha7 == io_sel ? io_ins_167 : _GEN_166; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_168 = 9'ha8 == io_sel ? io_ins_168 : _GEN_167; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_169 = 9'ha9 == io_sel ? io_ins_169 : _GEN_168; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_170 = 9'haa == io_sel ? io_ins_170 : _GEN_169; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_171 = 9'hab == io_sel ? io_ins_171 : _GEN_170; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_172 = 9'hac == io_sel ? io_ins_172 : _GEN_171; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_173 = 9'had == io_sel ? io_ins_173 : _GEN_172; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_174 = 9'hae == io_sel ? io_ins_174 : _GEN_173; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_175 = 9'haf == io_sel ? io_ins_175 : _GEN_174; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_176 = 9'hb0 == io_sel ? io_ins_176 : _GEN_175; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_177 = 9'hb1 == io_sel ? io_ins_177 : _GEN_176; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_178 = 9'hb2 == io_sel ? io_ins_178 : _GEN_177; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_179 = 9'hb3 == io_sel ? io_ins_179 : _GEN_178; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_180 = 9'hb4 == io_sel ? io_ins_180 : _GEN_179; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_181 = 9'hb5 == io_sel ? io_ins_181 : _GEN_180; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_182 = 9'hb6 == io_sel ? io_ins_182 : _GEN_181; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_183 = 9'hb7 == io_sel ? io_ins_183 : _GEN_182; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_184 = 9'hb8 == io_sel ? io_ins_184 : _GEN_183; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_185 = 9'hb9 == io_sel ? io_ins_185 : _GEN_184; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_186 = 9'hba == io_sel ? io_ins_186 : _GEN_185; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_187 = 9'hbb == io_sel ? io_ins_187 : _GEN_186; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_188 = 9'hbc == io_sel ? io_ins_188 : _GEN_187; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_189 = 9'hbd == io_sel ? io_ins_189 : _GEN_188; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_190 = 9'hbe == io_sel ? io_ins_190 : _GEN_189; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_191 = 9'hbf == io_sel ? io_ins_191 : _GEN_190; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_192 = 9'hc0 == io_sel ? io_ins_192 : _GEN_191; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_193 = 9'hc1 == io_sel ? io_ins_193 : _GEN_192; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_194 = 9'hc2 == io_sel ? io_ins_194 : _GEN_193; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_195 = 9'hc3 == io_sel ? io_ins_195 : _GEN_194; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_196 = 9'hc4 == io_sel ? io_ins_196 : _GEN_195; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_197 = 9'hc5 == io_sel ? io_ins_197 : _GEN_196; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_198 = 9'hc6 == io_sel ? io_ins_198 : _GEN_197; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_199 = 9'hc7 == io_sel ? io_ins_199 : _GEN_198; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_200 = 9'hc8 == io_sel ? io_ins_200 : _GEN_199; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_201 = 9'hc9 == io_sel ? io_ins_201 : _GEN_200; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_202 = 9'hca == io_sel ? io_ins_202 : _GEN_201; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_203 = 9'hcb == io_sel ? io_ins_203 : _GEN_202; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_204 = 9'hcc == io_sel ? io_ins_204 : _GEN_203; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_205 = 9'hcd == io_sel ? io_ins_205 : _GEN_204; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_206 = 9'hce == io_sel ? io_ins_206 : _GEN_205; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_207 = 9'hcf == io_sel ? io_ins_207 : _GEN_206; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_208 = 9'hd0 == io_sel ? io_ins_208 : _GEN_207; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_209 = 9'hd1 == io_sel ? io_ins_209 : _GEN_208; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_210 = 9'hd2 == io_sel ? io_ins_210 : _GEN_209; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_211 = 9'hd3 == io_sel ? io_ins_211 : _GEN_210; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_212 = 9'hd4 == io_sel ? io_ins_212 : _GEN_211; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_213 = 9'hd5 == io_sel ? io_ins_213 : _GEN_212; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_214 = 9'hd6 == io_sel ? io_ins_214 : _GEN_213; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_215 = 9'hd7 == io_sel ? io_ins_215 : _GEN_214; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_216 = 9'hd8 == io_sel ? io_ins_216 : _GEN_215; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_217 = 9'hd9 == io_sel ? io_ins_217 : _GEN_216; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_218 = 9'hda == io_sel ? io_ins_218 : _GEN_217; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_219 = 9'hdb == io_sel ? io_ins_219 : _GEN_218; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_220 = 9'hdc == io_sel ? io_ins_220 : _GEN_219; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_221 = 9'hdd == io_sel ? io_ins_221 : _GEN_220; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_222 = 9'hde == io_sel ? io_ins_222 : _GEN_221; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_223 = 9'hdf == io_sel ? io_ins_223 : _GEN_222; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_224 = 9'he0 == io_sel ? io_ins_224 : _GEN_223; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_225 = 9'he1 == io_sel ? io_ins_225 : _GEN_224; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_226 = 9'he2 == io_sel ? io_ins_226 : _GEN_225; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_227 = 9'he3 == io_sel ? io_ins_227 : _GEN_226; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_228 = 9'he4 == io_sel ? io_ins_228 : _GEN_227; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_229 = 9'he5 == io_sel ? io_ins_229 : _GEN_228; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_230 = 9'he6 == io_sel ? io_ins_230 : _GEN_229; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_231 = 9'he7 == io_sel ? io_ins_231 : _GEN_230; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_232 = 9'he8 == io_sel ? io_ins_232 : _GEN_231; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_233 = 9'he9 == io_sel ? io_ins_233 : _GEN_232; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_234 = 9'hea == io_sel ? io_ins_234 : _GEN_233; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_235 = 9'heb == io_sel ? io_ins_235 : _GEN_234; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_236 = 9'hec == io_sel ? io_ins_236 : _GEN_235; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_237 = 9'hed == io_sel ? io_ins_237 : _GEN_236; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_238 = 9'hee == io_sel ? io_ins_238 : _GEN_237; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_239 = 9'hef == io_sel ? io_ins_239 : _GEN_238; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_240 = 9'hf0 == io_sel ? io_ins_240 : _GEN_239; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_241 = 9'hf1 == io_sel ? io_ins_241 : _GEN_240; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_242 = 9'hf2 == io_sel ? io_ins_242 : _GEN_241; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_243 = 9'hf3 == io_sel ? io_ins_243 : _GEN_242; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_244 = 9'hf4 == io_sel ? io_ins_244 : _GEN_243; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_245 = 9'hf5 == io_sel ? io_ins_245 : _GEN_244; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_246 = 9'hf6 == io_sel ? io_ins_246 : _GEN_245; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_247 = 9'hf7 == io_sel ? io_ins_247 : _GEN_246; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_248 = 9'hf8 == io_sel ? io_ins_248 : _GEN_247; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_249 = 9'hf9 == io_sel ? io_ins_249 : _GEN_248; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_250 = 9'hfa == io_sel ? io_ins_250 : _GEN_249; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_251 = 9'hfb == io_sel ? io_ins_251 : _GEN_250; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_252 = 9'hfc == io_sel ? io_ins_252 : _GEN_251; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_253 = 9'hfd == io_sel ? io_ins_253 : _GEN_252; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_254 = 9'hfe == io_sel ? io_ins_254 : _GEN_253; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_255 = 9'hff == io_sel ? io_ins_255 : _GEN_254; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_256 = 9'h100 == io_sel ? io_ins_256 : _GEN_255; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_257 = 9'h101 == io_sel ? io_ins_257 : _GEN_256; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_258 = 9'h102 == io_sel ? io_ins_258 : _GEN_257; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_259 = 9'h103 == io_sel ? io_ins_259 : _GEN_258; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_260 = 9'h104 == io_sel ? io_ins_260 : _GEN_259; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_261 = 9'h105 == io_sel ? io_ins_261 : _GEN_260; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_262 = 9'h106 == io_sel ? io_ins_262 : _GEN_261; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_263 = 9'h107 == io_sel ? io_ins_263 : _GEN_262; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_264 = 9'h108 == io_sel ? io_ins_264 : _GEN_263; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_265 = 9'h109 == io_sel ? io_ins_265 : _GEN_264; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_266 = 9'h10a == io_sel ? io_ins_266 : _GEN_265; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_267 = 9'h10b == io_sel ? io_ins_267 : _GEN_266; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_268 = 9'h10c == io_sel ? io_ins_268 : _GEN_267; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_269 = 9'h10d == io_sel ? io_ins_269 : _GEN_268; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_270 = 9'h10e == io_sel ? io_ins_270 : _GEN_269; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_271 = 9'h10f == io_sel ? io_ins_271 : _GEN_270; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_272 = 9'h110 == io_sel ? io_ins_272 : _GEN_271; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_273 = 9'h111 == io_sel ? io_ins_273 : _GEN_272; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_274 = 9'h112 == io_sel ? io_ins_274 : _GEN_273; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_275 = 9'h113 == io_sel ? io_ins_275 : _GEN_274; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_276 = 9'h114 == io_sel ? io_ins_276 : _GEN_275; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_277 = 9'h115 == io_sel ? io_ins_277 : _GEN_276; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_278 = 9'h116 == io_sel ? io_ins_278 : _GEN_277; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_279 = 9'h117 == io_sel ? io_ins_279 : _GEN_278; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_280 = 9'h118 == io_sel ? io_ins_280 : _GEN_279; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_281 = 9'h119 == io_sel ? io_ins_281 : _GEN_280; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_282 = 9'h11a == io_sel ? io_ins_282 : _GEN_281; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_283 = 9'h11b == io_sel ? io_ins_283 : _GEN_282; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_284 = 9'h11c == io_sel ? io_ins_284 : _GEN_283; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_285 = 9'h11d == io_sel ? io_ins_285 : _GEN_284; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_286 = 9'h11e == io_sel ? io_ins_286 : _GEN_285; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_287 = 9'h11f == io_sel ? io_ins_287 : _GEN_286; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_288 = 9'h120 == io_sel ? io_ins_288 : _GEN_287; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_289 = 9'h121 == io_sel ? io_ins_289 : _GEN_288; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_290 = 9'h122 == io_sel ? io_ins_290 : _GEN_289; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_291 = 9'h123 == io_sel ? io_ins_291 : _GEN_290; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_292 = 9'h124 == io_sel ? io_ins_292 : _GEN_291; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_293 = 9'h125 == io_sel ? io_ins_293 : _GEN_292; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_294 = 9'h126 == io_sel ? io_ins_294 : _GEN_293; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_295 = 9'h127 == io_sel ? io_ins_295 : _GEN_294; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_296 = 9'h128 == io_sel ? io_ins_296 : _GEN_295; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_297 = 9'h129 == io_sel ? io_ins_297 : _GEN_296; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_298 = 9'h12a == io_sel ? io_ins_298 : _GEN_297; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_299 = 9'h12b == io_sel ? io_ins_299 : _GEN_298; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_300 = 9'h12c == io_sel ? io_ins_300 : _GEN_299; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_301 = 9'h12d == io_sel ? io_ins_301 : _GEN_300; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_302 = 9'h12e == io_sel ? io_ins_302 : _GEN_301; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_303 = 9'h12f == io_sel ? io_ins_303 : _GEN_302; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_304 = 9'h130 == io_sel ? io_ins_304 : _GEN_303; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_305 = 9'h131 == io_sel ? io_ins_305 : _GEN_304; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_306 = 9'h132 == io_sel ? io_ins_306 : _GEN_305; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_307 = 9'h133 == io_sel ? io_ins_307 : _GEN_306; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_308 = 9'h134 == io_sel ? io_ins_308 : _GEN_307; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_309 = 9'h135 == io_sel ? io_ins_309 : _GEN_308; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_310 = 9'h136 == io_sel ? io_ins_310 : _GEN_309; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_311 = 9'h137 == io_sel ? io_ins_311 : _GEN_310; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_312 = 9'h138 == io_sel ? io_ins_312 : _GEN_311; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_313 = 9'h139 == io_sel ? io_ins_313 : _GEN_312; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_314 = 9'h13a == io_sel ? io_ins_314 : _GEN_313; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_315 = 9'h13b == io_sel ? io_ins_315 : _GEN_314; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_316 = 9'h13c == io_sel ? io_ins_316 : _GEN_315; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_317 = 9'h13d == io_sel ? io_ins_317 : _GEN_316; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_318 = 9'h13e == io_sel ? io_ins_318 : _GEN_317; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_319 = 9'h13f == io_sel ? io_ins_319 : _GEN_318; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_320 = 9'h140 == io_sel ? io_ins_320 : _GEN_319; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_321 = 9'h141 == io_sel ? io_ins_321 : _GEN_320; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_322 = 9'h142 == io_sel ? io_ins_322 : _GEN_321; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_323 = 9'h143 == io_sel ? io_ins_323 : _GEN_322; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_324 = 9'h144 == io_sel ? io_ins_324 : _GEN_323; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_325 = 9'h145 == io_sel ? io_ins_325 : _GEN_324; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_326 = 9'h146 == io_sel ? io_ins_326 : _GEN_325; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_327 = 9'h147 == io_sel ? io_ins_327 : _GEN_326; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_328 = 9'h148 == io_sel ? io_ins_328 : _GEN_327; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_329 = 9'h149 == io_sel ? io_ins_329 : _GEN_328; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_330 = 9'h14a == io_sel ? io_ins_330 : _GEN_329; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_331 = 9'h14b == io_sel ? io_ins_331 : _GEN_330; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_332 = 9'h14c == io_sel ? io_ins_332 : _GEN_331; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_333 = 9'h14d == io_sel ? io_ins_333 : _GEN_332; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_334 = 9'h14e == io_sel ? io_ins_334 : _GEN_333; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_335 = 9'h14f == io_sel ? io_ins_335 : _GEN_334; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_336 = 9'h150 == io_sel ? io_ins_336 : _GEN_335; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_337 = 9'h151 == io_sel ? io_ins_337 : _GEN_336; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_338 = 9'h152 == io_sel ? io_ins_338 : _GEN_337; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_339 = 9'h153 == io_sel ? io_ins_339 : _GEN_338; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_340 = 9'h154 == io_sel ? io_ins_340 : _GEN_339; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_341 = 9'h155 == io_sel ? io_ins_341 : _GEN_340; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_342 = 9'h156 == io_sel ? io_ins_342 : _GEN_341; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_343 = 9'h157 == io_sel ? io_ins_343 : _GEN_342; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_344 = 9'h158 == io_sel ? io_ins_344 : _GEN_343; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_345 = 9'h159 == io_sel ? io_ins_345 : _GEN_344; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_346 = 9'h15a == io_sel ? io_ins_346 : _GEN_345; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_347 = 9'h15b == io_sel ? io_ins_347 : _GEN_346; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_348 = 9'h15c == io_sel ? io_ins_348 : _GEN_347; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_349 = 9'h15d == io_sel ? io_ins_349 : _GEN_348; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_350 = 9'h15e == io_sel ? io_ins_350 : _GEN_349; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_351 = 9'h15f == io_sel ? io_ins_351 : _GEN_350; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_352 = 9'h160 == io_sel ? io_ins_352 : _GEN_351; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_353 = 9'h161 == io_sel ? io_ins_353 : _GEN_352; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_354 = 9'h162 == io_sel ? io_ins_354 : _GEN_353; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_355 = 9'h163 == io_sel ? io_ins_355 : _GEN_354; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_356 = 9'h164 == io_sel ? io_ins_356 : _GEN_355; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_357 = 9'h165 == io_sel ? io_ins_357 : _GEN_356; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_358 = 9'h166 == io_sel ? io_ins_358 : _GEN_357; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_359 = 9'h167 == io_sel ? io_ins_359 : _GEN_358; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_360 = 9'h168 == io_sel ? io_ins_360 : _GEN_359; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_361 = 9'h169 == io_sel ? io_ins_361 : _GEN_360; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_362 = 9'h16a == io_sel ? io_ins_362 : _GEN_361; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_363 = 9'h16b == io_sel ? io_ins_363 : _GEN_362; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_364 = 9'h16c == io_sel ? io_ins_364 : _GEN_363; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_365 = 9'h16d == io_sel ? io_ins_365 : _GEN_364; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_366 = 9'h16e == io_sel ? io_ins_366 : _GEN_365; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_367 = 9'h16f == io_sel ? io_ins_367 : _GEN_366; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_368 = 9'h170 == io_sel ? io_ins_368 : _GEN_367; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_369 = 9'h171 == io_sel ? io_ins_369 : _GEN_368; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_370 = 9'h172 == io_sel ? io_ins_370 : _GEN_369; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_371 = 9'h173 == io_sel ? io_ins_371 : _GEN_370; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_372 = 9'h174 == io_sel ? io_ins_372 : _GEN_371; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_373 = 9'h175 == io_sel ? io_ins_373 : _GEN_372; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_374 = 9'h176 == io_sel ? io_ins_374 : _GEN_373; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_375 = 9'h177 == io_sel ? io_ins_375 : _GEN_374; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_376 = 9'h178 == io_sel ? io_ins_376 : _GEN_375; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_377 = 9'h179 == io_sel ? io_ins_377 : _GEN_376; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_378 = 9'h17a == io_sel ? io_ins_378 : _GEN_377; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_379 = 9'h17b == io_sel ? io_ins_379 : _GEN_378; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_380 = 9'h17c == io_sel ? io_ins_380 : _GEN_379; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_381 = 9'h17d == io_sel ? io_ins_381 : _GEN_380; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_382 = 9'h17e == io_sel ? io_ins_382 : _GEN_381; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_383 = 9'h17f == io_sel ? io_ins_383 : _GEN_382; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_384 = 9'h180 == io_sel ? io_ins_384 : _GEN_383; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_385 = 9'h181 == io_sel ? io_ins_385 : _GEN_384; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_386 = 9'h182 == io_sel ? io_ins_386 : _GEN_385; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_387 = 9'h183 == io_sel ? io_ins_387 : _GEN_386; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_388 = 9'h184 == io_sel ? io_ins_388 : _GEN_387; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_389 = 9'h185 == io_sel ? io_ins_389 : _GEN_388; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_390 = 9'h186 == io_sel ? io_ins_390 : _GEN_389; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_391 = 9'h187 == io_sel ? io_ins_391 : _GEN_390; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_392 = 9'h188 == io_sel ? io_ins_392 : _GEN_391; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_393 = 9'h189 == io_sel ? io_ins_393 : _GEN_392; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_394 = 9'h18a == io_sel ? io_ins_394 : _GEN_393; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_395 = 9'h18b == io_sel ? io_ins_395 : _GEN_394; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_396 = 9'h18c == io_sel ? io_ins_396 : _GEN_395; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_397 = 9'h18d == io_sel ? io_ins_397 : _GEN_396; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_398 = 9'h18e == io_sel ? io_ins_398 : _GEN_397; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_399 = 9'h18f == io_sel ? io_ins_399 : _GEN_398; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_400 = 9'h190 == io_sel ? io_ins_400 : _GEN_399; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_401 = 9'h191 == io_sel ? io_ins_401 : _GEN_400; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_402 = 9'h192 == io_sel ? io_ins_402 : _GEN_401; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_403 = 9'h193 == io_sel ? io_ins_403 : _GEN_402; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_404 = 9'h194 == io_sel ? io_ins_404 : _GEN_403; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_405 = 9'h195 == io_sel ? io_ins_405 : _GEN_404; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_406 = 9'h196 == io_sel ? io_ins_406 : _GEN_405; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_407 = 9'h197 == io_sel ? io_ins_407 : _GEN_406; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_408 = 9'h198 == io_sel ? io_ins_408 : _GEN_407; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_409 = 9'h199 == io_sel ? io_ins_409 : _GEN_408; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_410 = 9'h19a == io_sel ? io_ins_410 : _GEN_409; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_411 = 9'h19b == io_sel ? io_ins_411 : _GEN_410; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_412 = 9'h19c == io_sel ? io_ins_412 : _GEN_411; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_413 = 9'h19d == io_sel ? io_ins_413 : _GEN_412; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_414 = 9'h19e == io_sel ? io_ins_414 : _GEN_413; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_415 = 9'h19f == io_sel ? io_ins_415 : _GEN_414; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_416 = 9'h1a0 == io_sel ? io_ins_416 : _GEN_415; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_417 = 9'h1a1 == io_sel ? io_ins_417 : _GEN_416; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_418 = 9'h1a2 == io_sel ? io_ins_418 : _GEN_417; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_419 = 9'h1a3 == io_sel ? io_ins_419 : _GEN_418; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_420 = 9'h1a4 == io_sel ? io_ins_420 : _GEN_419; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_421 = 9'h1a5 == io_sel ? io_ins_421 : _GEN_420; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_422 = 9'h1a6 == io_sel ? io_ins_422 : _GEN_421; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_423 = 9'h1a7 == io_sel ? io_ins_423 : _GEN_422; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_424 = 9'h1a8 == io_sel ? io_ins_424 : _GEN_423; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_425 = 9'h1a9 == io_sel ? io_ins_425 : _GEN_424; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_426 = 9'h1aa == io_sel ? io_ins_426 : _GEN_425; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_427 = 9'h1ab == io_sel ? io_ins_427 : _GEN_426; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_428 = 9'h1ac == io_sel ? io_ins_428 : _GEN_427; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_429 = 9'h1ad == io_sel ? io_ins_429 : _GEN_428; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_430 = 9'h1ae == io_sel ? io_ins_430 : _GEN_429; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_431 = 9'h1af == io_sel ? io_ins_431 : _GEN_430; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_432 = 9'h1b0 == io_sel ? io_ins_432 : _GEN_431; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_433 = 9'h1b1 == io_sel ? io_ins_433 : _GEN_432; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_434 = 9'h1b2 == io_sel ? io_ins_434 : _GEN_433; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_435 = 9'h1b3 == io_sel ? io_ins_435 : _GEN_434; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_436 = 9'h1b4 == io_sel ? io_ins_436 : _GEN_435; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_437 = 9'h1b5 == io_sel ? io_ins_437 : _GEN_436; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_438 = 9'h1b6 == io_sel ? io_ins_438 : _GEN_437; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_439 = 9'h1b7 == io_sel ? io_ins_439 : _GEN_438; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_440 = 9'h1b8 == io_sel ? io_ins_440 : _GEN_439; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_441 = 9'h1b9 == io_sel ? io_ins_441 : _GEN_440; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_442 = 9'h1ba == io_sel ? io_ins_442 : _GEN_441; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_443 = 9'h1bb == io_sel ? io_ins_443 : _GEN_442; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_444 = 9'h1bc == io_sel ? io_ins_444 : _GEN_443; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_445 = 9'h1bd == io_sel ? io_ins_445 : _GEN_444; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_446 = 9'h1be == io_sel ? io_ins_446 : _GEN_445; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_447 = 9'h1bf == io_sel ? io_ins_447 : _GEN_446; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_448 = 9'h1c0 == io_sel ? io_ins_448 : _GEN_447; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_449 = 9'h1c1 == io_sel ? io_ins_449 : _GEN_448; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_450 = 9'h1c2 == io_sel ? io_ins_450 : _GEN_449; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_451 = 9'h1c3 == io_sel ? io_ins_451 : _GEN_450; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_452 = 9'h1c4 == io_sel ? io_ins_452 : _GEN_451; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_453 = 9'h1c5 == io_sel ? io_ins_453 : _GEN_452; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_454 = 9'h1c6 == io_sel ? io_ins_454 : _GEN_453; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_455 = 9'h1c7 == io_sel ? io_ins_455 : _GEN_454; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_456 = 9'h1c8 == io_sel ? io_ins_456 : _GEN_455; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_457 = 9'h1c9 == io_sel ? io_ins_457 : _GEN_456; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_458 = 9'h1ca == io_sel ? io_ins_458 : _GEN_457; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_459 = 9'h1cb == io_sel ? io_ins_459 : _GEN_458; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_460 = 9'h1cc == io_sel ? io_ins_460 : _GEN_459; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_461 = 9'h1cd == io_sel ? io_ins_461 : _GEN_460; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_462 = 9'h1ce == io_sel ? io_ins_462 : _GEN_461; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_463 = 9'h1cf == io_sel ? io_ins_463 : _GEN_462; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_464 = 9'h1d0 == io_sel ? io_ins_464 : _GEN_463; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_465 = 9'h1d1 == io_sel ? io_ins_465 : _GEN_464; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_466 = 9'h1d2 == io_sel ? io_ins_466 : _GEN_465; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_467 = 9'h1d3 == io_sel ? io_ins_467 : _GEN_466; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_468 = 9'h1d4 == io_sel ? io_ins_468 : _GEN_467; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_469 = 9'h1d5 == io_sel ? io_ins_469 : _GEN_468; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_470 = 9'h1d6 == io_sel ? io_ins_470 : _GEN_469; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_471 = 9'h1d7 == io_sel ? io_ins_471 : _GEN_470; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_472 = 9'h1d8 == io_sel ? io_ins_472 : _GEN_471; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_473 = 9'h1d9 == io_sel ? io_ins_473 : _GEN_472; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_474 = 9'h1da == io_sel ? io_ins_474 : _GEN_473; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_475 = 9'h1db == io_sel ? io_ins_475 : _GEN_474; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_476 = 9'h1dc == io_sel ? io_ins_476 : _GEN_475; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_477 = 9'h1dd == io_sel ? io_ins_477 : _GEN_476; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_478 = 9'h1de == io_sel ? io_ins_478 : _GEN_477; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_479 = 9'h1df == io_sel ? io_ins_479 : _GEN_478; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_480 = 9'h1e0 == io_sel ? io_ins_480 : _GEN_479; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_481 = 9'h1e1 == io_sel ? io_ins_481 : _GEN_480; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_482 = 9'h1e2 == io_sel ? io_ins_482 : _GEN_481; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_483 = 9'h1e3 == io_sel ? io_ins_483 : _GEN_482; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_484 = 9'h1e4 == io_sel ? io_ins_484 : _GEN_483; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_485 = 9'h1e5 == io_sel ? io_ins_485 : _GEN_484; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_486 = 9'h1e6 == io_sel ? io_ins_486 : _GEN_485; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_487 = 9'h1e7 == io_sel ? io_ins_487 : _GEN_486; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_488 = 9'h1e8 == io_sel ? io_ins_488 : _GEN_487; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_489 = 9'h1e9 == io_sel ? io_ins_489 : _GEN_488; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_490 = 9'h1ea == io_sel ? io_ins_490 : _GEN_489; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_491 = 9'h1eb == io_sel ? io_ins_491 : _GEN_490; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_492 = 9'h1ec == io_sel ? io_ins_492 : _GEN_491; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_493 = 9'h1ed == io_sel ? io_ins_493 : _GEN_492; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_494 = 9'h1ee == io_sel ? io_ins_494 : _GEN_493; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_495 = 9'h1ef == io_sel ? io_ins_495 : _GEN_494; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_496 = 9'h1f0 == io_sel ? io_ins_496 : _GEN_495; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_497 = 9'h1f1 == io_sel ? io_ins_497 : _GEN_496; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_498 = 9'h1f2 == io_sel ? io_ins_498 : _GEN_497; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_499 = 9'h1f3 == io_sel ? io_ins_499 : _GEN_498; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_500 = 9'h1f4 == io_sel ? io_ins_500 : _GEN_499; // @[MuxN.scala 16:10:@32240.4]
  assign _GEN_501 = 9'h1f5 == io_sel ? io_ins_501 : _GEN_500; // @[MuxN.scala 16:10:@32240.4]
  assign io_out = 9'h1f6 == io_sel ? io_ins_502 : _GEN_501; // @[MuxN.scala 16:10:@32240.4]
endmodule
module RegFile( // @[:@32242.2]
  input         clock, // @[:@32243.4]
  input         reset, // @[:@32244.4]
  input  [31:0] io_raddr, // @[:@32245.4]
  input         io_wen, // @[:@32245.4]
  input  [31:0] io_waddr, // @[:@32245.4]
  input  [63:0] io_wdata, // @[:@32245.4]
  output [63:0] io_rdata, // @[:@32245.4]
  input         io_reset, // @[:@32245.4]
  output [63:0] io_argIns_0, // @[:@32245.4]
  output [63:0] io_argIns_1, // @[:@32245.4]
  output [63:0] io_argIns_2, // @[:@32245.4]
  input         io_argOuts_0_valid, // @[:@32245.4]
  input  [63:0] io_argOuts_0_bits, // @[:@32245.4]
  input         io_argOuts_1_valid, // @[:@32245.4]
  input  [63:0] io_argOuts_1_bits // @[:@32245.4]
);
  wire  regs_0_clock; // @[RegFile.scala 66:20:@34255.4]
  wire  regs_0_reset; // @[RegFile.scala 66:20:@34255.4]
  wire [63:0] regs_0_io_in; // @[RegFile.scala 66:20:@34255.4]
  wire  regs_0_io_reset; // @[RegFile.scala 66:20:@34255.4]
  wire [63:0] regs_0_io_out; // @[RegFile.scala 66:20:@34255.4]
  wire  regs_0_io_enable; // @[RegFile.scala 66:20:@34255.4]
  wire  regs_1_clock; // @[RegFile.scala 66:20:@34267.4]
  wire  regs_1_reset; // @[RegFile.scala 66:20:@34267.4]
  wire [63:0] regs_1_io_in; // @[RegFile.scala 66:20:@34267.4]
  wire  regs_1_io_reset; // @[RegFile.scala 66:20:@34267.4]
  wire [63:0] regs_1_io_out; // @[RegFile.scala 66:20:@34267.4]
  wire  regs_1_io_enable; // @[RegFile.scala 66:20:@34267.4]
  wire  regs_2_clock; // @[RegFile.scala 66:20:@34286.4]
  wire  regs_2_reset; // @[RegFile.scala 66:20:@34286.4]
  wire [63:0] regs_2_io_in; // @[RegFile.scala 66:20:@34286.4]
  wire  regs_2_io_reset; // @[RegFile.scala 66:20:@34286.4]
  wire [63:0] regs_2_io_out; // @[RegFile.scala 66:20:@34286.4]
  wire  regs_2_io_enable; // @[RegFile.scala 66:20:@34286.4]
  wire  regs_3_clock; // @[RegFile.scala 66:20:@34298.4]
  wire  regs_3_reset; // @[RegFile.scala 66:20:@34298.4]
  wire [63:0] regs_3_io_in; // @[RegFile.scala 66:20:@34298.4]
  wire  regs_3_io_reset; // @[RegFile.scala 66:20:@34298.4]
  wire [63:0] regs_3_io_out; // @[RegFile.scala 66:20:@34298.4]
  wire  regs_3_io_enable; // @[RegFile.scala 66:20:@34298.4]
  wire  regs_4_clock; // @[RegFile.scala 66:20:@34312.4]
  wire  regs_4_reset; // @[RegFile.scala 66:20:@34312.4]
  wire [63:0] regs_4_io_in; // @[RegFile.scala 66:20:@34312.4]
  wire  regs_4_io_reset; // @[RegFile.scala 66:20:@34312.4]
  wire [63:0] regs_4_io_out; // @[RegFile.scala 66:20:@34312.4]
  wire  regs_4_io_enable; // @[RegFile.scala 66:20:@34312.4]
  wire  regs_5_clock; // @[RegFile.scala 66:20:@34326.4]
  wire  regs_5_reset; // @[RegFile.scala 66:20:@34326.4]
  wire [63:0] regs_5_io_in; // @[RegFile.scala 66:20:@34326.4]
  wire  regs_5_io_reset; // @[RegFile.scala 66:20:@34326.4]
  wire [63:0] regs_5_io_out; // @[RegFile.scala 66:20:@34326.4]
  wire  regs_5_io_enable; // @[RegFile.scala 66:20:@34326.4]
  wire  regs_6_clock; // @[RegFile.scala 66:20:@34340.4]
  wire  regs_6_reset; // @[RegFile.scala 66:20:@34340.4]
  wire [63:0] regs_6_io_in; // @[RegFile.scala 66:20:@34340.4]
  wire  regs_6_io_reset; // @[RegFile.scala 66:20:@34340.4]
  wire [63:0] regs_6_io_out; // @[RegFile.scala 66:20:@34340.4]
  wire  regs_6_io_enable; // @[RegFile.scala 66:20:@34340.4]
  wire  regs_7_clock; // @[RegFile.scala 66:20:@34354.4]
  wire  regs_7_reset; // @[RegFile.scala 66:20:@34354.4]
  wire [63:0] regs_7_io_in; // @[RegFile.scala 66:20:@34354.4]
  wire  regs_7_io_reset; // @[RegFile.scala 66:20:@34354.4]
  wire [63:0] regs_7_io_out; // @[RegFile.scala 66:20:@34354.4]
  wire  regs_7_io_enable; // @[RegFile.scala 66:20:@34354.4]
  wire  regs_8_clock; // @[RegFile.scala 66:20:@34368.4]
  wire  regs_8_reset; // @[RegFile.scala 66:20:@34368.4]
  wire [63:0] regs_8_io_in; // @[RegFile.scala 66:20:@34368.4]
  wire  regs_8_io_reset; // @[RegFile.scala 66:20:@34368.4]
  wire [63:0] regs_8_io_out; // @[RegFile.scala 66:20:@34368.4]
  wire  regs_8_io_enable; // @[RegFile.scala 66:20:@34368.4]
  wire  regs_9_clock; // @[RegFile.scala 66:20:@34382.4]
  wire  regs_9_reset; // @[RegFile.scala 66:20:@34382.4]
  wire [63:0] regs_9_io_in; // @[RegFile.scala 66:20:@34382.4]
  wire  regs_9_io_reset; // @[RegFile.scala 66:20:@34382.4]
  wire [63:0] regs_9_io_out; // @[RegFile.scala 66:20:@34382.4]
  wire  regs_9_io_enable; // @[RegFile.scala 66:20:@34382.4]
  wire  regs_10_clock; // @[RegFile.scala 66:20:@34396.4]
  wire  regs_10_reset; // @[RegFile.scala 66:20:@34396.4]
  wire [63:0] regs_10_io_in; // @[RegFile.scala 66:20:@34396.4]
  wire  regs_10_io_reset; // @[RegFile.scala 66:20:@34396.4]
  wire [63:0] regs_10_io_out; // @[RegFile.scala 66:20:@34396.4]
  wire  regs_10_io_enable; // @[RegFile.scala 66:20:@34396.4]
  wire  regs_11_clock; // @[RegFile.scala 66:20:@34410.4]
  wire  regs_11_reset; // @[RegFile.scala 66:20:@34410.4]
  wire [63:0] regs_11_io_in; // @[RegFile.scala 66:20:@34410.4]
  wire  regs_11_io_reset; // @[RegFile.scala 66:20:@34410.4]
  wire [63:0] regs_11_io_out; // @[RegFile.scala 66:20:@34410.4]
  wire  regs_11_io_enable; // @[RegFile.scala 66:20:@34410.4]
  wire  regs_12_clock; // @[RegFile.scala 66:20:@34424.4]
  wire  regs_12_reset; // @[RegFile.scala 66:20:@34424.4]
  wire [63:0] regs_12_io_in; // @[RegFile.scala 66:20:@34424.4]
  wire  regs_12_io_reset; // @[RegFile.scala 66:20:@34424.4]
  wire [63:0] regs_12_io_out; // @[RegFile.scala 66:20:@34424.4]
  wire  regs_12_io_enable; // @[RegFile.scala 66:20:@34424.4]
  wire  regs_13_clock; // @[RegFile.scala 66:20:@34438.4]
  wire  regs_13_reset; // @[RegFile.scala 66:20:@34438.4]
  wire [63:0] regs_13_io_in; // @[RegFile.scala 66:20:@34438.4]
  wire  regs_13_io_reset; // @[RegFile.scala 66:20:@34438.4]
  wire [63:0] regs_13_io_out; // @[RegFile.scala 66:20:@34438.4]
  wire  regs_13_io_enable; // @[RegFile.scala 66:20:@34438.4]
  wire  regs_14_clock; // @[RegFile.scala 66:20:@34452.4]
  wire  regs_14_reset; // @[RegFile.scala 66:20:@34452.4]
  wire [63:0] regs_14_io_in; // @[RegFile.scala 66:20:@34452.4]
  wire  regs_14_io_reset; // @[RegFile.scala 66:20:@34452.4]
  wire [63:0] regs_14_io_out; // @[RegFile.scala 66:20:@34452.4]
  wire  regs_14_io_enable; // @[RegFile.scala 66:20:@34452.4]
  wire  regs_15_clock; // @[RegFile.scala 66:20:@34466.4]
  wire  regs_15_reset; // @[RegFile.scala 66:20:@34466.4]
  wire [63:0] regs_15_io_in; // @[RegFile.scala 66:20:@34466.4]
  wire  regs_15_io_reset; // @[RegFile.scala 66:20:@34466.4]
  wire [63:0] regs_15_io_out; // @[RegFile.scala 66:20:@34466.4]
  wire  regs_15_io_enable; // @[RegFile.scala 66:20:@34466.4]
  wire  regs_16_clock; // @[RegFile.scala 66:20:@34480.4]
  wire  regs_16_reset; // @[RegFile.scala 66:20:@34480.4]
  wire [63:0] regs_16_io_in; // @[RegFile.scala 66:20:@34480.4]
  wire  regs_16_io_reset; // @[RegFile.scala 66:20:@34480.4]
  wire [63:0] regs_16_io_out; // @[RegFile.scala 66:20:@34480.4]
  wire  regs_16_io_enable; // @[RegFile.scala 66:20:@34480.4]
  wire  regs_17_clock; // @[RegFile.scala 66:20:@34494.4]
  wire  regs_17_reset; // @[RegFile.scala 66:20:@34494.4]
  wire [63:0] regs_17_io_in; // @[RegFile.scala 66:20:@34494.4]
  wire  regs_17_io_reset; // @[RegFile.scala 66:20:@34494.4]
  wire [63:0] regs_17_io_out; // @[RegFile.scala 66:20:@34494.4]
  wire  regs_17_io_enable; // @[RegFile.scala 66:20:@34494.4]
  wire  regs_18_clock; // @[RegFile.scala 66:20:@34508.4]
  wire  regs_18_reset; // @[RegFile.scala 66:20:@34508.4]
  wire [63:0] regs_18_io_in; // @[RegFile.scala 66:20:@34508.4]
  wire  regs_18_io_reset; // @[RegFile.scala 66:20:@34508.4]
  wire [63:0] regs_18_io_out; // @[RegFile.scala 66:20:@34508.4]
  wire  regs_18_io_enable; // @[RegFile.scala 66:20:@34508.4]
  wire  regs_19_clock; // @[RegFile.scala 66:20:@34522.4]
  wire  regs_19_reset; // @[RegFile.scala 66:20:@34522.4]
  wire [63:0] regs_19_io_in; // @[RegFile.scala 66:20:@34522.4]
  wire  regs_19_io_reset; // @[RegFile.scala 66:20:@34522.4]
  wire [63:0] regs_19_io_out; // @[RegFile.scala 66:20:@34522.4]
  wire  regs_19_io_enable; // @[RegFile.scala 66:20:@34522.4]
  wire  regs_20_clock; // @[RegFile.scala 66:20:@34536.4]
  wire  regs_20_reset; // @[RegFile.scala 66:20:@34536.4]
  wire [63:0] regs_20_io_in; // @[RegFile.scala 66:20:@34536.4]
  wire  regs_20_io_reset; // @[RegFile.scala 66:20:@34536.4]
  wire [63:0] regs_20_io_out; // @[RegFile.scala 66:20:@34536.4]
  wire  regs_20_io_enable; // @[RegFile.scala 66:20:@34536.4]
  wire  regs_21_clock; // @[RegFile.scala 66:20:@34550.4]
  wire  regs_21_reset; // @[RegFile.scala 66:20:@34550.4]
  wire [63:0] regs_21_io_in; // @[RegFile.scala 66:20:@34550.4]
  wire  regs_21_io_reset; // @[RegFile.scala 66:20:@34550.4]
  wire [63:0] regs_21_io_out; // @[RegFile.scala 66:20:@34550.4]
  wire  regs_21_io_enable; // @[RegFile.scala 66:20:@34550.4]
  wire  regs_22_clock; // @[RegFile.scala 66:20:@34564.4]
  wire  regs_22_reset; // @[RegFile.scala 66:20:@34564.4]
  wire [63:0] regs_22_io_in; // @[RegFile.scala 66:20:@34564.4]
  wire  regs_22_io_reset; // @[RegFile.scala 66:20:@34564.4]
  wire [63:0] regs_22_io_out; // @[RegFile.scala 66:20:@34564.4]
  wire  regs_22_io_enable; // @[RegFile.scala 66:20:@34564.4]
  wire  regs_23_clock; // @[RegFile.scala 66:20:@34578.4]
  wire  regs_23_reset; // @[RegFile.scala 66:20:@34578.4]
  wire [63:0] regs_23_io_in; // @[RegFile.scala 66:20:@34578.4]
  wire  regs_23_io_reset; // @[RegFile.scala 66:20:@34578.4]
  wire [63:0] regs_23_io_out; // @[RegFile.scala 66:20:@34578.4]
  wire  regs_23_io_enable; // @[RegFile.scala 66:20:@34578.4]
  wire  regs_24_clock; // @[RegFile.scala 66:20:@34592.4]
  wire  regs_24_reset; // @[RegFile.scala 66:20:@34592.4]
  wire [63:0] regs_24_io_in; // @[RegFile.scala 66:20:@34592.4]
  wire  regs_24_io_reset; // @[RegFile.scala 66:20:@34592.4]
  wire [63:0] regs_24_io_out; // @[RegFile.scala 66:20:@34592.4]
  wire  regs_24_io_enable; // @[RegFile.scala 66:20:@34592.4]
  wire  regs_25_clock; // @[RegFile.scala 66:20:@34606.4]
  wire  regs_25_reset; // @[RegFile.scala 66:20:@34606.4]
  wire [63:0] regs_25_io_in; // @[RegFile.scala 66:20:@34606.4]
  wire  regs_25_io_reset; // @[RegFile.scala 66:20:@34606.4]
  wire [63:0] regs_25_io_out; // @[RegFile.scala 66:20:@34606.4]
  wire  regs_25_io_enable; // @[RegFile.scala 66:20:@34606.4]
  wire  regs_26_clock; // @[RegFile.scala 66:20:@34620.4]
  wire  regs_26_reset; // @[RegFile.scala 66:20:@34620.4]
  wire [63:0] regs_26_io_in; // @[RegFile.scala 66:20:@34620.4]
  wire  regs_26_io_reset; // @[RegFile.scala 66:20:@34620.4]
  wire [63:0] regs_26_io_out; // @[RegFile.scala 66:20:@34620.4]
  wire  regs_26_io_enable; // @[RegFile.scala 66:20:@34620.4]
  wire  regs_27_clock; // @[RegFile.scala 66:20:@34634.4]
  wire  regs_27_reset; // @[RegFile.scala 66:20:@34634.4]
  wire [63:0] regs_27_io_in; // @[RegFile.scala 66:20:@34634.4]
  wire  regs_27_io_reset; // @[RegFile.scala 66:20:@34634.4]
  wire [63:0] regs_27_io_out; // @[RegFile.scala 66:20:@34634.4]
  wire  regs_27_io_enable; // @[RegFile.scala 66:20:@34634.4]
  wire  regs_28_clock; // @[RegFile.scala 66:20:@34648.4]
  wire  regs_28_reset; // @[RegFile.scala 66:20:@34648.4]
  wire [63:0] regs_28_io_in; // @[RegFile.scala 66:20:@34648.4]
  wire  regs_28_io_reset; // @[RegFile.scala 66:20:@34648.4]
  wire [63:0] regs_28_io_out; // @[RegFile.scala 66:20:@34648.4]
  wire  regs_28_io_enable; // @[RegFile.scala 66:20:@34648.4]
  wire  regs_29_clock; // @[RegFile.scala 66:20:@34662.4]
  wire  regs_29_reset; // @[RegFile.scala 66:20:@34662.4]
  wire [63:0] regs_29_io_in; // @[RegFile.scala 66:20:@34662.4]
  wire  regs_29_io_reset; // @[RegFile.scala 66:20:@34662.4]
  wire [63:0] regs_29_io_out; // @[RegFile.scala 66:20:@34662.4]
  wire  regs_29_io_enable; // @[RegFile.scala 66:20:@34662.4]
  wire  regs_30_clock; // @[RegFile.scala 66:20:@34676.4]
  wire  regs_30_reset; // @[RegFile.scala 66:20:@34676.4]
  wire [63:0] regs_30_io_in; // @[RegFile.scala 66:20:@34676.4]
  wire  regs_30_io_reset; // @[RegFile.scala 66:20:@34676.4]
  wire [63:0] regs_30_io_out; // @[RegFile.scala 66:20:@34676.4]
  wire  regs_30_io_enable; // @[RegFile.scala 66:20:@34676.4]
  wire  regs_31_clock; // @[RegFile.scala 66:20:@34690.4]
  wire  regs_31_reset; // @[RegFile.scala 66:20:@34690.4]
  wire [63:0] regs_31_io_in; // @[RegFile.scala 66:20:@34690.4]
  wire  regs_31_io_reset; // @[RegFile.scala 66:20:@34690.4]
  wire [63:0] regs_31_io_out; // @[RegFile.scala 66:20:@34690.4]
  wire  regs_31_io_enable; // @[RegFile.scala 66:20:@34690.4]
  wire  regs_32_clock; // @[RegFile.scala 66:20:@34704.4]
  wire  regs_32_reset; // @[RegFile.scala 66:20:@34704.4]
  wire [63:0] regs_32_io_in; // @[RegFile.scala 66:20:@34704.4]
  wire  regs_32_io_reset; // @[RegFile.scala 66:20:@34704.4]
  wire [63:0] regs_32_io_out; // @[RegFile.scala 66:20:@34704.4]
  wire  regs_32_io_enable; // @[RegFile.scala 66:20:@34704.4]
  wire  regs_33_clock; // @[RegFile.scala 66:20:@34718.4]
  wire  regs_33_reset; // @[RegFile.scala 66:20:@34718.4]
  wire [63:0] regs_33_io_in; // @[RegFile.scala 66:20:@34718.4]
  wire  regs_33_io_reset; // @[RegFile.scala 66:20:@34718.4]
  wire [63:0] regs_33_io_out; // @[RegFile.scala 66:20:@34718.4]
  wire  regs_33_io_enable; // @[RegFile.scala 66:20:@34718.4]
  wire  regs_34_clock; // @[RegFile.scala 66:20:@34732.4]
  wire  regs_34_reset; // @[RegFile.scala 66:20:@34732.4]
  wire [63:0] regs_34_io_in; // @[RegFile.scala 66:20:@34732.4]
  wire  regs_34_io_reset; // @[RegFile.scala 66:20:@34732.4]
  wire [63:0] regs_34_io_out; // @[RegFile.scala 66:20:@34732.4]
  wire  regs_34_io_enable; // @[RegFile.scala 66:20:@34732.4]
  wire  regs_35_clock; // @[RegFile.scala 66:20:@34746.4]
  wire  regs_35_reset; // @[RegFile.scala 66:20:@34746.4]
  wire [63:0] regs_35_io_in; // @[RegFile.scala 66:20:@34746.4]
  wire  regs_35_io_reset; // @[RegFile.scala 66:20:@34746.4]
  wire [63:0] regs_35_io_out; // @[RegFile.scala 66:20:@34746.4]
  wire  regs_35_io_enable; // @[RegFile.scala 66:20:@34746.4]
  wire  regs_36_clock; // @[RegFile.scala 66:20:@34760.4]
  wire  regs_36_reset; // @[RegFile.scala 66:20:@34760.4]
  wire [63:0] regs_36_io_in; // @[RegFile.scala 66:20:@34760.4]
  wire  regs_36_io_reset; // @[RegFile.scala 66:20:@34760.4]
  wire [63:0] regs_36_io_out; // @[RegFile.scala 66:20:@34760.4]
  wire  regs_36_io_enable; // @[RegFile.scala 66:20:@34760.4]
  wire  regs_37_clock; // @[RegFile.scala 66:20:@34774.4]
  wire  regs_37_reset; // @[RegFile.scala 66:20:@34774.4]
  wire [63:0] regs_37_io_in; // @[RegFile.scala 66:20:@34774.4]
  wire  regs_37_io_reset; // @[RegFile.scala 66:20:@34774.4]
  wire [63:0] regs_37_io_out; // @[RegFile.scala 66:20:@34774.4]
  wire  regs_37_io_enable; // @[RegFile.scala 66:20:@34774.4]
  wire  regs_38_clock; // @[RegFile.scala 66:20:@34788.4]
  wire  regs_38_reset; // @[RegFile.scala 66:20:@34788.4]
  wire [63:0] regs_38_io_in; // @[RegFile.scala 66:20:@34788.4]
  wire  regs_38_io_reset; // @[RegFile.scala 66:20:@34788.4]
  wire [63:0] regs_38_io_out; // @[RegFile.scala 66:20:@34788.4]
  wire  regs_38_io_enable; // @[RegFile.scala 66:20:@34788.4]
  wire  regs_39_clock; // @[RegFile.scala 66:20:@34802.4]
  wire  regs_39_reset; // @[RegFile.scala 66:20:@34802.4]
  wire [63:0] regs_39_io_in; // @[RegFile.scala 66:20:@34802.4]
  wire  regs_39_io_reset; // @[RegFile.scala 66:20:@34802.4]
  wire [63:0] regs_39_io_out; // @[RegFile.scala 66:20:@34802.4]
  wire  regs_39_io_enable; // @[RegFile.scala 66:20:@34802.4]
  wire  regs_40_clock; // @[RegFile.scala 66:20:@34816.4]
  wire  regs_40_reset; // @[RegFile.scala 66:20:@34816.4]
  wire [63:0] regs_40_io_in; // @[RegFile.scala 66:20:@34816.4]
  wire  regs_40_io_reset; // @[RegFile.scala 66:20:@34816.4]
  wire [63:0] regs_40_io_out; // @[RegFile.scala 66:20:@34816.4]
  wire  regs_40_io_enable; // @[RegFile.scala 66:20:@34816.4]
  wire  regs_41_clock; // @[RegFile.scala 66:20:@34830.4]
  wire  regs_41_reset; // @[RegFile.scala 66:20:@34830.4]
  wire [63:0] regs_41_io_in; // @[RegFile.scala 66:20:@34830.4]
  wire  regs_41_io_reset; // @[RegFile.scala 66:20:@34830.4]
  wire [63:0] regs_41_io_out; // @[RegFile.scala 66:20:@34830.4]
  wire  regs_41_io_enable; // @[RegFile.scala 66:20:@34830.4]
  wire  regs_42_clock; // @[RegFile.scala 66:20:@34844.4]
  wire  regs_42_reset; // @[RegFile.scala 66:20:@34844.4]
  wire [63:0] regs_42_io_in; // @[RegFile.scala 66:20:@34844.4]
  wire  regs_42_io_reset; // @[RegFile.scala 66:20:@34844.4]
  wire [63:0] regs_42_io_out; // @[RegFile.scala 66:20:@34844.4]
  wire  regs_42_io_enable; // @[RegFile.scala 66:20:@34844.4]
  wire  regs_43_clock; // @[RegFile.scala 66:20:@34858.4]
  wire  regs_43_reset; // @[RegFile.scala 66:20:@34858.4]
  wire [63:0] regs_43_io_in; // @[RegFile.scala 66:20:@34858.4]
  wire  regs_43_io_reset; // @[RegFile.scala 66:20:@34858.4]
  wire [63:0] regs_43_io_out; // @[RegFile.scala 66:20:@34858.4]
  wire  regs_43_io_enable; // @[RegFile.scala 66:20:@34858.4]
  wire  regs_44_clock; // @[RegFile.scala 66:20:@34872.4]
  wire  regs_44_reset; // @[RegFile.scala 66:20:@34872.4]
  wire [63:0] regs_44_io_in; // @[RegFile.scala 66:20:@34872.4]
  wire  regs_44_io_reset; // @[RegFile.scala 66:20:@34872.4]
  wire [63:0] regs_44_io_out; // @[RegFile.scala 66:20:@34872.4]
  wire  regs_44_io_enable; // @[RegFile.scala 66:20:@34872.4]
  wire  regs_45_clock; // @[RegFile.scala 66:20:@34886.4]
  wire  regs_45_reset; // @[RegFile.scala 66:20:@34886.4]
  wire [63:0] regs_45_io_in; // @[RegFile.scala 66:20:@34886.4]
  wire  regs_45_io_reset; // @[RegFile.scala 66:20:@34886.4]
  wire [63:0] regs_45_io_out; // @[RegFile.scala 66:20:@34886.4]
  wire  regs_45_io_enable; // @[RegFile.scala 66:20:@34886.4]
  wire  regs_46_clock; // @[RegFile.scala 66:20:@34900.4]
  wire  regs_46_reset; // @[RegFile.scala 66:20:@34900.4]
  wire [63:0] regs_46_io_in; // @[RegFile.scala 66:20:@34900.4]
  wire  regs_46_io_reset; // @[RegFile.scala 66:20:@34900.4]
  wire [63:0] regs_46_io_out; // @[RegFile.scala 66:20:@34900.4]
  wire  regs_46_io_enable; // @[RegFile.scala 66:20:@34900.4]
  wire  regs_47_clock; // @[RegFile.scala 66:20:@34914.4]
  wire  regs_47_reset; // @[RegFile.scala 66:20:@34914.4]
  wire [63:0] regs_47_io_in; // @[RegFile.scala 66:20:@34914.4]
  wire  regs_47_io_reset; // @[RegFile.scala 66:20:@34914.4]
  wire [63:0] regs_47_io_out; // @[RegFile.scala 66:20:@34914.4]
  wire  regs_47_io_enable; // @[RegFile.scala 66:20:@34914.4]
  wire  regs_48_clock; // @[RegFile.scala 66:20:@34928.4]
  wire  regs_48_reset; // @[RegFile.scala 66:20:@34928.4]
  wire [63:0] regs_48_io_in; // @[RegFile.scala 66:20:@34928.4]
  wire  regs_48_io_reset; // @[RegFile.scala 66:20:@34928.4]
  wire [63:0] regs_48_io_out; // @[RegFile.scala 66:20:@34928.4]
  wire  regs_48_io_enable; // @[RegFile.scala 66:20:@34928.4]
  wire  regs_49_clock; // @[RegFile.scala 66:20:@34942.4]
  wire  regs_49_reset; // @[RegFile.scala 66:20:@34942.4]
  wire [63:0] regs_49_io_in; // @[RegFile.scala 66:20:@34942.4]
  wire  regs_49_io_reset; // @[RegFile.scala 66:20:@34942.4]
  wire [63:0] regs_49_io_out; // @[RegFile.scala 66:20:@34942.4]
  wire  regs_49_io_enable; // @[RegFile.scala 66:20:@34942.4]
  wire  regs_50_clock; // @[RegFile.scala 66:20:@34956.4]
  wire  regs_50_reset; // @[RegFile.scala 66:20:@34956.4]
  wire [63:0] regs_50_io_in; // @[RegFile.scala 66:20:@34956.4]
  wire  regs_50_io_reset; // @[RegFile.scala 66:20:@34956.4]
  wire [63:0] regs_50_io_out; // @[RegFile.scala 66:20:@34956.4]
  wire  regs_50_io_enable; // @[RegFile.scala 66:20:@34956.4]
  wire  regs_51_clock; // @[RegFile.scala 66:20:@34970.4]
  wire  regs_51_reset; // @[RegFile.scala 66:20:@34970.4]
  wire [63:0] regs_51_io_in; // @[RegFile.scala 66:20:@34970.4]
  wire  regs_51_io_reset; // @[RegFile.scala 66:20:@34970.4]
  wire [63:0] regs_51_io_out; // @[RegFile.scala 66:20:@34970.4]
  wire  regs_51_io_enable; // @[RegFile.scala 66:20:@34970.4]
  wire  regs_52_clock; // @[RegFile.scala 66:20:@34984.4]
  wire  regs_52_reset; // @[RegFile.scala 66:20:@34984.4]
  wire [63:0] regs_52_io_in; // @[RegFile.scala 66:20:@34984.4]
  wire  regs_52_io_reset; // @[RegFile.scala 66:20:@34984.4]
  wire [63:0] regs_52_io_out; // @[RegFile.scala 66:20:@34984.4]
  wire  regs_52_io_enable; // @[RegFile.scala 66:20:@34984.4]
  wire  regs_53_clock; // @[RegFile.scala 66:20:@34998.4]
  wire  regs_53_reset; // @[RegFile.scala 66:20:@34998.4]
  wire [63:0] regs_53_io_in; // @[RegFile.scala 66:20:@34998.4]
  wire  regs_53_io_reset; // @[RegFile.scala 66:20:@34998.4]
  wire [63:0] regs_53_io_out; // @[RegFile.scala 66:20:@34998.4]
  wire  regs_53_io_enable; // @[RegFile.scala 66:20:@34998.4]
  wire  regs_54_clock; // @[RegFile.scala 66:20:@35012.4]
  wire  regs_54_reset; // @[RegFile.scala 66:20:@35012.4]
  wire [63:0] regs_54_io_in; // @[RegFile.scala 66:20:@35012.4]
  wire  regs_54_io_reset; // @[RegFile.scala 66:20:@35012.4]
  wire [63:0] regs_54_io_out; // @[RegFile.scala 66:20:@35012.4]
  wire  regs_54_io_enable; // @[RegFile.scala 66:20:@35012.4]
  wire  regs_55_clock; // @[RegFile.scala 66:20:@35026.4]
  wire  regs_55_reset; // @[RegFile.scala 66:20:@35026.4]
  wire [63:0] regs_55_io_in; // @[RegFile.scala 66:20:@35026.4]
  wire  regs_55_io_reset; // @[RegFile.scala 66:20:@35026.4]
  wire [63:0] regs_55_io_out; // @[RegFile.scala 66:20:@35026.4]
  wire  regs_55_io_enable; // @[RegFile.scala 66:20:@35026.4]
  wire  regs_56_clock; // @[RegFile.scala 66:20:@35040.4]
  wire  regs_56_reset; // @[RegFile.scala 66:20:@35040.4]
  wire [63:0] regs_56_io_in; // @[RegFile.scala 66:20:@35040.4]
  wire  regs_56_io_reset; // @[RegFile.scala 66:20:@35040.4]
  wire [63:0] regs_56_io_out; // @[RegFile.scala 66:20:@35040.4]
  wire  regs_56_io_enable; // @[RegFile.scala 66:20:@35040.4]
  wire  regs_57_clock; // @[RegFile.scala 66:20:@35054.4]
  wire  regs_57_reset; // @[RegFile.scala 66:20:@35054.4]
  wire [63:0] regs_57_io_in; // @[RegFile.scala 66:20:@35054.4]
  wire  regs_57_io_reset; // @[RegFile.scala 66:20:@35054.4]
  wire [63:0] regs_57_io_out; // @[RegFile.scala 66:20:@35054.4]
  wire  regs_57_io_enable; // @[RegFile.scala 66:20:@35054.4]
  wire  regs_58_clock; // @[RegFile.scala 66:20:@35068.4]
  wire  regs_58_reset; // @[RegFile.scala 66:20:@35068.4]
  wire [63:0] regs_58_io_in; // @[RegFile.scala 66:20:@35068.4]
  wire  regs_58_io_reset; // @[RegFile.scala 66:20:@35068.4]
  wire [63:0] regs_58_io_out; // @[RegFile.scala 66:20:@35068.4]
  wire  regs_58_io_enable; // @[RegFile.scala 66:20:@35068.4]
  wire  regs_59_clock; // @[RegFile.scala 66:20:@35082.4]
  wire  regs_59_reset; // @[RegFile.scala 66:20:@35082.4]
  wire [63:0] regs_59_io_in; // @[RegFile.scala 66:20:@35082.4]
  wire  regs_59_io_reset; // @[RegFile.scala 66:20:@35082.4]
  wire [63:0] regs_59_io_out; // @[RegFile.scala 66:20:@35082.4]
  wire  regs_59_io_enable; // @[RegFile.scala 66:20:@35082.4]
  wire  regs_60_clock; // @[RegFile.scala 66:20:@35096.4]
  wire  regs_60_reset; // @[RegFile.scala 66:20:@35096.4]
  wire [63:0] regs_60_io_in; // @[RegFile.scala 66:20:@35096.4]
  wire  regs_60_io_reset; // @[RegFile.scala 66:20:@35096.4]
  wire [63:0] regs_60_io_out; // @[RegFile.scala 66:20:@35096.4]
  wire  regs_60_io_enable; // @[RegFile.scala 66:20:@35096.4]
  wire  regs_61_clock; // @[RegFile.scala 66:20:@35110.4]
  wire  regs_61_reset; // @[RegFile.scala 66:20:@35110.4]
  wire [63:0] regs_61_io_in; // @[RegFile.scala 66:20:@35110.4]
  wire  regs_61_io_reset; // @[RegFile.scala 66:20:@35110.4]
  wire [63:0] regs_61_io_out; // @[RegFile.scala 66:20:@35110.4]
  wire  regs_61_io_enable; // @[RegFile.scala 66:20:@35110.4]
  wire  regs_62_clock; // @[RegFile.scala 66:20:@35124.4]
  wire  regs_62_reset; // @[RegFile.scala 66:20:@35124.4]
  wire [63:0] regs_62_io_in; // @[RegFile.scala 66:20:@35124.4]
  wire  regs_62_io_reset; // @[RegFile.scala 66:20:@35124.4]
  wire [63:0] regs_62_io_out; // @[RegFile.scala 66:20:@35124.4]
  wire  regs_62_io_enable; // @[RegFile.scala 66:20:@35124.4]
  wire  regs_63_clock; // @[RegFile.scala 66:20:@35138.4]
  wire  regs_63_reset; // @[RegFile.scala 66:20:@35138.4]
  wire [63:0] regs_63_io_in; // @[RegFile.scala 66:20:@35138.4]
  wire  regs_63_io_reset; // @[RegFile.scala 66:20:@35138.4]
  wire [63:0] regs_63_io_out; // @[RegFile.scala 66:20:@35138.4]
  wire  regs_63_io_enable; // @[RegFile.scala 66:20:@35138.4]
  wire  regs_64_clock; // @[RegFile.scala 66:20:@35152.4]
  wire  regs_64_reset; // @[RegFile.scala 66:20:@35152.4]
  wire [63:0] regs_64_io_in; // @[RegFile.scala 66:20:@35152.4]
  wire  regs_64_io_reset; // @[RegFile.scala 66:20:@35152.4]
  wire [63:0] regs_64_io_out; // @[RegFile.scala 66:20:@35152.4]
  wire  regs_64_io_enable; // @[RegFile.scala 66:20:@35152.4]
  wire  regs_65_clock; // @[RegFile.scala 66:20:@35166.4]
  wire  regs_65_reset; // @[RegFile.scala 66:20:@35166.4]
  wire [63:0] regs_65_io_in; // @[RegFile.scala 66:20:@35166.4]
  wire  regs_65_io_reset; // @[RegFile.scala 66:20:@35166.4]
  wire [63:0] regs_65_io_out; // @[RegFile.scala 66:20:@35166.4]
  wire  regs_65_io_enable; // @[RegFile.scala 66:20:@35166.4]
  wire  regs_66_clock; // @[RegFile.scala 66:20:@35180.4]
  wire  regs_66_reset; // @[RegFile.scala 66:20:@35180.4]
  wire [63:0] regs_66_io_in; // @[RegFile.scala 66:20:@35180.4]
  wire  regs_66_io_reset; // @[RegFile.scala 66:20:@35180.4]
  wire [63:0] regs_66_io_out; // @[RegFile.scala 66:20:@35180.4]
  wire  regs_66_io_enable; // @[RegFile.scala 66:20:@35180.4]
  wire  regs_67_clock; // @[RegFile.scala 66:20:@35194.4]
  wire  regs_67_reset; // @[RegFile.scala 66:20:@35194.4]
  wire [63:0] regs_67_io_in; // @[RegFile.scala 66:20:@35194.4]
  wire  regs_67_io_reset; // @[RegFile.scala 66:20:@35194.4]
  wire [63:0] regs_67_io_out; // @[RegFile.scala 66:20:@35194.4]
  wire  regs_67_io_enable; // @[RegFile.scala 66:20:@35194.4]
  wire  regs_68_clock; // @[RegFile.scala 66:20:@35208.4]
  wire  regs_68_reset; // @[RegFile.scala 66:20:@35208.4]
  wire [63:0] regs_68_io_in; // @[RegFile.scala 66:20:@35208.4]
  wire  regs_68_io_reset; // @[RegFile.scala 66:20:@35208.4]
  wire [63:0] regs_68_io_out; // @[RegFile.scala 66:20:@35208.4]
  wire  regs_68_io_enable; // @[RegFile.scala 66:20:@35208.4]
  wire  regs_69_clock; // @[RegFile.scala 66:20:@35222.4]
  wire  regs_69_reset; // @[RegFile.scala 66:20:@35222.4]
  wire [63:0] regs_69_io_in; // @[RegFile.scala 66:20:@35222.4]
  wire  regs_69_io_reset; // @[RegFile.scala 66:20:@35222.4]
  wire [63:0] regs_69_io_out; // @[RegFile.scala 66:20:@35222.4]
  wire  regs_69_io_enable; // @[RegFile.scala 66:20:@35222.4]
  wire  regs_70_clock; // @[RegFile.scala 66:20:@35236.4]
  wire  regs_70_reset; // @[RegFile.scala 66:20:@35236.4]
  wire [63:0] regs_70_io_in; // @[RegFile.scala 66:20:@35236.4]
  wire  regs_70_io_reset; // @[RegFile.scala 66:20:@35236.4]
  wire [63:0] regs_70_io_out; // @[RegFile.scala 66:20:@35236.4]
  wire  regs_70_io_enable; // @[RegFile.scala 66:20:@35236.4]
  wire  regs_71_clock; // @[RegFile.scala 66:20:@35250.4]
  wire  regs_71_reset; // @[RegFile.scala 66:20:@35250.4]
  wire [63:0] regs_71_io_in; // @[RegFile.scala 66:20:@35250.4]
  wire  regs_71_io_reset; // @[RegFile.scala 66:20:@35250.4]
  wire [63:0] regs_71_io_out; // @[RegFile.scala 66:20:@35250.4]
  wire  regs_71_io_enable; // @[RegFile.scala 66:20:@35250.4]
  wire  regs_72_clock; // @[RegFile.scala 66:20:@35264.4]
  wire  regs_72_reset; // @[RegFile.scala 66:20:@35264.4]
  wire [63:0] regs_72_io_in; // @[RegFile.scala 66:20:@35264.4]
  wire  regs_72_io_reset; // @[RegFile.scala 66:20:@35264.4]
  wire [63:0] regs_72_io_out; // @[RegFile.scala 66:20:@35264.4]
  wire  regs_72_io_enable; // @[RegFile.scala 66:20:@35264.4]
  wire  regs_73_clock; // @[RegFile.scala 66:20:@35278.4]
  wire  regs_73_reset; // @[RegFile.scala 66:20:@35278.4]
  wire [63:0] regs_73_io_in; // @[RegFile.scala 66:20:@35278.4]
  wire  regs_73_io_reset; // @[RegFile.scala 66:20:@35278.4]
  wire [63:0] regs_73_io_out; // @[RegFile.scala 66:20:@35278.4]
  wire  regs_73_io_enable; // @[RegFile.scala 66:20:@35278.4]
  wire  regs_74_clock; // @[RegFile.scala 66:20:@35292.4]
  wire  regs_74_reset; // @[RegFile.scala 66:20:@35292.4]
  wire [63:0] regs_74_io_in; // @[RegFile.scala 66:20:@35292.4]
  wire  regs_74_io_reset; // @[RegFile.scala 66:20:@35292.4]
  wire [63:0] regs_74_io_out; // @[RegFile.scala 66:20:@35292.4]
  wire  regs_74_io_enable; // @[RegFile.scala 66:20:@35292.4]
  wire  regs_75_clock; // @[RegFile.scala 66:20:@35306.4]
  wire  regs_75_reset; // @[RegFile.scala 66:20:@35306.4]
  wire [63:0] regs_75_io_in; // @[RegFile.scala 66:20:@35306.4]
  wire  regs_75_io_reset; // @[RegFile.scala 66:20:@35306.4]
  wire [63:0] regs_75_io_out; // @[RegFile.scala 66:20:@35306.4]
  wire  regs_75_io_enable; // @[RegFile.scala 66:20:@35306.4]
  wire  regs_76_clock; // @[RegFile.scala 66:20:@35320.4]
  wire  regs_76_reset; // @[RegFile.scala 66:20:@35320.4]
  wire [63:0] regs_76_io_in; // @[RegFile.scala 66:20:@35320.4]
  wire  regs_76_io_reset; // @[RegFile.scala 66:20:@35320.4]
  wire [63:0] regs_76_io_out; // @[RegFile.scala 66:20:@35320.4]
  wire  regs_76_io_enable; // @[RegFile.scala 66:20:@35320.4]
  wire  regs_77_clock; // @[RegFile.scala 66:20:@35334.4]
  wire  regs_77_reset; // @[RegFile.scala 66:20:@35334.4]
  wire [63:0] regs_77_io_in; // @[RegFile.scala 66:20:@35334.4]
  wire  regs_77_io_reset; // @[RegFile.scala 66:20:@35334.4]
  wire [63:0] regs_77_io_out; // @[RegFile.scala 66:20:@35334.4]
  wire  regs_77_io_enable; // @[RegFile.scala 66:20:@35334.4]
  wire  regs_78_clock; // @[RegFile.scala 66:20:@35348.4]
  wire  regs_78_reset; // @[RegFile.scala 66:20:@35348.4]
  wire [63:0] regs_78_io_in; // @[RegFile.scala 66:20:@35348.4]
  wire  regs_78_io_reset; // @[RegFile.scala 66:20:@35348.4]
  wire [63:0] regs_78_io_out; // @[RegFile.scala 66:20:@35348.4]
  wire  regs_78_io_enable; // @[RegFile.scala 66:20:@35348.4]
  wire  regs_79_clock; // @[RegFile.scala 66:20:@35362.4]
  wire  regs_79_reset; // @[RegFile.scala 66:20:@35362.4]
  wire [63:0] regs_79_io_in; // @[RegFile.scala 66:20:@35362.4]
  wire  regs_79_io_reset; // @[RegFile.scala 66:20:@35362.4]
  wire [63:0] regs_79_io_out; // @[RegFile.scala 66:20:@35362.4]
  wire  regs_79_io_enable; // @[RegFile.scala 66:20:@35362.4]
  wire  regs_80_clock; // @[RegFile.scala 66:20:@35376.4]
  wire  regs_80_reset; // @[RegFile.scala 66:20:@35376.4]
  wire [63:0] regs_80_io_in; // @[RegFile.scala 66:20:@35376.4]
  wire  regs_80_io_reset; // @[RegFile.scala 66:20:@35376.4]
  wire [63:0] regs_80_io_out; // @[RegFile.scala 66:20:@35376.4]
  wire  regs_80_io_enable; // @[RegFile.scala 66:20:@35376.4]
  wire  regs_81_clock; // @[RegFile.scala 66:20:@35390.4]
  wire  regs_81_reset; // @[RegFile.scala 66:20:@35390.4]
  wire [63:0] regs_81_io_in; // @[RegFile.scala 66:20:@35390.4]
  wire  regs_81_io_reset; // @[RegFile.scala 66:20:@35390.4]
  wire [63:0] regs_81_io_out; // @[RegFile.scala 66:20:@35390.4]
  wire  regs_81_io_enable; // @[RegFile.scala 66:20:@35390.4]
  wire  regs_82_clock; // @[RegFile.scala 66:20:@35404.4]
  wire  regs_82_reset; // @[RegFile.scala 66:20:@35404.4]
  wire [63:0] regs_82_io_in; // @[RegFile.scala 66:20:@35404.4]
  wire  regs_82_io_reset; // @[RegFile.scala 66:20:@35404.4]
  wire [63:0] regs_82_io_out; // @[RegFile.scala 66:20:@35404.4]
  wire  regs_82_io_enable; // @[RegFile.scala 66:20:@35404.4]
  wire  regs_83_clock; // @[RegFile.scala 66:20:@35418.4]
  wire  regs_83_reset; // @[RegFile.scala 66:20:@35418.4]
  wire [63:0] regs_83_io_in; // @[RegFile.scala 66:20:@35418.4]
  wire  regs_83_io_reset; // @[RegFile.scala 66:20:@35418.4]
  wire [63:0] regs_83_io_out; // @[RegFile.scala 66:20:@35418.4]
  wire  regs_83_io_enable; // @[RegFile.scala 66:20:@35418.4]
  wire  regs_84_clock; // @[RegFile.scala 66:20:@35432.4]
  wire  regs_84_reset; // @[RegFile.scala 66:20:@35432.4]
  wire [63:0] regs_84_io_in; // @[RegFile.scala 66:20:@35432.4]
  wire  regs_84_io_reset; // @[RegFile.scala 66:20:@35432.4]
  wire [63:0] regs_84_io_out; // @[RegFile.scala 66:20:@35432.4]
  wire  regs_84_io_enable; // @[RegFile.scala 66:20:@35432.4]
  wire  regs_85_clock; // @[RegFile.scala 66:20:@35446.4]
  wire  regs_85_reset; // @[RegFile.scala 66:20:@35446.4]
  wire [63:0] regs_85_io_in; // @[RegFile.scala 66:20:@35446.4]
  wire  regs_85_io_reset; // @[RegFile.scala 66:20:@35446.4]
  wire [63:0] regs_85_io_out; // @[RegFile.scala 66:20:@35446.4]
  wire  regs_85_io_enable; // @[RegFile.scala 66:20:@35446.4]
  wire  regs_86_clock; // @[RegFile.scala 66:20:@35460.4]
  wire  regs_86_reset; // @[RegFile.scala 66:20:@35460.4]
  wire [63:0] regs_86_io_in; // @[RegFile.scala 66:20:@35460.4]
  wire  regs_86_io_reset; // @[RegFile.scala 66:20:@35460.4]
  wire [63:0] regs_86_io_out; // @[RegFile.scala 66:20:@35460.4]
  wire  regs_86_io_enable; // @[RegFile.scala 66:20:@35460.4]
  wire  regs_87_clock; // @[RegFile.scala 66:20:@35474.4]
  wire  regs_87_reset; // @[RegFile.scala 66:20:@35474.4]
  wire [63:0] regs_87_io_in; // @[RegFile.scala 66:20:@35474.4]
  wire  regs_87_io_reset; // @[RegFile.scala 66:20:@35474.4]
  wire [63:0] regs_87_io_out; // @[RegFile.scala 66:20:@35474.4]
  wire  regs_87_io_enable; // @[RegFile.scala 66:20:@35474.4]
  wire  regs_88_clock; // @[RegFile.scala 66:20:@35488.4]
  wire  regs_88_reset; // @[RegFile.scala 66:20:@35488.4]
  wire [63:0] regs_88_io_in; // @[RegFile.scala 66:20:@35488.4]
  wire  regs_88_io_reset; // @[RegFile.scala 66:20:@35488.4]
  wire [63:0] regs_88_io_out; // @[RegFile.scala 66:20:@35488.4]
  wire  regs_88_io_enable; // @[RegFile.scala 66:20:@35488.4]
  wire  regs_89_clock; // @[RegFile.scala 66:20:@35502.4]
  wire  regs_89_reset; // @[RegFile.scala 66:20:@35502.4]
  wire [63:0] regs_89_io_in; // @[RegFile.scala 66:20:@35502.4]
  wire  regs_89_io_reset; // @[RegFile.scala 66:20:@35502.4]
  wire [63:0] regs_89_io_out; // @[RegFile.scala 66:20:@35502.4]
  wire  regs_89_io_enable; // @[RegFile.scala 66:20:@35502.4]
  wire  regs_90_clock; // @[RegFile.scala 66:20:@35516.4]
  wire  regs_90_reset; // @[RegFile.scala 66:20:@35516.4]
  wire [63:0] regs_90_io_in; // @[RegFile.scala 66:20:@35516.4]
  wire  regs_90_io_reset; // @[RegFile.scala 66:20:@35516.4]
  wire [63:0] regs_90_io_out; // @[RegFile.scala 66:20:@35516.4]
  wire  regs_90_io_enable; // @[RegFile.scala 66:20:@35516.4]
  wire  regs_91_clock; // @[RegFile.scala 66:20:@35530.4]
  wire  regs_91_reset; // @[RegFile.scala 66:20:@35530.4]
  wire [63:0] regs_91_io_in; // @[RegFile.scala 66:20:@35530.4]
  wire  regs_91_io_reset; // @[RegFile.scala 66:20:@35530.4]
  wire [63:0] regs_91_io_out; // @[RegFile.scala 66:20:@35530.4]
  wire  regs_91_io_enable; // @[RegFile.scala 66:20:@35530.4]
  wire  regs_92_clock; // @[RegFile.scala 66:20:@35544.4]
  wire  regs_92_reset; // @[RegFile.scala 66:20:@35544.4]
  wire [63:0] regs_92_io_in; // @[RegFile.scala 66:20:@35544.4]
  wire  regs_92_io_reset; // @[RegFile.scala 66:20:@35544.4]
  wire [63:0] regs_92_io_out; // @[RegFile.scala 66:20:@35544.4]
  wire  regs_92_io_enable; // @[RegFile.scala 66:20:@35544.4]
  wire  regs_93_clock; // @[RegFile.scala 66:20:@35558.4]
  wire  regs_93_reset; // @[RegFile.scala 66:20:@35558.4]
  wire [63:0] regs_93_io_in; // @[RegFile.scala 66:20:@35558.4]
  wire  regs_93_io_reset; // @[RegFile.scala 66:20:@35558.4]
  wire [63:0] regs_93_io_out; // @[RegFile.scala 66:20:@35558.4]
  wire  regs_93_io_enable; // @[RegFile.scala 66:20:@35558.4]
  wire  regs_94_clock; // @[RegFile.scala 66:20:@35572.4]
  wire  regs_94_reset; // @[RegFile.scala 66:20:@35572.4]
  wire [63:0] regs_94_io_in; // @[RegFile.scala 66:20:@35572.4]
  wire  regs_94_io_reset; // @[RegFile.scala 66:20:@35572.4]
  wire [63:0] regs_94_io_out; // @[RegFile.scala 66:20:@35572.4]
  wire  regs_94_io_enable; // @[RegFile.scala 66:20:@35572.4]
  wire  regs_95_clock; // @[RegFile.scala 66:20:@35586.4]
  wire  regs_95_reset; // @[RegFile.scala 66:20:@35586.4]
  wire [63:0] regs_95_io_in; // @[RegFile.scala 66:20:@35586.4]
  wire  regs_95_io_reset; // @[RegFile.scala 66:20:@35586.4]
  wire [63:0] regs_95_io_out; // @[RegFile.scala 66:20:@35586.4]
  wire  regs_95_io_enable; // @[RegFile.scala 66:20:@35586.4]
  wire  regs_96_clock; // @[RegFile.scala 66:20:@35600.4]
  wire  regs_96_reset; // @[RegFile.scala 66:20:@35600.4]
  wire [63:0] regs_96_io_in; // @[RegFile.scala 66:20:@35600.4]
  wire  regs_96_io_reset; // @[RegFile.scala 66:20:@35600.4]
  wire [63:0] regs_96_io_out; // @[RegFile.scala 66:20:@35600.4]
  wire  regs_96_io_enable; // @[RegFile.scala 66:20:@35600.4]
  wire  regs_97_clock; // @[RegFile.scala 66:20:@35614.4]
  wire  regs_97_reset; // @[RegFile.scala 66:20:@35614.4]
  wire [63:0] regs_97_io_in; // @[RegFile.scala 66:20:@35614.4]
  wire  regs_97_io_reset; // @[RegFile.scala 66:20:@35614.4]
  wire [63:0] regs_97_io_out; // @[RegFile.scala 66:20:@35614.4]
  wire  regs_97_io_enable; // @[RegFile.scala 66:20:@35614.4]
  wire  regs_98_clock; // @[RegFile.scala 66:20:@35628.4]
  wire  regs_98_reset; // @[RegFile.scala 66:20:@35628.4]
  wire [63:0] regs_98_io_in; // @[RegFile.scala 66:20:@35628.4]
  wire  regs_98_io_reset; // @[RegFile.scala 66:20:@35628.4]
  wire [63:0] regs_98_io_out; // @[RegFile.scala 66:20:@35628.4]
  wire  regs_98_io_enable; // @[RegFile.scala 66:20:@35628.4]
  wire  regs_99_clock; // @[RegFile.scala 66:20:@35642.4]
  wire  regs_99_reset; // @[RegFile.scala 66:20:@35642.4]
  wire [63:0] regs_99_io_in; // @[RegFile.scala 66:20:@35642.4]
  wire  regs_99_io_reset; // @[RegFile.scala 66:20:@35642.4]
  wire [63:0] regs_99_io_out; // @[RegFile.scala 66:20:@35642.4]
  wire  regs_99_io_enable; // @[RegFile.scala 66:20:@35642.4]
  wire  regs_100_clock; // @[RegFile.scala 66:20:@35656.4]
  wire  regs_100_reset; // @[RegFile.scala 66:20:@35656.4]
  wire [63:0] regs_100_io_in; // @[RegFile.scala 66:20:@35656.4]
  wire  regs_100_io_reset; // @[RegFile.scala 66:20:@35656.4]
  wire [63:0] regs_100_io_out; // @[RegFile.scala 66:20:@35656.4]
  wire  regs_100_io_enable; // @[RegFile.scala 66:20:@35656.4]
  wire  regs_101_clock; // @[RegFile.scala 66:20:@35670.4]
  wire  regs_101_reset; // @[RegFile.scala 66:20:@35670.4]
  wire [63:0] regs_101_io_in; // @[RegFile.scala 66:20:@35670.4]
  wire  regs_101_io_reset; // @[RegFile.scala 66:20:@35670.4]
  wire [63:0] regs_101_io_out; // @[RegFile.scala 66:20:@35670.4]
  wire  regs_101_io_enable; // @[RegFile.scala 66:20:@35670.4]
  wire  regs_102_clock; // @[RegFile.scala 66:20:@35684.4]
  wire  regs_102_reset; // @[RegFile.scala 66:20:@35684.4]
  wire [63:0] regs_102_io_in; // @[RegFile.scala 66:20:@35684.4]
  wire  regs_102_io_reset; // @[RegFile.scala 66:20:@35684.4]
  wire [63:0] regs_102_io_out; // @[RegFile.scala 66:20:@35684.4]
  wire  regs_102_io_enable; // @[RegFile.scala 66:20:@35684.4]
  wire  regs_103_clock; // @[RegFile.scala 66:20:@35698.4]
  wire  regs_103_reset; // @[RegFile.scala 66:20:@35698.4]
  wire [63:0] regs_103_io_in; // @[RegFile.scala 66:20:@35698.4]
  wire  regs_103_io_reset; // @[RegFile.scala 66:20:@35698.4]
  wire [63:0] regs_103_io_out; // @[RegFile.scala 66:20:@35698.4]
  wire  regs_103_io_enable; // @[RegFile.scala 66:20:@35698.4]
  wire  regs_104_clock; // @[RegFile.scala 66:20:@35712.4]
  wire  regs_104_reset; // @[RegFile.scala 66:20:@35712.4]
  wire [63:0] regs_104_io_in; // @[RegFile.scala 66:20:@35712.4]
  wire  regs_104_io_reset; // @[RegFile.scala 66:20:@35712.4]
  wire [63:0] regs_104_io_out; // @[RegFile.scala 66:20:@35712.4]
  wire  regs_104_io_enable; // @[RegFile.scala 66:20:@35712.4]
  wire  regs_105_clock; // @[RegFile.scala 66:20:@35726.4]
  wire  regs_105_reset; // @[RegFile.scala 66:20:@35726.4]
  wire [63:0] regs_105_io_in; // @[RegFile.scala 66:20:@35726.4]
  wire  regs_105_io_reset; // @[RegFile.scala 66:20:@35726.4]
  wire [63:0] regs_105_io_out; // @[RegFile.scala 66:20:@35726.4]
  wire  regs_105_io_enable; // @[RegFile.scala 66:20:@35726.4]
  wire  regs_106_clock; // @[RegFile.scala 66:20:@35740.4]
  wire  regs_106_reset; // @[RegFile.scala 66:20:@35740.4]
  wire [63:0] regs_106_io_in; // @[RegFile.scala 66:20:@35740.4]
  wire  regs_106_io_reset; // @[RegFile.scala 66:20:@35740.4]
  wire [63:0] regs_106_io_out; // @[RegFile.scala 66:20:@35740.4]
  wire  regs_106_io_enable; // @[RegFile.scala 66:20:@35740.4]
  wire  regs_107_clock; // @[RegFile.scala 66:20:@35754.4]
  wire  regs_107_reset; // @[RegFile.scala 66:20:@35754.4]
  wire [63:0] regs_107_io_in; // @[RegFile.scala 66:20:@35754.4]
  wire  regs_107_io_reset; // @[RegFile.scala 66:20:@35754.4]
  wire [63:0] regs_107_io_out; // @[RegFile.scala 66:20:@35754.4]
  wire  regs_107_io_enable; // @[RegFile.scala 66:20:@35754.4]
  wire  regs_108_clock; // @[RegFile.scala 66:20:@35768.4]
  wire  regs_108_reset; // @[RegFile.scala 66:20:@35768.4]
  wire [63:0] regs_108_io_in; // @[RegFile.scala 66:20:@35768.4]
  wire  regs_108_io_reset; // @[RegFile.scala 66:20:@35768.4]
  wire [63:0] regs_108_io_out; // @[RegFile.scala 66:20:@35768.4]
  wire  regs_108_io_enable; // @[RegFile.scala 66:20:@35768.4]
  wire  regs_109_clock; // @[RegFile.scala 66:20:@35782.4]
  wire  regs_109_reset; // @[RegFile.scala 66:20:@35782.4]
  wire [63:0] regs_109_io_in; // @[RegFile.scala 66:20:@35782.4]
  wire  regs_109_io_reset; // @[RegFile.scala 66:20:@35782.4]
  wire [63:0] regs_109_io_out; // @[RegFile.scala 66:20:@35782.4]
  wire  regs_109_io_enable; // @[RegFile.scala 66:20:@35782.4]
  wire  regs_110_clock; // @[RegFile.scala 66:20:@35796.4]
  wire  regs_110_reset; // @[RegFile.scala 66:20:@35796.4]
  wire [63:0] regs_110_io_in; // @[RegFile.scala 66:20:@35796.4]
  wire  regs_110_io_reset; // @[RegFile.scala 66:20:@35796.4]
  wire [63:0] regs_110_io_out; // @[RegFile.scala 66:20:@35796.4]
  wire  regs_110_io_enable; // @[RegFile.scala 66:20:@35796.4]
  wire  regs_111_clock; // @[RegFile.scala 66:20:@35810.4]
  wire  regs_111_reset; // @[RegFile.scala 66:20:@35810.4]
  wire [63:0] regs_111_io_in; // @[RegFile.scala 66:20:@35810.4]
  wire  regs_111_io_reset; // @[RegFile.scala 66:20:@35810.4]
  wire [63:0] regs_111_io_out; // @[RegFile.scala 66:20:@35810.4]
  wire  regs_111_io_enable; // @[RegFile.scala 66:20:@35810.4]
  wire  regs_112_clock; // @[RegFile.scala 66:20:@35824.4]
  wire  regs_112_reset; // @[RegFile.scala 66:20:@35824.4]
  wire [63:0] regs_112_io_in; // @[RegFile.scala 66:20:@35824.4]
  wire  regs_112_io_reset; // @[RegFile.scala 66:20:@35824.4]
  wire [63:0] regs_112_io_out; // @[RegFile.scala 66:20:@35824.4]
  wire  regs_112_io_enable; // @[RegFile.scala 66:20:@35824.4]
  wire  regs_113_clock; // @[RegFile.scala 66:20:@35838.4]
  wire  regs_113_reset; // @[RegFile.scala 66:20:@35838.4]
  wire [63:0] regs_113_io_in; // @[RegFile.scala 66:20:@35838.4]
  wire  regs_113_io_reset; // @[RegFile.scala 66:20:@35838.4]
  wire [63:0] regs_113_io_out; // @[RegFile.scala 66:20:@35838.4]
  wire  regs_113_io_enable; // @[RegFile.scala 66:20:@35838.4]
  wire  regs_114_clock; // @[RegFile.scala 66:20:@35852.4]
  wire  regs_114_reset; // @[RegFile.scala 66:20:@35852.4]
  wire [63:0] regs_114_io_in; // @[RegFile.scala 66:20:@35852.4]
  wire  regs_114_io_reset; // @[RegFile.scala 66:20:@35852.4]
  wire [63:0] regs_114_io_out; // @[RegFile.scala 66:20:@35852.4]
  wire  regs_114_io_enable; // @[RegFile.scala 66:20:@35852.4]
  wire  regs_115_clock; // @[RegFile.scala 66:20:@35866.4]
  wire  regs_115_reset; // @[RegFile.scala 66:20:@35866.4]
  wire [63:0] regs_115_io_in; // @[RegFile.scala 66:20:@35866.4]
  wire  regs_115_io_reset; // @[RegFile.scala 66:20:@35866.4]
  wire [63:0] regs_115_io_out; // @[RegFile.scala 66:20:@35866.4]
  wire  regs_115_io_enable; // @[RegFile.scala 66:20:@35866.4]
  wire  regs_116_clock; // @[RegFile.scala 66:20:@35880.4]
  wire  regs_116_reset; // @[RegFile.scala 66:20:@35880.4]
  wire [63:0] regs_116_io_in; // @[RegFile.scala 66:20:@35880.4]
  wire  regs_116_io_reset; // @[RegFile.scala 66:20:@35880.4]
  wire [63:0] regs_116_io_out; // @[RegFile.scala 66:20:@35880.4]
  wire  regs_116_io_enable; // @[RegFile.scala 66:20:@35880.4]
  wire  regs_117_clock; // @[RegFile.scala 66:20:@35894.4]
  wire  regs_117_reset; // @[RegFile.scala 66:20:@35894.4]
  wire [63:0] regs_117_io_in; // @[RegFile.scala 66:20:@35894.4]
  wire  regs_117_io_reset; // @[RegFile.scala 66:20:@35894.4]
  wire [63:0] regs_117_io_out; // @[RegFile.scala 66:20:@35894.4]
  wire  regs_117_io_enable; // @[RegFile.scala 66:20:@35894.4]
  wire  regs_118_clock; // @[RegFile.scala 66:20:@35908.4]
  wire  regs_118_reset; // @[RegFile.scala 66:20:@35908.4]
  wire [63:0] regs_118_io_in; // @[RegFile.scala 66:20:@35908.4]
  wire  regs_118_io_reset; // @[RegFile.scala 66:20:@35908.4]
  wire [63:0] regs_118_io_out; // @[RegFile.scala 66:20:@35908.4]
  wire  regs_118_io_enable; // @[RegFile.scala 66:20:@35908.4]
  wire  regs_119_clock; // @[RegFile.scala 66:20:@35922.4]
  wire  regs_119_reset; // @[RegFile.scala 66:20:@35922.4]
  wire [63:0] regs_119_io_in; // @[RegFile.scala 66:20:@35922.4]
  wire  regs_119_io_reset; // @[RegFile.scala 66:20:@35922.4]
  wire [63:0] regs_119_io_out; // @[RegFile.scala 66:20:@35922.4]
  wire  regs_119_io_enable; // @[RegFile.scala 66:20:@35922.4]
  wire  regs_120_clock; // @[RegFile.scala 66:20:@35936.4]
  wire  regs_120_reset; // @[RegFile.scala 66:20:@35936.4]
  wire [63:0] regs_120_io_in; // @[RegFile.scala 66:20:@35936.4]
  wire  regs_120_io_reset; // @[RegFile.scala 66:20:@35936.4]
  wire [63:0] regs_120_io_out; // @[RegFile.scala 66:20:@35936.4]
  wire  regs_120_io_enable; // @[RegFile.scala 66:20:@35936.4]
  wire  regs_121_clock; // @[RegFile.scala 66:20:@35950.4]
  wire  regs_121_reset; // @[RegFile.scala 66:20:@35950.4]
  wire [63:0] regs_121_io_in; // @[RegFile.scala 66:20:@35950.4]
  wire  regs_121_io_reset; // @[RegFile.scala 66:20:@35950.4]
  wire [63:0] regs_121_io_out; // @[RegFile.scala 66:20:@35950.4]
  wire  regs_121_io_enable; // @[RegFile.scala 66:20:@35950.4]
  wire  regs_122_clock; // @[RegFile.scala 66:20:@35964.4]
  wire  regs_122_reset; // @[RegFile.scala 66:20:@35964.4]
  wire [63:0] regs_122_io_in; // @[RegFile.scala 66:20:@35964.4]
  wire  regs_122_io_reset; // @[RegFile.scala 66:20:@35964.4]
  wire [63:0] regs_122_io_out; // @[RegFile.scala 66:20:@35964.4]
  wire  regs_122_io_enable; // @[RegFile.scala 66:20:@35964.4]
  wire  regs_123_clock; // @[RegFile.scala 66:20:@35978.4]
  wire  regs_123_reset; // @[RegFile.scala 66:20:@35978.4]
  wire [63:0] regs_123_io_in; // @[RegFile.scala 66:20:@35978.4]
  wire  regs_123_io_reset; // @[RegFile.scala 66:20:@35978.4]
  wire [63:0] regs_123_io_out; // @[RegFile.scala 66:20:@35978.4]
  wire  regs_123_io_enable; // @[RegFile.scala 66:20:@35978.4]
  wire  regs_124_clock; // @[RegFile.scala 66:20:@35992.4]
  wire  regs_124_reset; // @[RegFile.scala 66:20:@35992.4]
  wire [63:0] regs_124_io_in; // @[RegFile.scala 66:20:@35992.4]
  wire  regs_124_io_reset; // @[RegFile.scala 66:20:@35992.4]
  wire [63:0] regs_124_io_out; // @[RegFile.scala 66:20:@35992.4]
  wire  regs_124_io_enable; // @[RegFile.scala 66:20:@35992.4]
  wire  regs_125_clock; // @[RegFile.scala 66:20:@36006.4]
  wire  regs_125_reset; // @[RegFile.scala 66:20:@36006.4]
  wire [63:0] regs_125_io_in; // @[RegFile.scala 66:20:@36006.4]
  wire  regs_125_io_reset; // @[RegFile.scala 66:20:@36006.4]
  wire [63:0] regs_125_io_out; // @[RegFile.scala 66:20:@36006.4]
  wire  regs_125_io_enable; // @[RegFile.scala 66:20:@36006.4]
  wire  regs_126_clock; // @[RegFile.scala 66:20:@36020.4]
  wire  regs_126_reset; // @[RegFile.scala 66:20:@36020.4]
  wire [63:0] regs_126_io_in; // @[RegFile.scala 66:20:@36020.4]
  wire  regs_126_io_reset; // @[RegFile.scala 66:20:@36020.4]
  wire [63:0] regs_126_io_out; // @[RegFile.scala 66:20:@36020.4]
  wire  regs_126_io_enable; // @[RegFile.scala 66:20:@36020.4]
  wire  regs_127_clock; // @[RegFile.scala 66:20:@36034.4]
  wire  regs_127_reset; // @[RegFile.scala 66:20:@36034.4]
  wire [63:0] regs_127_io_in; // @[RegFile.scala 66:20:@36034.4]
  wire  regs_127_io_reset; // @[RegFile.scala 66:20:@36034.4]
  wire [63:0] regs_127_io_out; // @[RegFile.scala 66:20:@36034.4]
  wire  regs_127_io_enable; // @[RegFile.scala 66:20:@36034.4]
  wire  regs_128_clock; // @[RegFile.scala 66:20:@36048.4]
  wire  regs_128_reset; // @[RegFile.scala 66:20:@36048.4]
  wire [63:0] regs_128_io_in; // @[RegFile.scala 66:20:@36048.4]
  wire  regs_128_io_reset; // @[RegFile.scala 66:20:@36048.4]
  wire [63:0] regs_128_io_out; // @[RegFile.scala 66:20:@36048.4]
  wire  regs_128_io_enable; // @[RegFile.scala 66:20:@36048.4]
  wire  regs_129_clock; // @[RegFile.scala 66:20:@36062.4]
  wire  regs_129_reset; // @[RegFile.scala 66:20:@36062.4]
  wire [63:0] regs_129_io_in; // @[RegFile.scala 66:20:@36062.4]
  wire  regs_129_io_reset; // @[RegFile.scala 66:20:@36062.4]
  wire [63:0] regs_129_io_out; // @[RegFile.scala 66:20:@36062.4]
  wire  regs_129_io_enable; // @[RegFile.scala 66:20:@36062.4]
  wire  regs_130_clock; // @[RegFile.scala 66:20:@36076.4]
  wire  regs_130_reset; // @[RegFile.scala 66:20:@36076.4]
  wire [63:0] regs_130_io_in; // @[RegFile.scala 66:20:@36076.4]
  wire  regs_130_io_reset; // @[RegFile.scala 66:20:@36076.4]
  wire [63:0] regs_130_io_out; // @[RegFile.scala 66:20:@36076.4]
  wire  regs_130_io_enable; // @[RegFile.scala 66:20:@36076.4]
  wire  regs_131_clock; // @[RegFile.scala 66:20:@36090.4]
  wire  regs_131_reset; // @[RegFile.scala 66:20:@36090.4]
  wire [63:0] regs_131_io_in; // @[RegFile.scala 66:20:@36090.4]
  wire  regs_131_io_reset; // @[RegFile.scala 66:20:@36090.4]
  wire [63:0] regs_131_io_out; // @[RegFile.scala 66:20:@36090.4]
  wire  regs_131_io_enable; // @[RegFile.scala 66:20:@36090.4]
  wire  regs_132_clock; // @[RegFile.scala 66:20:@36104.4]
  wire  regs_132_reset; // @[RegFile.scala 66:20:@36104.4]
  wire [63:0] regs_132_io_in; // @[RegFile.scala 66:20:@36104.4]
  wire  regs_132_io_reset; // @[RegFile.scala 66:20:@36104.4]
  wire [63:0] regs_132_io_out; // @[RegFile.scala 66:20:@36104.4]
  wire  regs_132_io_enable; // @[RegFile.scala 66:20:@36104.4]
  wire  regs_133_clock; // @[RegFile.scala 66:20:@36118.4]
  wire  regs_133_reset; // @[RegFile.scala 66:20:@36118.4]
  wire [63:0] regs_133_io_in; // @[RegFile.scala 66:20:@36118.4]
  wire  regs_133_io_reset; // @[RegFile.scala 66:20:@36118.4]
  wire [63:0] regs_133_io_out; // @[RegFile.scala 66:20:@36118.4]
  wire  regs_133_io_enable; // @[RegFile.scala 66:20:@36118.4]
  wire  regs_134_clock; // @[RegFile.scala 66:20:@36132.4]
  wire  regs_134_reset; // @[RegFile.scala 66:20:@36132.4]
  wire [63:0] regs_134_io_in; // @[RegFile.scala 66:20:@36132.4]
  wire  regs_134_io_reset; // @[RegFile.scala 66:20:@36132.4]
  wire [63:0] regs_134_io_out; // @[RegFile.scala 66:20:@36132.4]
  wire  regs_134_io_enable; // @[RegFile.scala 66:20:@36132.4]
  wire  regs_135_clock; // @[RegFile.scala 66:20:@36146.4]
  wire  regs_135_reset; // @[RegFile.scala 66:20:@36146.4]
  wire [63:0] regs_135_io_in; // @[RegFile.scala 66:20:@36146.4]
  wire  regs_135_io_reset; // @[RegFile.scala 66:20:@36146.4]
  wire [63:0] regs_135_io_out; // @[RegFile.scala 66:20:@36146.4]
  wire  regs_135_io_enable; // @[RegFile.scala 66:20:@36146.4]
  wire  regs_136_clock; // @[RegFile.scala 66:20:@36160.4]
  wire  regs_136_reset; // @[RegFile.scala 66:20:@36160.4]
  wire [63:0] regs_136_io_in; // @[RegFile.scala 66:20:@36160.4]
  wire  regs_136_io_reset; // @[RegFile.scala 66:20:@36160.4]
  wire [63:0] regs_136_io_out; // @[RegFile.scala 66:20:@36160.4]
  wire  regs_136_io_enable; // @[RegFile.scala 66:20:@36160.4]
  wire  regs_137_clock; // @[RegFile.scala 66:20:@36174.4]
  wire  regs_137_reset; // @[RegFile.scala 66:20:@36174.4]
  wire [63:0] regs_137_io_in; // @[RegFile.scala 66:20:@36174.4]
  wire  regs_137_io_reset; // @[RegFile.scala 66:20:@36174.4]
  wire [63:0] regs_137_io_out; // @[RegFile.scala 66:20:@36174.4]
  wire  regs_137_io_enable; // @[RegFile.scala 66:20:@36174.4]
  wire  regs_138_clock; // @[RegFile.scala 66:20:@36188.4]
  wire  regs_138_reset; // @[RegFile.scala 66:20:@36188.4]
  wire [63:0] regs_138_io_in; // @[RegFile.scala 66:20:@36188.4]
  wire  regs_138_io_reset; // @[RegFile.scala 66:20:@36188.4]
  wire [63:0] regs_138_io_out; // @[RegFile.scala 66:20:@36188.4]
  wire  regs_138_io_enable; // @[RegFile.scala 66:20:@36188.4]
  wire  regs_139_clock; // @[RegFile.scala 66:20:@36202.4]
  wire  regs_139_reset; // @[RegFile.scala 66:20:@36202.4]
  wire [63:0] regs_139_io_in; // @[RegFile.scala 66:20:@36202.4]
  wire  regs_139_io_reset; // @[RegFile.scala 66:20:@36202.4]
  wire [63:0] regs_139_io_out; // @[RegFile.scala 66:20:@36202.4]
  wire  regs_139_io_enable; // @[RegFile.scala 66:20:@36202.4]
  wire  regs_140_clock; // @[RegFile.scala 66:20:@36216.4]
  wire  regs_140_reset; // @[RegFile.scala 66:20:@36216.4]
  wire [63:0] regs_140_io_in; // @[RegFile.scala 66:20:@36216.4]
  wire  regs_140_io_reset; // @[RegFile.scala 66:20:@36216.4]
  wire [63:0] regs_140_io_out; // @[RegFile.scala 66:20:@36216.4]
  wire  regs_140_io_enable; // @[RegFile.scala 66:20:@36216.4]
  wire  regs_141_clock; // @[RegFile.scala 66:20:@36230.4]
  wire  regs_141_reset; // @[RegFile.scala 66:20:@36230.4]
  wire [63:0] regs_141_io_in; // @[RegFile.scala 66:20:@36230.4]
  wire  regs_141_io_reset; // @[RegFile.scala 66:20:@36230.4]
  wire [63:0] regs_141_io_out; // @[RegFile.scala 66:20:@36230.4]
  wire  regs_141_io_enable; // @[RegFile.scala 66:20:@36230.4]
  wire  regs_142_clock; // @[RegFile.scala 66:20:@36244.4]
  wire  regs_142_reset; // @[RegFile.scala 66:20:@36244.4]
  wire [63:0] regs_142_io_in; // @[RegFile.scala 66:20:@36244.4]
  wire  regs_142_io_reset; // @[RegFile.scala 66:20:@36244.4]
  wire [63:0] regs_142_io_out; // @[RegFile.scala 66:20:@36244.4]
  wire  regs_142_io_enable; // @[RegFile.scala 66:20:@36244.4]
  wire  regs_143_clock; // @[RegFile.scala 66:20:@36258.4]
  wire  regs_143_reset; // @[RegFile.scala 66:20:@36258.4]
  wire [63:0] regs_143_io_in; // @[RegFile.scala 66:20:@36258.4]
  wire  regs_143_io_reset; // @[RegFile.scala 66:20:@36258.4]
  wire [63:0] regs_143_io_out; // @[RegFile.scala 66:20:@36258.4]
  wire  regs_143_io_enable; // @[RegFile.scala 66:20:@36258.4]
  wire  regs_144_clock; // @[RegFile.scala 66:20:@36272.4]
  wire  regs_144_reset; // @[RegFile.scala 66:20:@36272.4]
  wire [63:0] regs_144_io_in; // @[RegFile.scala 66:20:@36272.4]
  wire  regs_144_io_reset; // @[RegFile.scala 66:20:@36272.4]
  wire [63:0] regs_144_io_out; // @[RegFile.scala 66:20:@36272.4]
  wire  regs_144_io_enable; // @[RegFile.scala 66:20:@36272.4]
  wire  regs_145_clock; // @[RegFile.scala 66:20:@36286.4]
  wire  regs_145_reset; // @[RegFile.scala 66:20:@36286.4]
  wire [63:0] regs_145_io_in; // @[RegFile.scala 66:20:@36286.4]
  wire  regs_145_io_reset; // @[RegFile.scala 66:20:@36286.4]
  wire [63:0] regs_145_io_out; // @[RegFile.scala 66:20:@36286.4]
  wire  regs_145_io_enable; // @[RegFile.scala 66:20:@36286.4]
  wire  regs_146_clock; // @[RegFile.scala 66:20:@36300.4]
  wire  regs_146_reset; // @[RegFile.scala 66:20:@36300.4]
  wire [63:0] regs_146_io_in; // @[RegFile.scala 66:20:@36300.4]
  wire  regs_146_io_reset; // @[RegFile.scala 66:20:@36300.4]
  wire [63:0] regs_146_io_out; // @[RegFile.scala 66:20:@36300.4]
  wire  regs_146_io_enable; // @[RegFile.scala 66:20:@36300.4]
  wire  regs_147_clock; // @[RegFile.scala 66:20:@36314.4]
  wire  regs_147_reset; // @[RegFile.scala 66:20:@36314.4]
  wire [63:0] regs_147_io_in; // @[RegFile.scala 66:20:@36314.4]
  wire  regs_147_io_reset; // @[RegFile.scala 66:20:@36314.4]
  wire [63:0] regs_147_io_out; // @[RegFile.scala 66:20:@36314.4]
  wire  regs_147_io_enable; // @[RegFile.scala 66:20:@36314.4]
  wire  regs_148_clock; // @[RegFile.scala 66:20:@36328.4]
  wire  regs_148_reset; // @[RegFile.scala 66:20:@36328.4]
  wire [63:0] regs_148_io_in; // @[RegFile.scala 66:20:@36328.4]
  wire  regs_148_io_reset; // @[RegFile.scala 66:20:@36328.4]
  wire [63:0] regs_148_io_out; // @[RegFile.scala 66:20:@36328.4]
  wire  regs_148_io_enable; // @[RegFile.scala 66:20:@36328.4]
  wire  regs_149_clock; // @[RegFile.scala 66:20:@36342.4]
  wire  regs_149_reset; // @[RegFile.scala 66:20:@36342.4]
  wire [63:0] regs_149_io_in; // @[RegFile.scala 66:20:@36342.4]
  wire  regs_149_io_reset; // @[RegFile.scala 66:20:@36342.4]
  wire [63:0] regs_149_io_out; // @[RegFile.scala 66:20:@36342.4]
  wire  regs_149_io_enable; // @[RegFile.scala 66:20:@36342.4]
  wire  regs_150_clock; // @[RegFile.scala 66:20:@36356.4]
  wire  regs_150_reset; // @[RegFile.scala 66:20:@36356.4]
  wire [63:0] regs_150_io_in; // @[RegFile.scala 66:20:@36356.4]
  wire  regs_150_io_reset; // @[RegFile.scala 66:20:@36356.4]
  wire [63:0] regs_150_io_out; // @[RegFile.scala 66:20:@36356.4]
  wire  regs_150_io_enable; // @[RegFile.scala 66:20:@36356.4]
  wire  regs_151_clock; // @[RegFile.scala 66:20:@36370.4]
  wire  regs_151_reset; // @[RegFile.scala 66:20:@36370.4]
  wire [63:0] regs_151_io_in; // @[RegFile.scala 66:20:@36370.4]
  wire  regs_151_io_reset; // @[RegFile.scala 66:20:@36370.4]
  wire [63:0] regs_151_io_out; // @[RegFile.scala 66:20:@36370.4]
  wire  regs_151_io_enable; // @[RegFile.scala 66:20:@36370.4]
  wire  regs_152_clock; // @[RegFile.scala 66:20:@36384.4]
  wire  regs_152_reset; // @[RegFile.scala 66:20:@36384.4]
  wire [63:0] regs_152_io_in; // @[RegFile.scala 66:20:@36384.4]
  wire  regs_152_io_reset; // @[RegFile.scala 66:20:@36384.4]
  wire [63:0] regs_152_io_out; // @[RegFile.scala 66:20:@36384.4]
  wire  regs_152_io_enable; // @[RegFile.scala 66:20:@36384.4]
  wire  regs_153_clock; // @[RegFile.scala 66:20:@36398.4]
  wire  regs_153_reset; // @[RegFile.scala 66:20:@36398.4]
  wire [63:0] regs_153_io_in; // @[RegFile.scala 66:20:@36398.4]
  wire  regs_153_io_reset; // @[RegFile.scala 66:20:@36398.4]
  wire [63:0] regs_153_io_out; // @[RegFile.scala 66:20:@36398.4]
  wire  regs_153_io_enable; // @[RegFile.scala 66:20:@36398.4]
  wire  regs_154_clock; // @[RegFile.scala 66:20:@36412.4]
  wire  regs_154_reset; // @[RegFile.scala 66:20:@36412.4]
  wire [63:0] regs_154_io_in; // @[RegFile.scala 66:20:@36412.4]
  wire  regs_154_io_reset; // @[RegFile.scala 66:20:@36412.4]
  wire [63:0] regs_154_io_out; // @[RegFile.scala 66:20:@36412.4]
  wire  regs_154_io_enable; // @[RegFile.scala 66:20:@36412.4]
  wire  regs_155_clock; // @[RegFile.scala 66:20:@36426.4]
  wire  regs_155_reset; // @[RegFile.scala 66:20:@36426.4]
  wire [63:0] regs_155_io_in; // @[RegFile.scala 66:20:@36426.4]
  wire  regs_155_io_reset; // @[RegFile.scala 66:20:@36426.4]
  wire [63:0] regs_155_io_out; // @[RegFile.scala 66:20:@36426.4]
  wire  regs_155_io_enable; // @[RegFile.scala 66:20:@36426.4]
  wire  regs_156_clock; // @[RegFile.scala 66:20:@36440.4]
  wire  regs_156_reset; // @[RegFile.scala 66:20:@36440.4]
  wire [63:0] regs_156_io_in; // @[RegFile.scala 66:20:@36440.4]
  wire  regs_156_io_reset; // @[RegFile.scala 66:20:@36440.4]
  wire [63:0] regs_156_io_out; // @[RegFile.scala 66:20:@36440.4]
  wire  regs_156_io_enable; // @[RegFile.scala 66:20:@36440.4]
  wire  regs_157_clock; // @[RegFile.scala 66:20:@36454.4]
  wire  regs_157_reset; // @[RegFile.scala 66:20:@36454.4]
  wire [63:0] regs_157_io_in; // @[RegFile.scala 66:20:@36454.4]
  wire  regs_157_io_reset; // @[RegFile.scala 66:20:@36454.4]
  wire [63:0] regs_157_io_out; // @[RegFile.scala 66:20:@36454.4]
  wire  regs_157_io_enable; // @[RegFile.scala 66:20:@36454.4]
  wire  regs_158_clock; // @[RegFile.scala 66:20:@36468.4]
  wire  regs_158_reset; // @[RegFile.scala 66:20:@36468.4]
  wire [63:0] regs_158_io_in; // @[RegFile.scala 66:20:@36468.4]
  wire  regs_158_io_reset; // @[RegFile.scala 66:20:@36468.4]
  wire [63:0] regs_158_io_out; // @[RegFile.scala 66:20:@36468.4]
  wire  regs_158_io_enable; // @[RegFile.scala 66:20:@36468.4]
  wire  regs_159_clock; // @[RegFile.scala 66:20:@36482.4]
  wire  regs_159_reset; // @[RegFile.scala 66:20:@36482.4]
  wire [63:0] regs_159_io_in; // @[RegFile.scala 66:20:@36482.4]
  wire  regs_159_io_reset; // @[RegFile.scala 66:20:@36482.4]
  wire [63:0] regs_159_io_out; // @[RegFile.scala 66:20:@36482.4]
  wire  regs_159_io_enable; // @[RegFile.scala 66:20:@36482.4]
  wire  regs_160_clock; // @[RegFile.scala 66:20:@36496.4]
  wire  regs_160_reset; // @[RegFile.scala 66:20:@36496.4]
  wire [63:0] regs_160_io_in; // @[RegFile.scala 66:20:@36496.4]
  wire  regs_160_io_reset; // @[RegFile.scala 66:20:@36496.4]
  wire [63:0] regs_160_io_out; // @[RegFile.scala 66:20:@36496.4]
  wire  regs_160_io_enable; // @[RegFile.scala 66:20:@36496.4]
  wire  regs_161_clock; // @[RegFile.scala 66:20:@36510.4]
  wire  regs_161_reset; // @[RegFile.scala 66:20:@36510.4]
  wire [63:0] regs_161_io_in; // @[RegFile.scala 66:20:@36510.4]
  wire  regs_161_io_reset; // @[RegFile.scala 66:20:@36510.4]
  wire [63:0] regs_161_io_out; // @[RegFile.scala 66:20:@36510.4]
  wire  regs_161_io_enable; // @[RegFile.scala 66:20:@36510.4]
  wire  regs_162_clock; // @[RegFile.scala 66:20:@36524.4]
  wire  regs_162_reset; // @[RegFile.scala 66:20:@36524.4]
  wire [63:0] regs_162_io_in; // @[RegFile.scala 66:20:@36524.4]
  wire  regs_162_io_reset; // @[RegFile.scala 66:20:@36524.4]
  wire [63:0] regs_162_io_out; // @[RegFile.scala 66:20:@36524.4]
  wire  regs_162_io_enable; // @[RegFile.scala 66:20:@36524.4]
  wire  regs_163_clock; // @[RegFile.scala 66:20:@36538.4]
  wire  regs_163_reset; // @[RegFile.scala 66:20:@36538.4]
  wire [63:0] regs_163_io_in; // @[RegFile.scala 66:20:@36538.4]
  wire  regs_163_io_reset; // @[RegFile.scala 66:20:@36538.4]
  wire [63:0] regs_163_io_out; // @[RegFile.scala 66:20:@36538.4]
  wire  regs_163_io_enable; // @[RegFile.scala 66:20:@36538.4]
  wire  regs_164_clock; // @[RegFile.scala 66:20:@36552.4]
  wire  regs_164_reset; // @[RegFile.scala 66:20:@36552.4]
  wire [63:0] regs_164_io_in; // @[RegFile.scala 66:20:@36552.4]
  wire  regs_164_io_reset; // @[RegFile.scala 66:20:@36552.4]
  wire [63:0] regs_164_io_out; // @[RegFile.scala 66:20:@36552.4]
  wire  regs_164_io_enable; // @[RegFile.scala 66:20:@36552.4]
  wire  regs_165_clock; // @[RegFile.scala 66:20:@36566.4]
  wire  regs_165_reset; // @[RegFile.scala 66:20:@36566.4]
  wire [63:0] regs_165_io_in; // @[RegFile.scala 66:20:@36566.4]
  wire  regs_165_io_reset; // @[RegFile.scala 66:20:@36566.4]
  wire [63:0] regs_165_io_out; // @[RegFile.scala 66:20:@36566.4]
  wire  regs_165_io_enable; // @[RegFile.scala 66:20:@36566.4]
  wire  regs_166_clock; // @[RegFile.scala 66:20:@36580.4]
  wire  regs_166_reset; // @[RegFile.scala 66:20:@36580.4]
  wire [63:0] regs_166_io_in; // @[RegFile.scala 66:20:@36580.4]
  wire  regs_166_io_reset; // @[RegFile.scala 66:20:@36580.4]
  wire [63:0] regs_166_io_out; // @[RegFile.scala 66:20:@36580.4]
  wire  regs_166_io_enable; // @[RegFile.scala 66:20:@36580.4]
  wire  regs_167_clock; // @[RegFile.scala 66:20:@36594.4]
  wire  regs_167_reset; // @[RegFile.scala 66:20:@36594.4]
  wire [63:0] regs_167_io_in; // @[RegFile.scala 66:20:@36594.4]
  wire  regs_167_io_reset; // @[RegFile.scala 66:20:@36594.4]
  wire [63:0] regs_167_io_out; // @[RegFile.scala 66:20:@36594.4]
  wire  regs_167_io_enable; // @[RegFile.scala 66:20:@36594.4]
  wire  regs_168_clock; // @[RegFile.scala 66:20:@36608.4]
  wire  regs_168_reset; // @[RegFile.scala 66:20:@36608.4]
  wire [63:0] regs_168_io_in; // @[RegFile.scala 66:20:@36608.4]
  wire  regs_168_io_reset; // @[RegFile.scala 66:20:@36608.4]
  wire [63:0] regs_168_io_out; // @[RegFile.scala 66:20:@36608.4]
  wire  regs_168_io_enable; // @[RegFile.scala 66:20:@36608.4]
  wire  regs_169_clock; // @[RegFile.scala 66:20:@36622.4]
  wire  regs_169_reset; // @[RegFile.scala 66:20:@36622.4]
  wire [63:0] regs_169_io_in; // @[RegFile.scala 66:20:@36622.4]
  wire  regs_169_io_reset; // @[RegFile.scala 66:20:@36622.4]
  wire [63:0] regs_169_io_out; // @[RegFile.scala 66:20:@36622.4]
  wire  regs_169_io_enable; // @[RegFile.scala 66:20:@36622.4]
  wire  regs_170_clock; // @[RegFile.scala 66:20:@36636.4]
  wire  regs_170_reset; // @[RegFile.scala 66:20:@36636.4]
  wire [63:0] regs_170_io_in; // @[RegFile.scala 66:20:@36636.4]
  wire  regs_170_io_reset; // @[RegFile.scala 66:20:@36636.4]
  wire [63:0] regs_170_io_out; // @[RegFile.scala 66:20:@36636.4]
  wire  regs_170_io_enable; // @[RegFile.scala 66:20:@36636.4]
  wire  regs_171_clock; // @[RegFile.scala 66:20:@36650.4]
  wire  regs_171_reset; // @[RegFile.scala 66:20:@36650.4]
  wire [63:0] regs_171_io_in; // @[RegFile.scala 66:20:@36650.4]
  wire  regs_171_io_reset; // @[RegFile.scala 66:20:@36650.4]
  wire [63:0] regs_171_io_out; // @[RegFile.scala 66:20:@36650.4]
  wire  regs_171_io_enable; // @[RegFile.scala 66:20:@36650.4]
  wire  regs_172_clock; // @[RegFile.scala 66:20:@36664.4]
  wire  regs_172_reset; // @[RegFile.scala 66:20:@36664.4]
  wire [63:0] regs_172_io_in; // @[RegFile.scala 66:20:@36664.4]
  wire  regs_172_io_reset; // @[RegFile.scala 66:20:@36664.4]
  wire [63:0] regs_172_io_out; // @[RegFile.scala 66:20:@36664.4]
  wire  regs_172_io_enable; // @[RegFile.scala 66:20:@36664.4]
  wire  regs_173_clock; // @[RegFile.scala 66:20:@36678.4]
  wire  regs_173_reset; // @[RegFile.scala 66:20:@36678.4]
  wire [63:0] regs_173_io_in; // @[RegFile.scala 66:20:@36678.4]
  wire  regs_173_io_reset; // @[RegFile.scala 66:20:@36678.4]
  wire [63:0] regs_173_io_out; // @[RegFile.scala 66:20:@36678.4]
  wire  regs_173_io_enable; // @[RegFile.scala 66:20:@36678.4]
  wire  regs_174_clock; // @[RegFile.scala 66:20:@36692.4]
  wire  regs_174_reset; // @[RegFile.scala 66:20:@36692.4]
  wire [63:0] regs_174_io_in; // @[RegFile.scala 66:20:@36692.4]
  wire  regs_174_io_reset; // @[RegFile.scala 66:20:@36692.4]
  wire [63:0] regs_174_io_out; // @[RegFile.scala 66:20:@36692.4]
  wire  regs_174_io_enable; // @[RegFile.scala 66:20:@36692.4]
  wire  regs_175_clock; // @[RegFile.scala 66:20:@36706.4]
  wire  regs_175_reset; // @[RegFile.scala 66:20:@36706.4]
  wire [63:0] regs_175_io_in; // @[RegFile.scala 66:20:@36706.4]
  wire  regs_175_io_reset; // @[RegFile.scala 66:20:@36706.4]
  wire [63:0] regs_175_io_out; // @[RegFile.scala 66:20:@36706.4]
  wire  regs_175_io_enable; // @[RegFile.scala 66:20:@36706.4]
  wire  regs_176_clock; // @[RegFile.scala 66:20:@36720.4]
  wire  regs_176_reset; // @[RegFile.scala 66:20:@36720.4]
  wire [63:0] regs_176_io_in; // @[RegFile.scala 66:20:@36720.4]
  wire  regs_176_io_reset; // @[RegFile.scala 66:20:@36720.4]
  wire [63:0] regs_176_io_out; // @[RegFile.scala 66:20:@36720.4]
  wire  regs_176_io_enable; // @[RegFile.scala 66:20:@36720.4]
  wire  regs_177_clock; // @[RegFile.scala 66:20:@36734.4]
  wire  regs_177_reset; // @[RegFile.scala 66:20:@36734.4]
  wire [63:0] regs_177_io_in; // @[RegFile.scala 66:20:@36734.4]
  wire  regs_177_io_reset; // @[RegFile.scala 66:20:@36734.4]
  wire [63:0] regs_177_io_out; // @[RegFile.scala 66:20:@36734.4]
  wire  regs_177_io_enable; // @[RegFile.scala 66:20:@36734.4]
  wire  regs_178_clock; // @[RegFile.scala 66:20:@36748.4]
  wire  regs_178_reset; // @[RegFile.scala 66:20:@36748.4]
  wire [63:0] regs_178_io_in; // @[RegFile.scala 66:20:@36748.4]
  wire  regs_178_io_reset; // @[RegFile.scala 66:20:@36748.4]
  wire [63:0] regs_178_io_out; // @[RegFile.scala 66:20:@36748.4]
  wire  regs_178_io_enable; // @[RegFile.scala 66:20:@36748.4]
  wire  regs_179_clock; // @[RegFile.scala 66:20:@36762.4]
  wire  regs_179_reset; // @[RegFile.scala 66:20:@36762.4]
  wire [63:0] regs_179_io_in; // @[RegFile.scala 66:20:@36762.4]
  wire  regs_179_io_reset; // @[RegFile.scala 66:20:@36762.4]
  wire [63:0] regs_179_io_out; // @[RegFile.scala 66:20:@36762.4]
  wire  regs_179_io_enable; // @[RegFile.scala 66:20:@36762.4]
  wire  regs_180_clock; // @[RegFile.scala 66:20:@36776.4]
  wire  regs_180_reset; // @[RegFile.scala 66:20:@36776.4]
  wire [63:0] regs_180_io_in; // @[RegFile.scala 66:20:@36776.4]
  wire  regs_180_io_reset; // @[RegFile.scala 66:20:@36776.4]
  wire [63:0] regs_180_io_out; // @[RegFile.scala 66:20:@36776.4]
  wire  regs_180_io_enable; // @[RegFile.scala 66:20:@36776.4]
  wire  regs_181_clock; // @[RegFile.scala 66:20:@36790.4]
  wire  regs_181_reset; // @[RegFile.scala 66:20:@36790.4]
  wire [63:0] regs_181_io_in; // @[RegFile.scala 66:20:@36790.4]
  wire  regs_181_io_reset; // @[RegFile.scala 66:20:@36790.4]
  wire [63:0] regs_181_io_out; // @[RegFile.scala 66:20:@36790.4]
  wire  regs_181_io_enable; // @[RegFile.scala 66:20:@36790.4]
  wire  regs_182_clock; // @[RegFile.scala 66:20:@36804.4]
  wire  regs_182_reset; // @[RegFile.scala 66:20:@36804.4]
  wire [63:0] regs_182_io_in; // @[RegFile.scala 66:20:@36804.4]
  wire  regs_182_io_reset; // @[RegFile.scala 66:20:@36804.4]
  wire [63:0] regs_182_io_out; // @[RegFile.scala 66:20:@36804.4]
  wire  regs_182_io_enable; // @[RegFile.scala 66:20:@36804.4]
  wire  regs_183_clock; // @[RegFile.scala 66:20:@36818.4]
  wire  regs_183_reset; // @[RegFile.scala 66:20:@36818.4]
  wire [63:0] regs_183_io_in; // @[RegFile.scala 66:20:@36818.4]
  wire  regs_183_io_reset; // @[RegFile.scala 66:20:@36818.4]
  wire [63:0] regs_183_io_out; // @[RegFile.scala 66:20:@36818.4]
  wire  regs_183_io_enable; // @[RegFile.scala 66:20:@36818.4]
  wire  regs_184_clock; // @[RegFile.scala 66:20:@36832.4]
  wire  regs_184_reset; // @[RegFile.scala 66:20:@36832.4]
  wire [63:0] regs_184_io_in; // @[RegFile.scala 66:20:@36832.4]
  wire  regs_184_io_reset; // @[RegFile.scala 66:20:@36832.4]
  wire [63:0] regs_184_io_out; // @[RegFile.scala 66:20:@36832.4]
  wire  regs_184_io_enable; // @[RegFile.scala 66:20:@36832.4]
  wire  regs_185_clock; // @[RegFile.scala 66:20:@36846.4]
  wire  regs_185_reset; // @[RegFile.scala 66:20:@36846.4]
  wire [63:0] regs_185_io_in; // @[RegFile.scala 66:20:@36846.4]
  wire  regs_185_io_reset; // @[RegFile.scala 66:20:@36846.4]
  wire [63:0] regs_185_io_out; // @[RegFile.scala 66:20:@36846.4]
  wire  regs_185_io_enable; // @[RegFile.scala 66:20:@36846.4]
  wire  regs_186_clock; // @[RegFile.scala 66:20:@36860.4]
  wire  regs_186_reset; // @[RegFile.scala 66:20:@36860.4]
  wire [63:0] regs_186_io_in; // @[RegFile.scala 66:20:@36860.4]
  wire  regs_186_io_reset; // @[RegFile.scala 66:20:@36860.4]
  wire [63:0] regs_186_io_out; // @[RegFile.scala 66:20:@36860.4]
  wire  regs_186_io_enable; // @[RegFile.scala 66:20:@36860.4]
  wire  regs_187_clock; // @[RegFile.scala 66:20:@36874.4]
  wire  regs_187_reset; // @[RegFile.scala 66:20:@36874.4]
  wire [63:0] regs_187_io_in; // @[RegFile.scala 66:20:@36874.4]
  wire  regs_187_io_reset; // @[RegFile.scala 66:20:@36874.4]
  wire [63:0] regs_187_io_out; // @[RegFile.scala 66:20:@36874.4]
  wire  regs_187_io_enable; // @[RegFile.scala 66:20:@36874.4]
  wire  regs_188_clock; // @[RegFile.scala 66:20:@36888.4]
  wire  regs_188_reset; // @[RegFile.scala 66:20:@36888.4]
  wire [63:0] regs_188_io_in; // @[RegFile.scala 66:20:@36888.4]
  wire  regs_188_io_reset; // @[RegFile.scala 66:20:@36888.4]
  wire [63:0] regs_188_io_out; // @[RegFile.scala 66:20:@36888.4]
  wire  regs_188_io_enable; // @[RegFile.scala 66:20:@36888.4]
  wire  regs_189_clock; // @[RegFile.scala 66:20:@36902.4]
  wire  regs_189_reset; // @[RegFile.scala 66:20:@36902.4]
  wire [63:0] regs_189_io_in; // @[RegFile.scala 66:20:@36902.4]
  wire  regs_189_io_reset; // @[RegFile.scala 66:20:@36902.4]
  wire [63:0] regs_189_io_out; // @[RegFile.scala 66:20:@36902.4]
  wire  regs_189_io_enable; // @[RegFile.scala 66:20:@36902.4]
  wire  regs_190_clock; // @[RegFile.scala 66:20:@36916.4]
  wire  regs_190_reset; // @[RegFile.scala 66:20:@36916.4]
  wire [63:0] regs_190_io_in; // @[RegFile.scala 66:20:@36916.4]
  wire  regs_190_io_reset; // @[RegFile.scala 66:20:@36916.4]
  wire [63:0] regs_190_io_out; // @[RegFile.scala 66:20:@36916.4]
  wire  regs_190_io_enable; // @[RegFile.scala 66:20:@36916.4]
  wire  regs_191_clock; // @[RegFile.scala 66:20:@36930.4]
  wire  regs_191_reset; // @[RegFile.scala 66:20:@36930.4]
  wire [63:0] regs_191_io_in; // @[RegFile.scala 66:20:@36930.4]
  wire  regs_191_io_reset; // @[RegFile.scala 66:20:@36930.4]
  wire [63:0] regs_191_io_out; // @[RegFile.scala 66:20:@36930.4]
  wire  regs_191_io_enable; // @[RegFile.scala 66:20:@36930.4]
  wire  regs_192_clock; // @[RegFile.scala 66:20:@36944.4]
  wire  regs_192_reset; // @[RegFile.scala 66:20:@36944.4]
  wire [63:0] regs_192_io_in; // @[RegFile.scala 66:20:@36944.4]
  wire  regs_192_io_reset; // @[RegFile.scala 66:20:@36944.4]
  wire [63:0] regs_192_io_out; // @[RegFile.scala 66:20:@36944.4]
  wire  regs_192_io_enable; // @[RegFile.scala 66:20:@36944.4]
  wire  regs_193_clock; // @[RegFile.scala 66:20:@36958.4]
  wire  regs_193_reset; // @[RegFile.scala 66:20:@36958.4]
  wire [63:0] regs_193_io_in; // @[RegFile.scala 66:20:@36958.4]
  wire  regs_193_io_reset; // @[RegFile.scala 66:20:@36958.4]
  wire [63:0] regs_193_io_out; // @[RegFile.scala 66:20:@36958.4]
  wire  regs_193_io_enable; // @[RegFile.scala 66:20:@36958.4]
  wire  regs_194_clock; // @[RegFile.scala 66:20:@36972.4]
  wire  regs_194_reset; // @[RegFile.scala 66:20:@36972.4]
  wire [63:0] regs_194_io_in; // @[RegFile.scala 66:20:@36972.4]
  wire  regs_194_io_reset; // @[RegFile.scala 66:20:@36972.4]
  wire [63:0] regs_194_io_out; // @[RegFile.scala 66:20:@36972.4]
  wire  regs_194_io_enable; // @[RegFile.scala 66:20:@36972.4]
  wire  regs_195_clock; // @[RegFile.scala 66:20:@36986.4]
  wire  regs_195_reset; // @[RegFile.scala 66:20:@36986.4]
  wire [63:0] regs_195_io_in; // @[RegFile.scala 66:20:@36986.4]
  wire  regs_195_io_reset; // @[RegFile.scala 66:20:@36986.4]
  wire [63:0] regs_195_io_out; // @[RegFile.scala 66:20:@36986.4]
  wire  regs_195_io_enable; // @[RegFile.scala 66:20:@36986.4]
  wire  regs_196_clock; // @[RegFile.scala 66:20:@37000.4]
  wire  regs_196_reset; // @[RegFile.scala 66:20:@37000.4]
  wire [63:0] regs_196_io_in; // @[RegFile.scala 66:20:@37000.4]
  wire  regs_196_io_reset; // @[RegFile.scala 66:20:@37000.4]
  wire [63:0] regs_196_io_out; // @[RegFile.scala 66:20:@37000.4]
  wire  regs_196_io_enable; // @[RegFile.scala 66:20:@37000.4]
  wire  regs_197_clock; // @[RegFile.scala 66:20:@37014.4]
  wire  regs_197_reset; // @[RegFile.scala 66:20:@37014.4]
  wire [63:0] regs_197_io_in; // @[RegFile.scala 66:20:@37014.4]
  wire  regs_197_io_reset; // @[RegFile.scala 66:20:@37014.4]
  wire [63:0] regs_197_io_out; // @[RegFile.scala 66:20:@37014.4]
  wire  regs_197_io_enable; // @[RegFile.scala 66:20:@37014.4]
  wire  regs_198_clock; // @[RegFile.scala 66:20:@37028.4]
  wire  regs_198_reset; // @[RegFile.scala 66:20:@37028.4]
  wire [63:0] regs_198_io_in; // @[RegFile.scala 66:20:@37028.4]
  wire  regs_198_io_reset; // @[RegFile.scala 66:20:@37028.4]
  wire [63:0] regs_198_io_out; // @[RegFile.scala 66:20:@37028.4]
  wire  regs_198_io_enable; // @[RegFile.scala 66:20:@37028.4]
  wire  regs_199_clock; // @[RegFile.scala 66:20:@37042.4]
  wire  regs_199_reset; // @[RegFile.scala 66:20:@37042.4]
  wire [63:0] regs_199_io_in; // @[RegFile.scala 66:20:@37042.4]
  wire  regs_199_io_reset; // @[RegFile.scala 66:20:@37042.4]
  wire [63:0] regs_199_io_out; // @[RegFile.scala 66:20:@37042.4]
  wire  regs_199_io_enable; // @[RegFile.scala 66:20:@37042.4]
  wire  regs_200_clock; // @[RegFile.scala 66:20:@37056.4]
  wire  regs_200_reset; // @[RegFile.scala 66:20:@37056.4]
  wire [63:0] regs_200_io_in; // @[RegFile.scala 66:20:@37056.4]
  wire  regs_200_io_reset; // @[RegFile.scala 66:20:@37056.4]
  wire [63:0] regs_200_io_out; // @[RegFile.scala 66:20:@37056.4]
  wire  regs_200_io_enable; // @[RegFile.scala 66:20:@37056.4]
  wire  regs_201_clock; // @[RegFile.scala 66:20:@37070.4]
  wire  regs_201_reset; // @[RegFile.scala 66:20:@37070.4]
  wire [63:0] regs_201_io_in; // @[RegFile.scala 66:20:@37070.4]
  wire  regs_201_io_reset; // @[RegFile.scala 66:20:@37070.4]
  wire [63:0] regs_201_io_out; // @[RegFile.scala 66:20:@37070.4]
  wire  regs_201_io_enable; // @[RegFile.scala 66:20:@37070.4]
  wire  regs_202_clock; // @[RegFile.scala 66:20:@37084.4]
  wire  regs_202_reset; // @[RegFile.scala 66:20:@37084.4]
  wire [63:0] regs_202_io_in; // @[RegFile.scala 66:20:@37084.4]
  wire  regs_202_io_reset; // @[RegFile.scala 66:20:@37084.4]
  wire [63:0] regs_202_io_out; // @[RegFile.scala 66:20:@37084.4]
  wire  regs_202_io_enable; // @[RegFile.scala 66:20:@37084.4]
  wire  regs_203_clock; // @[RegFile.scala 66:20:@37098.4]
  wire  regs_203_reset; // @[RegFile.scala 66:20:@37098.4]
  wire [63:0] regs_203_io_in; // @[RegFile.scala 66:20:@37098.4]
  wire  regs_203_io_reset; // @[RegFile.scala 66:20:@37098.4]
  wire [63:0] regs_203_io_out; // @[RegFile.scala 66:20:@37098.4]
  wire  regs_203_io_enable; // @[RegFile.scala 66:20:@37098.4]
  wire  regs_204_clock; // @[RegFile.scala 66:20:@37112.4]
  wire  regs_204_reset; // @[RegFile.scala 66:20:@37112.4]
  wire [63:0] regs_204_io_in; // @[RegFile.scala 66:20:@37112.4]
  wire  regs_204_io_reset; // @[RegFile.scala 66:20:@37112.4]
  wire [63:0] regs_204_io_out; // @[RegFile.scala 66:20:@37112.4]
  wire  regs_204_io_enable; // @[RegFile.scala 66:20:@37112.4]
  wire  regs_205_clock; // @[RegFile.scala 66:20:@37126.4]
  wire  regs_205_reset; // @[RegFile.scala 66:20:@37126.4]
  wire [63:0] regs_205_io_in; // @[RegFile.scala 66:20:@37126.4]
  wire  regs_205_io_reset; // @[RegFile.scala 66:20:@37126.4]
  wire [63:0] regs_205_io_out; // @[RegFile.scala 66:20:@37126.4]
  wire  regs_205_io_enable; // @[RegFile.scala 66:20:@37126.4]
  wire  regs_206_clock; // @[RegFile.scala 66:20:@37140.4]
  wire  regs_206_reset; // @[RegFile.scala 66:20:@37140.4]
  wire [63:0] regs_206_io_in; // @[RegFile.scala 66:20:@37140.4]
  wire  regs_206_io_reset; // @[RegFile.scala 66:20:@37140.4]
  wire [63:0] regs_206_io_out; // @[RegFile.scala 66:20:@37140.4]
  wire  regs_206_io_enable; // @[RegFile.scala 66:20:@37140.4]
  wire  regs_207_clock; // @[RegFile.scala 66:20:@37154.4]
  wire  regs_207_reset; // @[RegFile.scala 66:20:@37154.4]
  wire [63:0] regs_207_io_in; // @[RegFile.scala 66:20:@37154.4]
  wire  regs_207_io_reset; // @[RegFile.scala 66:20:@37154.4]
  wire [63:0] regs_207_io_out; // @[RegFile.scala 66:20:@37154.4]
  wire  regs_207_io_enable; // @[RegFile.scala 66:20:@37154.4]
  wire  regs_208_clock; // @[RegFile.scala 66:20:@37168.4]
  wire  regs_208_reset; // @[RegFile.scala 66:20:@37168.4]
  wire [63:0] regs_208_io_in; // @[RegFile.scala 66:20:@37168.4]
  wire  regs_208_io_reset; // @[RegFile.scala 66:20:@37168.4]
  wire [63:0] regs_208_io_out; // @[RegFile.scala 66:20:@37168.4]
  wire  regs_208_io_enable; // @[RegFile.scala 66:20:@37168.4]
  wire  regs_209_clock; // @[RegFile.scala 66:20:@37182.4]
  wire  regs_209_reset; // @[RegFile.scala 66:20:@37182.4]
  wire [63:0] regs_209_io_in; // @[RegFile.scala 66:20:@37182.4]
  wire  regs_209_io_reset; // @[RegFile.scala 66:20:@37182.4]
  wire [63:0] regs_209_io_out; // @[RegFile.scala 66:20:@37182.4]
  wire  regs_209_io_enable; // @[RegFile.scala 66:20:@37182.4]
  wire  regs_210_clock; // @[RegFile.scala 66:20:@37196.4]
  wire  regs_210_reset; // @[RegFile.scala 66:20:@37196.4]
  wire [63:0] regs_210_io_in; // @[RegFile.scala 66:20:@37196.4]
  wire  regs_210_io_reset; // @[RegFile.scala 66:20:@37196.4]
  wire [63:0] regs_210_io_out; // @[RegFile.scala 66:20:@37196.4]
  wire  regs_210_io_enable; // @[RegFile.scala 66:20:@37196.4]
  wire  regs_211_clock; // @[RegFile.scala 66:20:@37210.4]
  wire  regs_211_reset; // @[RegFile.scala 66:20:@37210.4]
  wire [63:0] regs_211_io_in; // @[RegFile.scala 66:20:@37210.4]
  wire  regs_211_io_reset; // @[RegFile.scala 66:20:@37210.4]
  wire [63:0] regs_211_io_out; // @[RegFile.scala 66:20:@37210.4]
  wire  regs_211_io_enable; // @[RegFile.scala 66:20:@37210.4]
  wire  regs_212_clock; // @[RegFile.scala 66:20:@37224.4]
  wire  regs_212_reset; // @[RegFile.scala 66:20:@37224.4]
  wire [63:0] regs_212_io_in; // @[RegFile.scala 66:20:@37224.4]
  wire  regs_212_io_reset; // @[RegFile.scala 66:20:@37224.4]
  wire [63:0] regs_212_io_out; // @[RegFile.scala 66:20:@37224.4]
  wire  regs_212_io_enable; // @[RegFile.scala 66:20:@37224.4]
  wire  regs_213_clock; // @[RegFile.scala 66:20:@37238.4]
  wire  regs_213_reset; // @[RegFile.scala 66:20:@37238.4]
  wire [63:0] regs_213_io_in; // @[RegFile.scala 66:20:@37238.4]
  wire  regs_213_io_reset; // @[RegFile.scala 66:20:@37238.4]
  wire [63:0] regs_213_io_out; // @[RegFile.scala 66:20:@37238.4]
  wire  regs_213_io_enable; // @[RegFile.scala 66:20:@37238.4]
  wire  regs_214_clock; // @[RegFile.scala 66:20:@37252.4]
  wire  regs_214_reset; // @[RegFile.scala 66:20:@37252.4]
  wire [63:0] regs_214_io_in; // @[RegFile.scala 66:20:@37252.4]
  wire  regs_214_io_reset; // @[RegFile.scala 66:20:@37252.4]
  wire [63:0] regs_214_io_out; // @[RegFile.scala 66:20:@37252.4]
  wire  regs_214_io_enable; // @[RegFile.scala 66:20:@37252.4]
  wire  regs_215_clock; // @[RegFile.scala 66:20:@37266.4]
  wire  regs_215_reset; // @[RegFile.scala 66:20:@37266.4]
  wire [63:0] regs_215_io_in; // @[RegFile.scala 66:20:@37266.4]
  wire  regs_215_io_reset; // @[RegFile.scala 66:20:@37266.4]
  wire [63:0] regs_215_io_out; // @[RegFile.scala 66:20:@37266.4]
  wire  regs_215_io_enable; // @[RegFile.scala 66:20:@37266.4]
  wire  regs_216_clock; // @[RegFile.scala 66:20:@37280.4]
  wire  regs_216_reset; // @[RegFile.scala 66:20:@37280.4]
  wire [63:0] regs_216_io_in; // @[RegFile.scala 66:20:@37280.4]
  wire  regs_216_io_reset; // @[RegFile.scala 66:20:@37280.4]
  wire [63:0] regs_216_io_out; // @[RegFile.scala 66:20:@37280.4]
  wire  regs_216_io_enable; // @[RegFile.scala 66:20:@37280.4]
  wire  regs_217_clock; // @[RegFile.scala 66:20:@37294.4]
  wire  regs_217_reset; // @[RegFile.scala 66:20:@37294.4]
  wire [63:0] regs_217_io_in; // @[RegFile.scala 66:20:@37294.4]
  wire  regs_217_io_reset; // @[RegFile.scala 66:20:@37294.4]
  wire [63:0] regs_217_io_out; // @[RegFile.scala 66:20:@37294.4]
  wire  regs_217_io_enable; // @[RegFile.scala 66:20:@37294.4]
  wire  regs_218_clock; // @[RegFile.scala 66:20:@37308.4]
  wire  regs_218_reset; // @[RegFile.scala 66:20:@37308.4]
  wire [63:0] regs_218_io_in; // @[RegFile.scala 66:20:@37308.4]
  wire  regs_218_io_reset; // @[RegFile.scala 66:20:@37308.4]
  wire [63:0] regs_218_io_out; // @[RegFile.scala 66:20:@37308.4]
  wire  regs_218_io_enable; // @[RegFile.scala 66:20:@37308.4]
  wire  regs_219_clock; // @[RegFile.scala 66:20:@37322.4]
  wire  regs_219_reset; // @[RegFile.scala 66:20:@37322.4]
  wire [63:0] regs_219_io_in; // @[RegFile.scala 66:20:@37322.4]
  wire  regs_219_io_reset; // @[RegFile.scala 66:20:@37322.4]
  wire [63:0] regs_219_io_out; // @[RegFile.scala 66:20:@37322.4]
  wire  regs_219_io_enable; // @[RegFile.scala 66:20:@37322.4]
  wire  regs_220_clock; // @[RegFile.scala 66:20:@37336.4]
  wire  regs_220_reset; // @[RegFile.scala 66:20:@37336.4]
  wire [63:0] regs_220_io_in; // @[RegFile.scala 66:20:@37336.4]
  wire  regs_220_io_reset; // @[RegFile.scala 66:20:@37336.4]
  wire [63:0] regs_220_io_out; // @[RegFile.scala 66:20:@37336.4]
  wire  regs_220_io_enable; // @[RegFile.scala 66:20:@37336.4]
  wire  regs_221_clock; // @[RegFile.scala 66:20:@37350.4]
  wire  regs_221_reset; // @[RegFile.scala 66:20:@37350.4]
  wire [63:0] regs_221_io_in; // @[RegFile.scala 66:20:@37350.4]
  wire  regs_221_io_reset; // @[RegFile.scala 66:20:@37350.4]
  wire [63:0] regs_221_io_out; // @[RegFile.scala 66:20:@37350.4]
  wire  regs_221_io_enable; // @[RegFile.scala 66:20:@37350.4]
  wire  regs_222_clock; // @[RegFile.scala 66:20:@37364.4]
  wire  regs_222_reset; // @[RegFile.scala 66:20:@37364.4]
  wire [63:0] regs_222_io_in; // @[RegFile.scala 66:20:@37364.4]
  wire  regs_222_io_reset; // @[RegFile.scala 66:20:@37364.4]
  wire [63:0] regs_222_io_out; // @[RegFile.scala 66:20:@37364.4]
  wire  regs_222_io_enable; // @[RegFile.scala 66:20:@37364.4]
  wire  regs_223_clock; // @[RegFile.scala 66:20:@37378.4]
  wire  regs_223_reset; // @[RegFile.scala 66:20:@37378.4]
  wire [63:0] regs_223_io_in; // @[RegFile.scala 66:20:@37378.4]
  wire  regs_223_io_reset; // @[RegFile.scala 66:20:@37378.4]
  wire [63:0] regs_223_io_out; // @[RegFile.scala 66:20:@37378.4]
  wire  regs_223_io_enable; // @[RegFile.scala 66:20:@37378.4]
  wire  regs_224_clock; // @[RegFile.scala 66:20:@37392.4]
  wire  regs_224_reset; // @[RegFile.scala 66:20:@37392.4]
  wire [63:0] regs_224_io_in; // @[RegFile.scala 66:20:@37392.4]
  wire  regs_224_io_reset; // @[RegFile.scala 66:20:@37392.4]
  wire [63:0] regs_224_io_out; // @[RegFile.scala 66:20:@37392.4]
  wire  regs_224_io_enable; // @[RegFile.scala 66:20:@37392.4]
  wire  regs_225_clock; // @[RegFile.scala 66:20:@37406.4]
  wire  regs_225_reset; // @[RegFile.scala 66:20:@37406.4]
  wire [63:0] regs_225_io_in; // @[RegFile.scala 66:20:@37406.4]
  wire  regs_225_io_reset; // @[RegFile.scala 66:20:@37406.4]
  wire [63:0] regs_225_io_out; // @[RegFile.scala 66:20:@37406.4]
  wire  regs_225_io_enable; // @[RegFile.scala 66:20:@37406.4]
  wire  regs_226_clock; // @[RegFile.scala 66:20:@37420.4]
  wire  regs_226_reset; // @[RegFile.scala 66:20:@37420.4]
  wire [63:0] regs_226_io_in; // @[RegFile.scala 66:20:@37420.4]
  wire  regs_226_io_reset; // @[RegFile.scala 66:20:@37420.4]
  wire [63:0] regs_226_io_out; // @[RegFile.scala 66:20:@37420.4]
  wire  regs_226_io_enable; // @[RegFile.scala 66:20:@37420.4]
  wire  regs_227_clock; // @[RegFile.scala 66:20:@37434.4]
  wire  regs_227_reset; // @[RegFile.scala 66:20:@37434.4]
  wire [63:0] regs_227_io_in; // @[RegFile.scala 66:20:@37434.4]
  wire  regs_227_io_reset; // @[RegFile.scala 66:20:@37434.4]
  wire [63:0] regs_227_io_out; // @[RegFile.scala 66:20:@37434.4]
  wire  regs_227_io_enable; // @[RegFile.scala 66:20:@37434.4]
  wire  regs_228_clock; // @[RegFile.scala 66:20:@37448.4]
  wire  regs_228_reset; // @[RegFile.scala 66:20:@37448.4]
  wire [63:0] regs_228_io_in; // @[RegFile.scala 66:20:@37448.4]
  wire  regs_228_io_reset; // @[RegFile.scala 66:20:@37448.4]
  wire [63:0] regs_228_io_out; // @[RegFile.scala 66:20:@37448.4]
  wire  regs_228_io_enable; // @[RegFile.scala 66:20:@37448.4]
  wire  regs_229_clock; // @[RegFile.scala 66:20:@37462.4]
  wire  regs_229_reset; // @[RegFile.scala 66:20:@37462.4]
  wire [63:0] regs_229_io_in; // @[RegFile.scala 66:20:@37462.4]
  wire  regs_229_io_reset; // @[RegFile.scala 66:20:@37462.4]
  wire [63:0] regs_229_io_out; // @[RegFile.scala 66:20:@37462.4]
  wire  regs_229_io_enable; // @[RegFile.scala 66:20:@37462.4]
  wire  regs_230_clock; // @[RegFile.scala 66:20:@37476.4]
  wire  regs_230_reset; // @[RegFile.scala 66:20:@37476.4]
  wire [63:0] regs_230_io_in; // @[RegFile.scala 66:20:@37476.4]
  wire  regs_230_io_reset; // @[RegFile.scala 66:20:@37476.4]
  wire [63:0] regs_230_io_out; // @[RegFile.scala 66:20:@37476.4]
  wire  regs_230_io_enable; // @[RegFile.scala 66:20:@37476.4]
  wire  regs_231_clock; // @[RegFile.scala 66:20:@37490.4]
  wire  regs_231_reset; // @[RegFile.scala 66:20:@37490.4]
  wire [63:0] regs_231_io_in; // @[RegFile.scala 66:20:@37490.4]
  wire  regs_231_io_reset; // @[RegFile.scala 66:20:@37490.4]
  wire [63:0] regs_231_io_out; // @[RegFile.scala 66:20:@37490.4]
  wire  regs_231_io_enable; // @[RegFile.scala 66:20:@37490.4]
  wire  regs_232_clock; // @[RegFile.scala 66:20:@37504.4]
  wire  regs_232_reset; // @[RegFile.scala 66:20:@37504.4]
  wire [63:0] regs_232_io_in; // @[RegFile.scala 66:20:@37504.4]
  wire  regs_232_io_reset; // @[RegFile.scala 66:20:@37504.4]
  wire [63:0] regs_232_io_out; // @[RegFile.scala 66:20:@37504.4]
  wire  regs_232_io_enable; // @[RegFile.scala 66:20:@37504.4]
  wire  regs_233_clock; // @[RegFile.scala 66:20:@37518.4]
  wire  regs_233_reset; // @[RegFile.scala 66:20:@37518.4]
  wire [63:0] regs_233_io_in; // @[RegFile.scala 66:20:@37518.4]
  wire  regs_233_io_reset; // @[RegFile.scala 66:20:@37518.4]
  wire [63:0] regs_233_io_out; // @[RegFile.scala 66:20:@37518.4]
  wire  regs_233_io_enable; // @[RegFile.scala 66:20:@37518.4]
  wire  regs_234_clock; // @[RegFile.scala 66:20:@37532.4]
  wire  regs_234_reset; // @[RegFile.scala 66:20:@37532.4]
  wire [63:0] regs_234_io_in; // @[RegFile.scala 66:20:@37532.4]
  wire  regs_234_io_reset; // @[RegFile.scala 66:20:@37532.4]
  wire [63:0] regs_234_io_out; // @[RegFile.scala 66:20:@37532.4]
  wire  regs_234_io_enable; // @[RegFile.scala 66:20:@37532.4]
  wire  regs_235_clock; // @[RegFile.scala 66:20:@37546.4]
  wire  regs_235_reset; // @[RegFile.scala 66:20:@37546.4]
  wire [63:0] regs_235_io_in; // @[RegFile.scala 66:20:@37546.4]
  wire  regs_235_io_reset; // @[RegFile.scala 66:20:@37546.4]
  wire [63:0] regs_235_io_out; // @[RegFile.scala 66:20:@37546.4]
  wire  regs_235_io_enable; // @[RegFile.scala 66:20:@37546.4]
  wire  regs_236_clock; // @[RegFile.scala 66:20:@37560.4]
  wire  regs_236_reset; // @[RegFile.scala 66:20:@37560.4]
  wire [63:0] regs_236_io_in; // @[RegFile.scala 66:20:@37560.4]
  wire  regs_236_io_reset; // @[RegFile.scala 66:20:@37560.4]
  wire [63:0] regs_236_io_out; // @[RegFile.scala 66:20:@37560.4]
  wire  regs_236_io_enable; // @[RegFile.scala 66:20:@37560.4]
  wire  regs_237_clock; // @[RegFile.scala 66:20:@37574.4]
  wire  regs_237_reset; // @[RegFile.scala 66:20:@37574.4]
  wire [63:0] regs_237_io_in; // @[RegFile.scala 66:20:@37574.4]
  wire  regs_237_io_reset; // @[RegFile.scala 66:20:@37574.4]
  wire [63:0] regs_237_io_out; // @[RegFile.scala 66:20:@37574.4]
  wire  regs_237_io_enable; // @[RegFile.scala 66:20:@37574.4]
  wire  regs_238_clock; // @[RegFile.scala 66:20:@37588.4]
  wire  regs_238_reset; // @[RegFile.scala 66:20:@37588.4]
  wire [63:0] regs_238_io_in; // @[RegFile.scala 66:20:@37588.4]
  wire  regs_238_io_reset; // @[RegFile.scala 66:20:@37588.4]
  wire [63:0] regs_238_io_out; // @[RegFile.scala 66:20:@37588.4]
  wire  regs_238_io_enable; // @[RegFile.scala 66:20:@37588.4]
  wire  regs_239_clock; // @[RegFile.scala 66:20:@37602.4]
  wire  regs_239_reset; // @[RegFile.scala 66:20:@37602.4]
  wire [63:0] regs_239_io_in; // @[RegFile.scala 66:20:@37602.4]
  wire  regs_239_io_reset; // @[RegFile.scala 66:20:@37602.4]
  wire [63:0] regs_239_io_out; // @[RegFile.scala 66:20:@37602.4]
  wire  regs_239_io_enable; // @[RegFile.scala 66:20:@37602.4]
  wire  regs_240_clock; // @[RegFile.scala 66:20:@37616.4]
  wire  regs_240_reset; // @[RegFile.scala 66:20:@37616.4]
  wire [63:0] regs_240_io_in; // @[RegFile.scala 66:20:@37616.4]
  wire  regs_240_io_reset; // @[RegFile.scala 66:20:@37616.4]
  wire [63:0] regs_240_io_out; // @[RegFile.scala 66:20:@37616.4]
  wire  regs_240_io_enable; // @[RegFile.scala 66:20:@37616.4]
  wire  regs_241_clock; // @[RegFile.scala 66:20:@37630.4]
  wire  regs_241_reset; // @[RegFile.scala 66:20:@37630.4]
  wire [63:0] regs_241_io_in; // @[RegFile.scala 66:20:@37630.4]
  wire  regs_241_io_reset; // @[RegFile.scala 66:20:@37630.4]
  wire [63:0] regs_241_io_out; // @[RegFile.scala 66:20:@37630.4]
  wire  regs_241_io_enable; // @[RegFile.scala 66:20:@37630.4]
  wire  regs_242_clock; // @[RegFile.scala 66:20:@37644.4]
  wire  regs_242_reset; // @[RegFile.scala 66:20:@37644.4]
  wire [63:0] regs_242_io_in; // @[RegFile.scala 66:20:@37644.4]
  wire  regs_242_io_reset; // @[RegFile.scala 66:20:@37644.4]
  wire [63:0] regs_242_io_out; // @[RegFile.scala 66:20:@37644.4]
  wire  regs_242_io_enable; // @[RegFile.scala 66:20:@37644.4]
  wire  regs_243_clock; // @[RegFile.scala 66:20:@37658.4]
  wire  regs_243_reset; // @[RegFile.scala 66:20:@37658.4]
  wire [63:0] regs_243_io_in; // @[RegFile.scala 66:20:@37658.4]
  wire  regs_243_io_reset; // @[RegFile.scala 66:20:@37658.4]
  wire [63:0] regs_243_io_out; // @[RegFile.scala 66:20:@37658.4]
  wire  regs_243_io_enable; // @[RegFile.scala 66:20:@37658.4]
  wire  regs_244_clock; // @[RegFile.scala 66:20:@37672.4]
  wire  regs_244_reset; // @[RegFile.scala 66:20:@37672.4]
  wire [63:0] regs_244_io_in; // @[RegFile.scala 66:20:@37672.4]
  wire  regs_244_io_reset; // @[RegFile.scala 66:20:@37672.4]
  wire [63:0] regs_244_io_out; // @[RegFile.scala 66:20:@37672.4]
  wire  regs_244_io_enable; // @[RegFile.scala 66:20:@37672.4]
  wire  regs_245_clock; // @[RegFile.scala 66:20:@37686.4]
  wire  regs_245_reset; // @[RegFile.scala 66:20:@37686.4]
  wire [63:0] regs_245_io_in; // @[RegFile.scala 66:20:@37686.4]
  wire  regs_245_io_reset; // @[RegFile.scala 66:20:@37686.4]
  wire [63:0] regs_245_io_out; // @[RegFile.scala 66:20:@37686.4]
  wire  regs_245_io_enable; // @[RegFile.scala 66:20:@37686.4]
  wire  regs_246_clock; // @[RegFile.scala 66:20:@37700.4]
  wire  regs_246_reset; // @[RegFile.scala 66:20:@37700.4]
  wire [63:0] regs_246_io_in; // @[RegFile.scala 66:20:@37700.4]
  wire  regs_246_io_reset; // @[RegFile.scala 66:20:@37700.4]
  wire [63:0] regs_246_io_out; // @[RegFile.scala 66:20:@37700.4]
  wire  regs_246_io_enable; // @[RegFile.scala 66:20:@37700.4]
  wire  regs_247_clock; // @[RegFile.scala 66:20:@37714.4]
  wire  regs_247_reset; // @[RegFile.scala 66:20:@37714.4]
  wire [63:0] regs_247_io_in; // @[RegFile.scala 66:20:@37714.4]
  wire  regs_247_io_reset; // @[RegFile.scala 66:20:@37714.4]
  wire [63:0] regs_247_io_out; // @[RegFile.scala 66:20:@37714.4]
  wire  regs_247_io_enable; // @[RegFile.scala 66:20:@37714.4]
  wire  regs_248_clock; // @[RegFile.scala 66:20:@37728.4]
  wire  regs_248_reset; // @[RegFile.scala 66:20:@37728.4]
  wire [63:0] regs_248_io_in; // @[RegFile.scala 66:20:@37728.4]
  wire  regs_248_io_reset; // @[RegFile.scala 66:20:@37728.4]
  wire [63:0] regs_248_io_out; // @[RegFile.scala 66:20:@37728.4]
  wire  regs_248_io_enable; // @[RegFile.scala 66:20:@37728.4]
  wire  regs_249_clock; // @[RegFile.scala 66:20:@37742.4]
  wire  regs_249_reset; // @[RegFile.scala 66:20:@37742.4]
  wire [63:0] regs_249_io_in; // @[RegFile.scala 66:20:@37742.4]
  wire  regs_249_io_reset; // @[RegFile.scala 66:20:@37742.4]
  wire [63:0] regs_249_io_out; // @[RegFile.scala 66:20:@37742.4]
  wire  regs_249_io_enable; // @[RegFile.scala 66:20:@37742.4]
  wire  regs_250_clock; // @[RegFile.scala 66:20:@37756.4]
  wire  regs_250_reset; // @[RegFile.scala 66:20:@37756.4]
  wire [63:0] regs_250_io_in; // @[RegFile.scala 66:20:@37756.4]
  wire  regs_250_io_reset; // @[RegFile.scala 66:20:@37756.4]
  wire [63:0] regs_250_io_out; // @[RegFile.scala 66:20:@37756.4]
  wire  regs_250_io_enable; // @[RegFile.scala 66:20:@37756.4]
  wire  regs_251_clock; // @[RegFile.scala 66:20:@37770.4]
  wire  regs_251_reset; // @[RegFile.scala 66:20:@37770.4]
  wire [63:0] regs_251_io_in; // @[RegFile.scala 66:20:@37770.4]
  wire  regs_251_io_reset; // @[RegFile.scala 66:20:@37770.4]
  wire [63:0] regs_251_io_out; // @[RegFile.scala 66:20:@37770.4]
  wire  regs_251_io_enable; // @[RegFile.scala 66:20:@37770.4]
  wire  regs_252_clock; // @[RegFile.scala 66:20:@37784.4]
  wire  regs_252_reset; // @[RegFile.scala 66:20:@37784.4]
  wire [63:0] regs_252_io_in; // @[RegFile.scala 66:20:@37784.4]
  wire  regs_252_io_reset; // @[RegFile.scala 66:20:@37784.4]
  wire [63:0] regs_252_io_out; // @[RegFile.scala 66:20:@37784.4]
  wire  regs_252_io_enable; // @[RegFile.scala 66:20:@37784.4]
  wire  regs_253_clock; // @[RegFile.scala 66:20:@37798.4]
  wire  regs_253_reset; // @[RegFile.scala 66:20:@37798.4]
  wire [63:0] regs_253_io_in; // @[RegFile.scala 66:20:@37798.4]
  wire  regs_253_io_reset; // @[RegFile.scala 66:20:@37798.4]
  wire [63:0] regs_253_io_out; // @[RegFile.scala 66:20:@37798.4]
  wire  regs_253_io_enable; // @[RegFile.scala 66:20:@37798.4]
  wire  regs_254_clock; // @[RegFile.scala 66:20:@37812.4]
  wire  regs_254_reset; // @[RegFile.scala 66:20:@37812.4]
  wire [63:0] regs_254_io_in; // @[RegFile.scala 66:20:@37812.4]
  wire  regs_254_io_reset; // @[RegFile.scala 66:20:@37812.4]
  wire [63:0] regs_254_io_out; // @[RegFile.scala 66:20:@37812.4]
  wire  regs_254_io_enable; // @[RegFile.scala 66:20:@37812.4]
  wire  regs_255_clock; // @[RegFile.scala 66:20:@37826.4]
  wire  regs_255_reset; // @[RegFile.scala 66:20:@37826.4]
  wire [63:0] regs_255_io_in; // @[RegFile.scala 66:20:@37826.4]
  wire  regs_255_io_reset; // @[RegFile.scala 66:20:@37826.4]
  wire [63:0] regs_255_io_out; // @[RegFile.scala 66:20:@37826.4]
  wire  regs_255_io_enable; // @[RegFile.scala 66:20:@37826.4]
  wire  regs_256_clock; // @[RegFile.scala 66:20:@37840.4]
  wire  regs_256_reset; // @[RegFile.scala 66:20:@37840.4]
  wire [63:0] regs_256_io_in; // @[RegFile.scala 66:20:@37840.4]
  wire  regs_256_io_reset; // @[RegFile.scala 66:20:@37840.4]
  wire [63:0] regs_256_io_out; // @[RegFile.scala 66:20:@37840.4]
  wire  regs_256_io_enable; // @[RegFile.scala 66:20:@37840.4]
  wire  regs_257_clock; // @[RegFile.scala 66:20:@37854.4]
  wire  regs_257_reset; // @[RegFile.scala 66:20:@37854.4]
  wire [63:0] regs_257_io_in; // @[RegFile.scala 66:20:@37854.4]
  wire  regs_257_io_reset; // @[RegFile.scala 66:20:@37854.4]
  wire [63:0] regs_257_io_out; // @[RegFile.scala 66:20:@37854.4]
  wire  regs_257_io_enable; // @[RegFile.scala 66:20:@37854.4]
  wire  regs_258_clock; // @[RegFile.scala 66:20:@37868.4]
  wire  regs_258_reset; // @[RegFile.scala 66:20:@37868.4]
  wire [63:0] regs_258_io_in; // @[RegFile.scala 66:20:@37868.4]
  wire  regs_258_io_reset; // @[RegFile.scala 66:20:@37868.4]
  wire [63:0] regs_258_io_out; // @[RegFile.scala 66:20:@37868.4]
  wire  regs_258_io_enable; // @[RegFile.scala 66:20:@37868.4]
  wire  regs_259_clock; // @[RegFile.scala 66:20:@37882.4]
  wire  regs_259_reset; // @[RegFile.scala 66:20:@37882.4]
  wire [63:0] regs_259_io_in; // @[RegFile.scala 66:20:@37882.4]
  wire  regs_259_io_reset; // @[RegFile.scala 66:20:@37882.4]
  wire [63:0] regs_259_io_out; // @[RegFile.scala 66:20:@37882.4]
  wire  regs_259_io_enable; // @[RegFile.scala 66:20:@37882.4]
  wire  regs_260_clock; // @[RegFile.scala 66:20:@37896.4]
  wire  regs_260_reset; // @[RegFile.scala 66:20:@37896.4]
  wire [63:0] regs_260_io_in; // @[RegFile.scala 66:20:@37896.4]
  wire  regs_260_io_reset; // @[RegFile.scala 66:20:@37896.4]
  wire [63:0] regs_260_io_out; // @[RegFile.scala 66:20:@37896.4]
  wire  regs_260_io_enable; // @[RegFile.scala 66:20:@37896.4]
  wire  regs_261_clock; // @[RegFile.scala 66:20:@37910.4]
  wire  regs_261_reset; // @[RegFile.scala 66:20:@37910.4]
  wire [63:0] regs_261_io_in; // @[RegFile.scala 66:20:@37910.4]
  wire  regs_261_io_reset; // @[RegFile.scala 66:20:@37910.4]
  wire [63:0] regs_261_io_out; // @[RegFile.scala 66:20:@37910.4]
  wire  regs_261_io_enable; // @[RegFile.scala 66:20:@37910.4]
  wire  regs_262_clock; // @[RegFile.scala 66:20:@37924.4]
  wire  regs_262_reset; // @[RegFile.scala 66:20:@37924.4]
  wire [63:0] regs_262_io_in; // @[RegFile.scala 66:20:@37924.4]
  wire  regs_262_io_reset; // @[RegFile.scala 66:20:@37924.4]
  wire [63:0] regs_262_io_out; // @[RegFile.scala 66:20:@37924.4]
  wire  regs_262_io_enable; // @[RegFile.scala 66:20:@37924.4]
  wire  regs_263_clock; // @[RegFile.scala 66:20:@37938.4]
  wire  regs_263_reset; // @[RegFile.scala 66:20:@37938.4]
  wire [63:0] regs_263_io_in; // @[RegFile.scala 66:20:@37938.4]
  wire  regs_263_io_reset; // @[RegFile.scala 66:20:@37938.4]
  wire [63:0] regs_263_io_out; // @[RegFile.scala 66:20:@37938.4]
  wire  regs_263_io_enable; // @[RegFile.scala 66:20:@37938.4]
  wire  regs_264_clock; // @[RegFile.scala 66:20:@37952.4]
  wire  regs_264_reset; // @[RegFile.scala 66:20:@37952.4]
  wire [63:0] regs_264_io_in; // @[RegFile.scala 66:20:@37952.4]
  wire  regs_264_io_reset; // @[RegFile.scala 66:20:@37952.4]
  wire [63:0] regs_264_io_out; // @[RegFile.scala 66:20:@37952.4]
  wire  regs_264_io_enable; // @[RegFile.scala 66:20:@37952.4]
  wire  regs_265_clock; // @[RegFile.scala 66:20:@37966.4]
  wire  regs_265_reset; // @[RegFile.scala 66:20:@37966.4]
  wire [63:0] regs_265_io_in; // @[RegFile.scala 66:20:@37966.4]
  wire  regs_265_io_reset; // @[RegFile.scala 66:20:@37966.4]
  wire [63:0] regs_265_io_out; // @[RegFile.scala 66:20:@37966.4]
  wire  regs_265_io_enable; // @[RegFile.scala 66:20:@37966.4]
  wire  regs_266_clock; // @[RegFile.scala 66:20:@37980.4]
  wire  regs_266_reset; // @[RegFile.scala 66:20:@37980.4]
  wire [63:0] regs_266_io_in; // @[RegFile.scala 66:20:@37980.4]
  wire  regs_266_io_reset; // @[RegFile.scala 66:20:@37980.4]
  wire [63:0] regs_266_io_out; // @[RegFile.scala 66:20:@37980.4]
  wire  regs_266_io_enable; // @[RegFile.scala 66:20:@37980.4]
  wire  regs_267_clock; // @[RegFile.scala 66:20:@37994.4]
  wire  regs_267_reset; // @[RegFile.scala 66:20:@37994.4]
  wire [63:0] regs_267_io_in; // @[RegFile.scala 66:20:@37994.4]
  wire  regs_267_io_reset; // @[RegFile.scala 66:20:@37994.4]
  wire [63:0] regs_267_io_out; // @[RegFile.scala 66:20:@37994.4]
  wire  regs_267_io_enable; // @[RegFile.scala 66:20:@37994.4]
  wire  regs_268_clock; // @[RegFile.scala 66:20:@38008.4]
  wire  regs_268_reset; // @[RegFile.scala 66:20:@38008.4]
  wire [63:0] regs_268_io_in; // @[RegFile.scala 66:20:@38008.4]
  wire  regs_268_io_reset; // @[RegFile.scala 66:20:@38008.4]
  wire [63:0] regs_268_io_out; // @[RegFile.scala 66:20:@38008.4]
  wire  regs_268_io_enable; // @[RegFile.scala 66:20:@38008.4]
  wire  regs_269_clock; // @[RegFile.scala 66:20:@38022.4]
  wire  regs_269_reset; // @[RegFile.scala 66:20:@38022.4]
  wire [63:0] regs_269_io_in; // @[RegFile.scala 66:20:@38022.4]
  wire  regs_269_io_reset; // @[RegFile.scala 66:20:@38022.4]
  wire [63:0] regs_269_io_out; // @[RegFile.scala 66:20:@38022.4]
  wire  regs_269_io_enable; // @[RegFile.scala 66:20:@38022.4]
  wire  regs_270_clock; // @[RegFile.scala 66:20:@38036.4]
  wire  regs_270_reset; // @[RegFile.scala 66:20:@38036.4]
  wire [63:0] regs_270_io_in; // @[RegFile.scala 66:20:@38036.4]
  wire  regs_270_io_reset; // @[RegFile.scala 66:20:@38036.4]
  wire [63:0] regs_270_io_out; // @[RegFile.scala 66:20:@38036.4]
  wire  regs_270_io_enable; // @[RegFile.scala 66:20:@38036.4]
  wire  regs_271_clock; // @[RegFile.scala 66:20:@38050.4]
  wire  regs_271_reset; // @[RegFile.scala 66:20:@38050.4]
  wire [63:0] regs_271_io_in; // @[RegFile.scala 66:20:@38050.4]
  wire  regs_271_io_reset; // @[RegFile.scala 66:20:@38050.4]
  wire [63:0] regs_271_io_out; // @[RegFile.scala 66:20:@38050.4]
  wire  regs_271_io_enable; // @[RegFile.scala 66:20:@38050.4]
  wire  regs_272_clock; // @[RegFile.scala 66:20:@38064.4]
  wire  regs_272_reset; // @[RegFile.scala 66:20:@38064.4]
  wire [63:0] regs_272_io_in; // @[RegFile.scala 66:20:@38064.4]
  wire  regs_272_io_reset; // @[RegFile.scala 66:20:@38064.4]
  wire [63:0] regs_272_io_out; // @[RegFile.scala 66:20:@38064.4]
  wire  regs_272_io_enable; // @[RegFile.scala 66:20:@38064.4]
  wire  regs_273_clock; // @[RegFile.scala 66:20:@38078.4]
  wire  regs_273_reset; // @[RegFile.scala 66:20:@38078.4]
  wire [63:0] regs_273_io_in; // @[RegFile.scala 66:20:@38078.4]
  wire  regs_273_io_reset; // @[RegFile.scala 66:20:@38078.4]
  wire [63:0] regs_273_io_out; // @[RegFile.scala 66:20:@38078.4]
  wire  regs_273_io_enable; // @[RegFile.scala 66:20:@38078.4]
  wire  regs_274_clock; // @[RegFile.scala 66:20:@38092.4]
  wire  regs_274_reset; // @[RegFile.scala 66:20:@38092.4]
  wire [63:0] regs_274_io_in; // @[RegFile.scala 66:20:@38092.4]
  wire  regs_274_io_reset; // @[RegFile.scala 66:20:@38092.4]
  wire [63:0] regs_274_io_out; // @[RegFile.scala 66:20:@38092.4]
  wire  regs_274_io_enable; // @[RegFile.scala 66:20:@38092.4]
  wire  regs_275_clock; // @[RegFile.scala 66:20:@38106.4]
  wire  regs_275_reset; // @[RegFile.scala 66:20:@38106.4]
  wire [63:0] regs_275_io_in; // @[RegFile.scala 66:20:@38106.4]
  wire  regs_275_io_reset; // @[RegFile.scala 66:20:@38106.4]
  wire [63:0] regs_275_io_out; // @[RegFile.scala 66:20:@38106.4]
  wire  regs_275_io_enable; // @[RegFile.scala 66:20:@38106.4]
  wire  regs_276_clock; // @[RegFile.scala 66:20:@38120.4]
  wire  regs_276_reset; // @[RegFile.scala 66:20:@38120.4]
  wire [63:0] regs_276_io_in; // @[RegFile.scala 66:20:@38120.4]
  wire  regs_276_io_reset; // @[RegFile.scala 66:20:@38120.4]
  wire [63:0] regs_276_io_out; // @[RegFile.scala 66:20:@38120.4]
  wire  regs_276_io_enable; // @[RegFile.scala 66:20:@38120.4]
  wire  regs_277_clock; // @[RegFile.scala 66:20:@38134.4]
  wire  regs_277_reset; // @[RegFile.scala 66:20:@38134.4]
  wire [63:0] regs_277_io_in; // @[RegFile.scala 66:20:@38134.4]
  wire  regs_277_io_reset; // @[RegFile.scala 66:20:@38134.4]
  wire [63:0] regs_277_io_out; // @[RegFile.scala 66:20:@38134.4]
  wire  regs_277_io_enable; // @[RegFile.scala 66:20:@38134.4]
  wire  regs_278_clock; // @[RegFile.scala 66:20:@38148.4]
  wire  regs_278_reset; // @[RegFile.scala 66:20:@38148.4]
  wire [63:0] regs_278_io_in; // @[RegFile.scala 66:20:@38148.4]
  wire  regs_278_io_reset; // @[RegFile.scala 66:20:@38148.4]
  wire [63:0] regs_278_io_out; // @[RegFile.scala 66:20:@38148.4]
  wire  regs_278_io_enable; // @[RegFile.scala 66:20:@38148.4]
  wire  regs_279_clock; // @[RegFile.scala 66:20:@38162.4]
  wire  regs_279_reset; // @[RegFile.scala 66:20:@38162.4]
  wire [63:0] regs_279_io_in; // @[RegFile.scala 66:20:@38162.4]
  wire  regs_279_io_reset; // @[RegFile.scala 66:20:@38162.4]
  wire [63:0] regs_279_io_out; // @[RegFile.scala 66:20:@38162.4]
  wire  regs_279_io_enable; // @[RegFile.scala 66:20:@38162.4]
  wire  regs_280_clock; // @[RegFile.scala 66:20:@38176.4]
  wire  regs_280_reset; // @[RegFile.scala 66:20:@38176.4]
  wire [63:0] regs_280_io_in; // @[RegFile.scala 66:20:@38176.4]
  wire  regs_280_io_reset; // @[RegFile.scala 66:20:@38176.4]
  wire [63:0] regs_280_io_out; // @[RegFile.scala 66:20:@38176.4]
  wire  regs_280_io_enable; // @[RegFile.scala 66:20:@38176.4]
  wire  regs_281_clock; // @[RegFile.scala 66:20:@38190.4]
  wire  regs_281_reset; // @[RegFile.scala 66:20:@38190.4]
  wire [63:0] regs_281_io_in; // @[RegFile.scala 66:20:@38190.4]
  wire  regs_281_io_reset; // @[RegFile.scala 66:20:@38190.4]
  wire [63:0] regs_281_io_out; // @[RegFile.scala 66:20:@38190.4]
  wire  regs_281_io_enable; // @[RegFile.scala 66:20:@38190.4]
  wire  regs_282_clock; // @[RegFile.scala 66:20:@38204.4]
  wire  regs_282_reset; // @[RegFile.scala 66:20:@38204.4]
  wire [63:0] regs_282_io_in; // @[RegFile.scala 66:20:@38204.4]
  wire  regs_282_io_reset; // @[RegFile.scala 66:20:@38204.4]
  wire [63:0] regs_282_io_out; // @[RegFile.scala 66:20:@38204.4]
  wire  regs_282_io_enable; // @[RegFile.scala 66:20:@38204.4]
  wire  regs_283_clock; // @[RegFile.scala 66:20:@38218.4]
  wire  regs_283_reset; // @[RegFile.scala 66:20:@38218.4]
  wire [63:0] regs_283_io_in; // @[RegFile.scala 66:20:@38218.4]
  wire  regs_283_io_reset; // @[RegFile.scala 66:20:@38218.4]
  wire [63:0] regs_283_io_out; // @[RegFile.scala 66:20:@38218.4]
  wire  regs_283_io_enable; // @[RegFile.scala 66:20:@38218.4]
  wire  regs_284_clock; // @[RegFile.scala 66:20:@38232.4]
  wire  regs_284_reset; // @[RegFile.scala 66:20:@38232.4]
  wire [63:0] regs_284_io_in; // @[RegFile.scala 66:20:@38232.4]
  wire  regs_284_io_reset; // @[RegFile.scala 66:20:@38232.4]
  wire [63:0] regs_284_io_out; // @[RegFile.scala 66:20:@38232.4]
  wire  regs_284_io_enable; // @[RegFile.scala 66:20:@38232.4]
  wire  regs_285_clock; // @[RegFile.scala 66:20:@38246.4]
  wire  regs_285_reset; // @[RegFile.scala 66:20:@38246.4]
  wire [63:0] regs_285_io_in; // @[RegFile.scala 66:20:@38246.4]
  wire  regs_285_io_reset; // @[RegFile.scala 66:20:@38246.4]
  wire [63:0] regs_285_io_out; // @[RegFile.scala 66:20:@38246.4]
  wire  regs_285_io_enable; // @[RegFile.scala 66:20:@38246.4]
  wire  regs_286_clock; // @[RegFile.scala 66:20:@38260.4]
  wire  regs_286_reset; // @[RegFile.scala 66:20:@38260.4]
  wire [63:0] regs_286_io_in; // @[RegFile.scala 66:20:@38260.4]
  wire  regs_286_io_reset; // @[RegFile.scala 66:20:@38260.4]
  wire [63:0] regs_286_io_out; // @[RegFile.scala 66:20:@38260.4]
  wire  regs_286_io_enable; // @[RegFile.scala 66:20:@38260.4]
  wire  regs_287_clock; // @[RegFile.scala 66:20:@38274.4]
  wire  regs_287_reset; // @[RegFile.scala 66:20:@38274.4]
  wire [63:0] regs_287_io_in; // @[RegFile.scala 66:20:@38274.4]
  wire  regs_287_io_reset; // @[RegFile.scala 66:20:@38274.4]
  wire [63:0] regs_287_io_out; // @[RegFile.scala 66:20:@38274.4]
  wire  regs_287_io_enable; // @[RegFile.scala 66:20:@38274.4]
  wire  regs_288_clock; // @[RegFile.scala 66:20:@38288.4]
  wire  regs_288_reset; // @[RegFile.scala 66:20:@38288.4]
  wire [63:0] regs_288_io_in; // @[RegFile.scala 66:20:@38288.4]
  wire  regs_288_io_reset; // @[RegFile.scala 66:20:@38288.4]
  wire [63:0] regs_288_io_out; // @[RegFile.scala 66:20:@38288.4]
  wire  regs_288_io_enable; // @[RegFile.scala 66:20:@38288.4]
  wire  regs_289_clock; // @[RegFile.scala 66:20:@38302.4]
  wire  regs_289_reset; // @[RegFile.scala 66:20:@38302.4]
  wire [63:0] regs_289_io_in; // @[RegFile.scala 66:20:@38302.4]
  wire  regs_289_io_reset; // @[RegFile.scala 66:20:@38302.4]
  wire [63:0] regs_289_io_out; // @[RegFile.scala 66:20:@38302.4]
  wire  regs_289_io_enable; // @[RegFile.scala 66:20:@38302.4]
  wire  regs_290_clock; // @[RegFile.scala 66:20:@38316.4]
  wire  regs_290_reset; // @[RegFile.scala 66:20:@38316.4]
  wire [63:0] regs_290_io_in; // @[RegFile.scala 66:20:@38316.4]
  wire  regs_290_io_reset; // @[RegFile.scala 66:20:@38316.4]
  wire [63:0] regs_290_io_out; // @[RegFile.scala 66:20:@38316.4]
  wire  regs_290_io_enable; // @[RegFile.scala 66:20:@38316.4]
  wire  regs_291_clock; // @[RegFile.scala 66:20:@38330.4]
  wire  regs_291_reset; // @[RegFile.scala 66:20:@38330.4]
  wire [63:0] regs_291_io_in; // @[RegFile.scala 66:20:@38330.4]
  wire  regs_291_io_reset; // @[RegFile.scala 66:20:@38330.4]
  wire [63:0] regs_291_io_out; // @[RegFile.scala 66:20:@38330.4]
  wire  regs_291_io_enable; // @[RegFile.scala 66:20:@38330.4]
  wire  regs_292_clock; // @[RegFile.scala 66:20:@38344.4]
  wire  regs_292_reset; // @[RegFile.scala 66:20:@38344.4]
  wire [63:0] regs_292_io_in; // @[RegFile.scala 66:20:@38344.4]
  wire  regs_292_io_reset; // @[RegFile.scala 66:20:@38344.4]
  wire [63:0] regs_292_io_out; // @[RegFile.scala 66:20:@38344.4]
  wire  regs_292_io_enable; // @[RegFile.scala 66:20:@38344.4]
  wire  regs_293_clock; // @[RegFile.scala 66:20:@38358.4]
  wire  regs_293_reset; // @[RegFile.scala 66:20:@38358.4]
  wire [63:0] regs_293_io_in; // @[RegFile.scala 66:20:@38358.4]
  wire  regs_293_io_reset; // @[RegFile.scala 66:20:@38358.4]
  wire [63:0] regs_293_io_out; // @[RegFile.scala 66:20:@38358.4]
  wire  regs_293_io_enable; // @[RegFile.scala 66:20:@38358.4]
  wire  regs_294_clock; // @[RegFile.scala 66:20:@38372.4]
  wire  regs_294_reset; // @[RegFile.scala 66:20:@38372.4]
  wire [63:0] regs_294_io_in; // @[RegFile.scala 66:20:@38372.4]
  wire  regs_294_io_reset; // @[RegFile.scala 66:20:@38372.4]
  wire [63:0] regs_294_io_out; // @[RegFile.scala 66:20:@38372.4]
  wire  regs_294_io_enable; // @[RegFile.scala 66:20:@38372.4]
  wire  regs_295_clock; // @[RegFile.scala 66:20:@38386.4]
  wire  regs_295_reset; // @[RegFile.scala 66:20:@38386.4]
  wire [63:0] regs_295_io_in; // @[RegFile.scala 66:20:@38386.4]
  wire  regs_295_io_reset; // @[RegFile.scala 66:20:@38386.4]
  wire [63:0] regs_295_io_out; // @[RegFile.scala 66:20:@38386.4]
  wire  regs_295_io_enable; // @[RegFile.scala 66:20:@38386.4]
  wire  regs_296_clock; // @[RegFile.scala 66:20:@38400.4]
  wire  regs_296_reset; // @[RegFile.scala 66:20:@38400.4]
  wire [63:0] regs_296_io_in; // @[RegFile.scala 66:20:@38400.4]
  wire  regs_296_io_reset; // @[RegFile.scala 66:20:@38400.4]
  wire [63:0] regs_296_io_out; // @[RegFile.scala 66:20:@38400.4]
  wire  regs_296_io_enable; // @[RegFile.scala 66:20:@38400.4]
  wire  regs_297_clock; // @[RegFile.scala 66:20:@38414.4]
  wire  regs_297_reset; // @[RegFile.scala 66:20:@38414.4]
  wire [63:0] regs_297_io_in; // @[RegFile.scala 66:20:@38414.4]
  wire  regs_297_io_reset; // @[RegFile.scala 66:20:@38414.4]
  wire [63:0] regs_297_io_out; // @[RegFile.scala 66:20:@38414.4]
  wire  regs_297_io_enable; // @[RegFile.scala 66:20:@38414.4]
  wire  regs_298_clock; // @[RegFile.scala 66:20:@38428.4]
  wire  regs_298_reset; // @[RegFile.scala 66:20:@38428.4]
  wire [63:0] regs_298_io_in; // @[RegFile.scala 66:20:@38428.4]
  wire  regs_298_io_reset; // @[RegFile.scala 66:20:@38428.4]
  wire [63:0] regs_298_io_out; // @[RegFile.scala 66:20:@38428.4]
  wire  regs_298_io_enable; // @[RegFile.scala 66:20:@38428.4]
  wire  regs_299_clock; // @[RegFile.scala 66:20:@38442.4]
  wire  regs_299_reset; // @[RegFile.scala 66:20:@38442.4]
  wire [63:0] regs_299_io_in; // @[RegFile.scala 66:20:@38442.4]
  wire  regs_299_io_reset; // @[RegFile.scala 66:20:@38442.4]
  wire [63:0] regs_299_io_out; // @[RegFile.scala 66:20:@38442.4]
  wire  regs_299_io_enable; // @[RegFile.scala 66:20:@38442.4]
  wire  regs_300_clock; // @[RegFile.scala 66:20:@38456.4]
  wire  regs_300_reset; // @[RegFile.scala 66:20:@38456.4]
  wire [63:0] regs_300_io_in; // @[RegFile.scala 66:20:@38456.4]
  wire  regs_300_io_reset; // @[RegFile.scala 66:20:@38456.4]
  wire [63:0] regs_300_io_out; // @[RegFile.scala 66:20:@38456.4]
  wire  regs_300_io_enable; // @[RegFile.scala 66:20:@38456.4]
  wire  regs_301_clock; // @[RegFile.scala 66:20:@38470.4]
  wire  regs_301_reset; // @[RegFile.scala 66:20:@38470.4]
  wire [63:0] regs_301_io_in; // @[RegFile.scala 66:20:@38470.4]
  wire  regs_301_io_reset; // @[RegFile.scala 66:20:@38470.4]
  wire [63:0] regs_301_io_out; // @[RegFile.scala 66:20:@38470.4]
  wire  regs_301_io_enable; // @[RegFile.scala 66:20:@38470.4]
  wire  regs_302_clock; // @[RegFile.scala 66:20:@38484.4]
  wire  regs_302_reset; // @[RegFile.scala 66:20:@38484.4]
  wire [63:0] regs_302_io_in; // @[RegFile.scala 66:20:@38484.4]
  wire  regs_302_io_reset; // @[RegFile.scala 66:20:@38484.4]
  wire [63:0] regs_302_io_out; // @[RegFile.scala 66:20:@38484.4]
  wire  regs_302_io_enable; // @[RegFile.scala 66:20:@38484.4]
  wire  regs_303_clock; // @[RegFile.scala 66:20:@38498.4]
  wire  regs_303_reset; // @[RegFile.scala 66:20:@38498.4]
  wire [63:0] regs_303_io_in; // @[RegFile.scala 66:20:@38498.4]
  wire  regs_303_io_reset; // @[RegFile.scala 66:20:@38498.4]
  wire [63:0] regs_303_io_out; // @[RegFile.scala 66:20:@38498.4]
  wire  regs_303_io_enable; // @[RegFile.scala 66:20:@38498.4]
  wire  regs_304_clock; // @[RegFile.scala 66:20:@38512.4]
  wire  regs_304_reset; // @[RegFile.scala 66:20:@38512.4]
  wire [63:0] regs_304_io_in; // @[RegFile.scala 66:20:@38512.4]
  wire  regs_304_io_reset; // @[RegFile.scala 66:20:@38512.4]
  wire [63:0] regs_304_io_out; // @[RegFile.scala 66:20:@38512.4]
  wire  regs_304_io_enable; // @[RegFile.scala 66:20:@38512.4]
  wire  regs_305_clock; // @[RegFile.scala 66:20:@38526.4]
  wire  regs_305_reset; // @[RegFile.scala 66:20:@38526.4]
  wire [63:0] regs_305_io_in; // @[RegFile.scala 66:20:@38526.4]
  wire  regs_305_io_reset; // @[RegFile.scala 66:20:@38526.4]
  wire [63:0] regs_305_io_out; // @[RegFile.scala 66:20:@38526.4]
  wire  regs_305_io_enable; // @[RegFile.scala 66:20:@38526.4]
  wire  regs_306_clock; // @[RegFile.scala 66:20:@38540.4]
  wire  regs_306_reset; // @[RegFile.scala 66:20:@38540.4]
  wire [63:0] regs_306_io_in; // @[RegFile.scala 66:20:@38540.4]
  wire  regs_306_io_reset; // @[RegFile.scala 66:20:@38540.4]
  wire [63:0] regs_306_io_out; // @[RegFile.scala 66:20:@38540.4]
  wire  regs_306_io_enable; // @[RegFile.scala 66:20:@38540.4]
  wire  regs_307_clock; // @[RegFile.scala 66:20:@38554.4]
  wire  regs_307_reset; // @[RegFile.scala 66:20:@38554.4]
  wire [63:0] regs_307_io_in; // @[RegFile.scala 66:20:@38554.4]
  wire  regs_307_io_reset; // @[RegFile.scala 66:20:@38554.4]
  wire [63:0] regs_307_io_out; // @[RegFile.scala 66:20:@38554.4]
  wire  regs_307_io_enable; // @[RegFile.scala 66:20:@38554.4]
  wire  regs_308_clock; // @[RegFile.scala 66:20:@38568.4]
  wire  regs_308_reset; // @[RegFile.scala 66:20:@38568.4]
  wire [63:0] regs_308_io_in; // @[RegFile.scala 66:20:@38568.4]
  wire  regs_308_io_reset; // @[RegFile.scala 66:20:@38568.4]
  wire [63:0] regs_308_io_out; // @[RegFile.scala 66:20:@38568.4]
  wire  regs_308_io_enable; // @[RegFile.scala 66:20:@38568.4]
  wire  regs_309_clock; // @[RegFile.scala 66:20:@38582.4]
  wire  regs_309_reset; // @[RegFile.scala 66:20:@38582.4]
  wire [63:0] regs_309_io_in; // @[RegFile.scala 66:20:@38582.4]
  wire  regs_309_io_reset; // @[RegFile.scala 66:20:@38582.4]
  wire [63:0] regs_309_io_out; // @[RegFile.scala 66:20:@38582.4]
  wire  regs_309_io_enable; // @[RegFile.scala 66:20:@38582.4]
  wire  regs_310_clock; // @[RegFile.scala 66:20:@38596.4]
  wire  regs_310_reset; // @[RegFile.scala 66:20:@38596.4]
  wire [63:0] regs_310_io_in; // @[RegFile.scala 66:20:@38596.4]
  wire  regs_310_io_reset; // @[RegFile.scala 66:20:@38596.4]
  wire [63:0] regs_310_io_out; // @[RegFile.scala 66:20:@38596.4]
  wire  regs_310_io_enable; // @[RegFile.scala 66:20:@38596.4]
  wire  regs_311_clock; // @[RegFile.scala 66:20:@38610.4]
  wire  regs_311_reset; // @[RegFile.scala 66:20:@38610.4]
  wire [63:0] regs_311_io_in; // @[RegFile.scala 66:20:@38610.4]
  wire  regs_311_io_reset; // @[RegFile.scala 66:20:@38610.4]
  wire [63:0] regs_311_io_out; // @[RegFile.scala 66:20:@38610.4]
  wire  regs_311_io_enable; // @[RegFile.scala 66:20:@38610.4]
  wire  regs_312_clock; // @[RegFile.scala 66:20:@38624.4]
  wire  regs_312_reset; // @[RegFile.scala 66:20:@38624.4]
  wire [63:0] regs_312_io_in; // @[RegFile.scala 66:20:@38624.4]
  wire  regs_312_io_reset; // @[RegFile.scala 66:20:@38624.4]
  wire [63:0] regs_312_io_out; // @[RegFile.scala 66:20:@38624.4]
  wire  regs_312_io_enable; // @[RegFile.scala 66:20:@38624.4]
  wire  regs_313_clock; // @[RegFile.scala 66:20:@38638.4]
  wire  regs_313_reset; // @[RegFile.scala 66:20:@38638.4]
  wire [63:0] regs_313_io_in; // @[RegFile.scala 66:20:@38638.4]
  wire  regs_313_io_reset; // @[RegFile.scala 66:20:@38638.4]
  wire [63:0] regs_313_io_out; // @[RegFile.scala 66:20:@38638.4]
  wire  regs_313_io_enable; // @[RegFile.scala 66:20:@38638.4]
  wire  regs_314_clock; // @[RegFile.scala 66:20:@38652.4]
  wire  regs_314_reset; // @[RegFile.scala 66:20:@38652.4]
  wire [63:0] regs_314_io_in; // @[RegFile.scala 66:20:@38652.4]
  wire  regs_314_io_reset; // @[RegFile.scala 66:20:@38652.4]
  wire [63:0] regs_314_io_out; // @[RegFile.scala 66:20:@38652.4]
  wire  regs_314_io_enable; // @[RegFile.scala 66:20:@38652.4]
  wire  regs_315_clock; // @[RegFile.scala 66:20:@38666.4]
  wire  regs_315_reset; // @[RegFile.scala 66:20:@38666.4]
  wire [63:0] regs_315_io_in; // @[RegFile.scala 66:20:@38666.4]
  wire  regs_315_io_reset; // @[RegFile.scala 66:20:@38666.4]
  wire [63:0] regs_315_io_out; // @[RegFile.scala 66:20:@38666.4]
  wire  regs_315_io_enable; // @[RegFile.scala 66:20:@38666.4]
  wire  regs_316_clock; // @[RegFile.scala 66:20:@38680.4]
  wire  regs_316_reset; // @[RegFile.scala 66:20:@38680.4]
  wire [63:0] regs_316_io_in; // @[RegFile.scala 66:20:@38680.4]
  wire  regs_316_io_reset; // @[RegFile.scala 66:20:@38680.4]
  wire [63:0] regs_316_io_out; // @[RegFile.scala 66:20:@38680.4]
  wire  regs_316_io_enable; // @[RegFile.scala 66:20:@38680.4]
  wire  regs_317_clock; // @[RegFile.scala 66:20:@38694.4]
  wire  regs_317_reset; // @[RegFile.scala 66:20:@38694.4]
  wire [63:0] regs_317_io_in; // @[RegFile.scala 66:20:@38694.4]
  wire  regs_317_io_reset; // @[RegFile.scala 66:20:@38694.4]
  wire [63:0] regs_317_io_out; // @[RegFile.scala 66:20:@38694.4]
  wire  regs_317_io_enable; // @[RegFile.scala 66:20:@38694.4]
  wire  regs_318_clock; // @[RegFile.scala 66:20:@38708.4]
  wire  regs_318_reset; // @[RegFile.scala 66:20:@38708.4]
  wire [63:0] regs_318_io_in; // @[RegFile.scala 66:20:@38708.4]
  wire  regs_318_io_reset; // @[RegFile.scala 66:20:@38708.4]
  wire [63:0] regs_318_io_out; // @[RegFile.scala 66:20:@38708.4]
  wire  regs_318_io_enable; // @[RegFile.scala 66:20:@38708.4]
  wire  regs_319_clock; // @[RegFile.scala 66:20:@38722.4]
  wire  regs_319_reset; // @[RegFile.scala 66:20:@38722.4]
  wire [63:0] regs_319_io_in; // @[RegFile.scala 66:20:@38722.4]
  wire  regs_319_io_reset; // @[RegFile.scala 66:20:@38722.4]
  wire [63:0] regs_319_io_out; // @[RegFile.scala 66:20:@38722.4]
  wire  regs_319_io_enable; // @[RegFile.scala 66:20:@38722.4]
  wire  regs_320_clock; // @[RegFile.scala 66:20:@38736.4]
  wire  regs_320_reset; // @[RegFile.scala 66:20:@38736.4]
  wire [63:0] regs_320_io_in; // @[RegFile.scala 66:20:@38736.4]
  wire  regs_320_io_reset; // @[RegFile.scala 66:20:@38736.4]
  wire [63:0] regs_320_io_out; // @[RegFile.scala 66:20:@38736.4]
  wire  regs_320_io_enable; // @[RegFile.scala 66:20:@38736.4]
  wire  regs_321_clock; // @[RegFile.scala 66:20:@38750.4]
  wire  regs_321_reset; // @[RegFile.scala 66:20:@38750.4]
  wire [63:0] regs_321_io_in; // @[RegFile.scala 66:20:@38750.4]
  wire  regs_321_io_reset; // @[RegFile.scala 66:20:@38750.4]
  wire [63:0] regs_321_io_out; // @[RegFile.scala 66:20:@38750.4]
  wire  regs_321_io_enable; // @[RegFile.scala 66:20:@38750.4]
  wire  regs_322_clock; // @[RegFile.scala 66:20:@38764.4]
  wire  regs_322_reset; // @[RegFile.scala 66:20:@38764.4]
  wire [63:0] regs_322_io_in; // @[RegFile.scala 66:20:@38764.4]
  wire  regs_322_io_reset; // @[RegFile.scala 66:20:@38764.4]
  wire [63:0] regs_322_io_out; // @[RegFile.scala 66:20:@38764.4]
  wire  regs_322_io_enable; // @[RegFile.scala 66:20:@38764.4]
  wire  regs_323_clock; // @[RegFile.scala 66:20:@38778.4]
  wire  regs_323_reset; // @[RegFile.scala 66:20:@38778.4]
  wire [63:0] regs_323_io_in; // @[RegFile.scala 66:20:@38778.4]
  wire  regs_323_io_reset; // @[RegFile.scala 66:20:@38778.4]
  wire [63:0] regs_323_io_out; // @[RegFile.scala 66:20:@38778.4]
  wire  regs_323_io_enable; // @[RegFile.scala 66:20:@38778.4]
  wire  regs_324_clock; // @[RegFile.scala 66:20:@38792.4]
  wire  regs_324_reset; // @[RegFile.scala 66:20:@38792.4]
  wire [63:0] regs_324_io_in; // @[RegFile.scala 66:20:@38792.4]
  wire  regs_324_io_reset; // @[RegFile.scala 66:20:@38792.4]
  wire [63:0] regs_324_io_out; // @[RegFile.scala 66:20:@38792.4]
  wire  regs_324_io_enable; // @[RegFile.scala 66:20:@38792.4]
  wire  regs_325_clock; // @[RegFile.scala 66:20:@38806.4]
  wire  regs_325_reset; // @[RegFile.scala 66:20:@38806.4]
  wire [63:0] regs_325_io_in; // @[RegFile.scala 66:20:@38806.4]
  wire  regs_325_io_reset; // @[RegFile.scala 66:20:@38806.4]
  wire [63:0] regs_325_io_out; // @[RegFile.scala 66:20:@38806.4]
  wire  regs_325_io_enable; // @[RegFile.scala 66:20:@38806.4]
  wire  regs_326_clock; // @[RegFile.scala 66:20:@38820.4]
  wire  regs_326_reset; // @[RegFile.scala 66:20:@38820.4]
  wire [63:0] regs_326_io_in; // @[RegFile.scala 66:20:@38820.4]
  wire  regs_326_io_reset; // @[RegFile.scala 66:20:@38820.4]
  wire [63:0] regs_326_io_out; // @[RegFile.scala 66:20:@38820.4]
  wire  regs_326_io_enable; // @[RegFile.scala 66:20:@38820.4]
  wire  regs_327_clock; // @[RegFile.scala 66:20:@38834.4]
  wire  regs_327_reset; // @[RegFile.scala 66:20:@38834.4]
  wire [63:0] regs_327_io_in; // @[RegFile.scala 66:20:@38834.4]
  wire  regs_327_io_reset; // @[RegFile.scala 66:20:@38834.4]
  wire [63:0] regs_327_io_out; // @[RegFile.scala 66:20:@38834.4]
  wire  regs_327_io_enable; // @[RegFile.scala 66:20:@38834.4]
  wire  regs_328_clock; // @[RegFile.scala 66:20:@38848.4]
  wire  regs_328_reset; // @[RegFile.scala 66:20:@38848.4]
  wire [63:0] regs_328_io_in; // @[RegFile.scala 66:20:@38848.4]
  wire  regs_328_io_reset; // @[RegFile.scala 66:20:@38848.4]
  wire [63:0] regs_328_io_out; // @[RegFile.scala 66:20:@38848.4]
  wire  regs_328_io_enable; // @[RegFile.scala 66:20:@38848.4]
  wire  regs_329_clock; // @[RegFile.scala 66:20:@38862.4]
  wire  regs_329_reset; // @[RegFile.scala 66:20:@38862.4]
  wire [63:0] regs_329_io_in; // @[RegFile.scala 66:20:@38862.4]
  wire  regs_329_io_reset; // @[RegFile.scala 66:20:@38862.4]
  wire [63:0] regs_329_io_out; // @[RegFile.scala 66:20:@38862.4]
  wire  regs_329_io_enable; // @[RegFile.scala 66:20:@38862.4]
  wire  regs_330_clock; // @[RegFile.scala 66:20:@38876.4]
  wire  regs_330_reset; // @[RegFile.scala 66:20:@38876.4]
  wire [63:0] regs_330_io_in; // @[RegFile.scala 66:20:@38876.4]
  wire  regs_330_io_reset; // @[RegFile.scala 66:20:@38876.4]
  wire [63:0] regs_330_io_out; // @[RegFile.scala 66:20:@38876.4]
  wire  regs_330_io_enable; // @[RegFile.scala 66:20:@38876.4]
  wire  regs_331_clock; // @[RegFile.scala 66:20:@38890.4]
  wire  regs_331_reset; // @[RegFile.scala 66:20:@38890.4]
  wire [63:0] regs_331_io_in; // @[RegFile.scala 66:20:@38890.4]
  wire  regs_331_io_reset; // @[RegFile.scala 66:20:@38890.4]
  wire [63:0] regs_331_io_out; // @[RegFile.scala 66:20:@38890.4]
  wire  regs_331_io_enable; // @[RegFile.scala 66:20:@38890.4]
  wire  regs_332_clock; // @[RegFile.scala 66:20:@38904.4]
  wire  regs_332_reset; // @[RegFile.scala 66:20:@38904.4]
  wire [63:0] regs_332_io_in; // @[RegFile.scala 66:20:@38904.4]
  wire  regs_332_io_reset; // @[RegFile.scala 66:20:@38904.4]
  wire [63:0] regs_332_io_out; // @[RegFile.scala 66:20:@38904.4]
  wire  regs_332_io_enable; // @[RegFile.scala 66:20:@38904.4]
  wire  regs_333_clock; // @[RegFile.scala 66:20:@38918.4]
  wire  regs_333_reset; // @[RegFile.scala 66:20:@38918.4]
  wire [63:0] regs_333_io_in; // @[RegFile.scala 66:20:@38918.4]
  wire  regs_333_io_reset; // @[RegFile.scala 66:20:@38918.4]
  wire [63:0] regs_333_io_out; // @[RegFile.scala 66:20:@38918.4]
  wire  regs_333_io_enable; // @[RegFile.scala 66:20:@38918.4]
  wire  regs_334_clock; // @[RegFile.scala 66:20:@38932.4]
  wire  regs_334_reset; // @[RegFile.scala 66:20:@38932.4]
  wire [63:0] regs_334_io_in; // @[RegFile.scala 66:20:@38932.4]
  wire  regs_334_io_reset; // @[RegFile.scala 66:20:@38932.4]
  wire [63:0] regs_334_io_out; // @[RegFile.scala 66:20:@38932.4]
  wire  regs_334_io_enable; // @[RegFile.scala 66:20:@38932.4]
  wire  regs_335_clock; // @[RegFile.scala 66:20:@38946.4]
  wire  regs_335_reset; // @[RegFile.scala 66:20:@38946.4]
  wire [63:0] regs_335_io_in; // @[RegFile.scala 66:20:@38946.4]
  wire  regs_335_io_reset; // @[RegFile.scala 66:20:@38946.4]
  wire [63:0] regs_335_io_out; // @[RegFile.scala 66:20:@38946.4]
  wire  regs_335_io_enable; // @[RegFile.scala 66:20:@38946.4]
  wire  regs_336_clock; // @[RegFile.scala 66:20:@38960.4]
  wire  regs_336_reset; // @[RegFile.scala 66:20:@38960.4]
  wire [63:0] regs_336_io_in; // @[RegFile.scala 66:20:@38960.4]
  wire  regs_336_io_reset; // @[RegFile.scala 66:20:@38960.4]
  wire [63:0] regs_336_io_out; // @[RegFile.scala 66:20:@38960.4]
  wire  regs_336_io_enable; // @[RegFile.scala 66:20:@38960.4]
  wire  regs_337_clock; // @[RegFile.scala 66:20:@38974.4]
  wire  regs_337_reset; // @[RegFile.scala 66:20:@38974.4]
  wire [63:0] regs_337_io_in; // @[RegFile.scala 66:20:@38974.4]
  wire  regs_337_io_reset; // @[RegFile.scala 66:20:@38974.4]
  wire [63:0] regs_337_io_out; // @[RegFile.scala 66:20:@38974.4]
  wire  regs_337_io_enable; // @[RegFile.scala 66:20:@38974.4]
  wire  regs_338_clock; // @[RegFile.scala 66:20:@38988.4]
  wire  regs_338_reset; // @[RegFile.scala 66:20:@38988.4]
  wire [63:0] regs_338_io_in; // @[RegFile.scala 66:20:@38988.4]
  wire  regs_338_io_reset; // @[RegFile.scala 66:20:@38988.4]
  wire [63:0] regs_338_io_out; // @[RegFile.scala 66:20:@38988.4]
  wire  regs_338_io_enable; // @[RegFile.scala 66:20:@38988.4]
  wire  regs_339_clock; // @[RegFile.scala 66:20:@39002.4]
  wire  regs_339_reset; // @[RegFile.scala 66:20:@39002.4]
  wire [63:0] regs_339_io_in; // @[RegFile.scala 66:20:@39002.4]
  wire  regs_339_io_reset; // @[RegFile.scala 66:20:@39002.4]
  wire [63:0] regs_339_io_out; // @[RegFile.scala 66:20:@39002.4]
  wire  regs_339_io_enable; // @[RegFile.scala 66:20:@39002.4]
  wire  regs_340_clock; // @[RegFile.scala 66:20:@39016.4]
  wire  regs_340_reset; // @[RegFile.scala 66:20:@39016.4]
  wire [63:0] regs_340_io_in; // @[RegFile.scala 66:20:@39016.4]
  wire  regs_340_io_reset; // @[RegFile.scala 66:20:@39016.4]
  wire [63:0] regs_340_io_out; // @[RegFile.scala 66:20:@39016.4]
  wire  regs_340_io_enable; // @[RegFile.scala 66:20:@39016.4]
  wire  regs_341_clock; // @[RegFile.scala 66:20:@39030.4]
  wire  regs_341_reset; // @[RegFile.scala 66:20:@39030.4]
  wire [63:0] regs_341_io_in; // @[RegFile.scala 66:20:@39030.4]
  wire  regs_341_io_reset; // @[RegFile.scala 66:20:@39030.4]
  wire [63:0] regs_341_io_out; // @[RegFile.scala 66:20:@39030.4]
  wire  regs_341_io_enable; // @[RegFile.scala 66:20:@39030.4]
  wire  regs_342_clock; // @[RegFile.scala 66:20:@39044.4]
  wire  regs_342_reset; // @[RegFile.scala 66:20:@39044.4]
  wire [63:0] regs_342_io_in; // @[RegFile.scala 66:20:@39044.4]
  wire  regs_342_io_reset; // @[RegFile.scala 66:20:@39044.4]
  wire [63:0] regs_342_io_out; // @[RegFile.scala 66:20:@39044.4]
  wire  regs_342_io_enable; // @[RegFile.scala 66:20:@39044.4]
  wire  regs_343_clock; // @[RegFile.scala 66:20:@39058.4]
  wire  regs_343_reset; // @[RegFile.scala 66:20:@39058.4]
  wire [63:0] regs_343_io_in; // @[RegFile.scala 66:20:@39058.4]
  wire  regs_343_io_reset; // @[RegFile.scala 66:20:@39058.4]
  wire [63:0] regs_343_io_out; // @[RegFile.scala 66:20:@39058.4]
  wire  regs_343_io_enable; // @[RegFile.scala 66:20:@39058.4]
  wire  regs_344_clock; // @[RegFile.scala 66:20:@39072.4]
  wire  regs_344_reset; // @[RegFile.scala 66:20:@39072.4]
  wire [63:0] regs_344_io_in; // @[RegFile.scala 66:20:@39072.4]
  wire  regs_344_io_reset; // @[RegFile.scala 66:20:@39072.4]
  wire [63:0] regs_344_io_out; // @[RegFile.scala 66:20:@39072.4]
  wire  regs_344_io_enable; // @[RegFile.scala 66:20:@39072.4]
  wire  regs_345_clock; // @[RegFile.scala 66:20:@39086.4]
  wire  regs_345_reset; // @[RegFile.scala 66:20:@39086.4]
  wire [63:0] regs_345_io_in; // @[RegFile.scala 66:20:@39086.4]
  wire  regs_345_io_reset; // @[RegFile.scala 66:20:@39086.4]
  wire [63:0] regs_345_io_out; // @[RegFile.scala 66:20:@39086.4]
  wire  regs_345_io_enable; // @[RegFile.scala 66:20:@39086.4]
  wire  regs_346_clock; // @[RegFile.scala 66:20:@39100.4]
  wire  regs_346_reset; // @[RegFile.scala 66:20:@39100.4]
  wire [63:0] regs_346_io_in; // @[RegFile.scala 66:20:@39100.4]
  wire  regs_346_io_reset; // @[RegFile.scala 66:20:@39100.4]
  wire [63:0] regs_346_io_out; // @[RegFile.scala 66:20:@39100.4]
  wire  regs_346_io_enable; // @[RegFile.scala 66:20:@39100.4]
  wire  regs_347_clock; // @[RegFile.scala 66:20:@39114.4]
  wire  regs_347_reset; // @[RegFile.scala 66:20:@39114.4]
  wire [63:0] regs_347_io_in; // @[RegFile.scala 66:20:@39114.4]
  wire  regs_347_io_reset; // @[RegFile.scala 66:20:@39114.4]
  wire [63:0] regs_347_io_out; // @[RegFile.scala 66:20:@39114.4]
  wire  regs_347_io_enable; // @[RegFile.scala 66:20:@39114.4]
  wire  regs_348_clock; // @[RegFile.scala 66:20:@39128.4]
  wire  regs_348_reset; // @[RegFile.scala 66:20:@39128.4]
  wire [63:0] regs_348_io_in; // @[RegFile.scala 66:20:@39128.4]
  wire  regs_348_io_reset; // @[RegFile.scala 66:20:@39128.4]
  wire [63:0] regs_348_io_out; // @[RegFile.scala 66:20:@39128.4]
  wire  regs_348_io_enable; // @[RegFile.scala 66:20:@39128.4]
  wire  regs_349_clock; // @[RegFile.scala 66:20:@39142.4]
  wire  regs_349_reset; // @[RegFile.scala 66:20:@39142.4]
  wire [63:0] regs_349_io_in; // @[RegFile.scala 66:20:@39142.4]
  wire  regs_349_io_reset; // @[RegFile.scala 66:20:@39142.4]
  wire [63:0] regs_349_io_out; // @[RegFile.scala 66:20:@39142.4]
  wire  regs_349_io_enable; // @[RegFile.scala 66:20:@39142.4]
  wire  regs_350_clock; // @[RegFile.scala 66:20:@39156.4]
  wire  regs_350_reset; // @[RegFile.scala 66:20:@39156.4]
  wire [63:0] regs_350_io_in; // @[RegFile.scala 66:20:@39156.4]
  wire  regs_350_io_reset; // @[RegFile.scala 66:20:@39156.4]
  wire [63:0] regs_350_io_out; // @[RegFile.scala 66:20:@39156.4]
  wire  regs_350_io_enable; // @[RegFile.scala 66:20:@39156.4]
  wire  regs_351_clock; // @[RegFile.scala 66:20:@39170.4]
  wire  regs_351_reset; // @[RegFile.scala 66:20:@39170.4]
  wire [63:0] regs_351_io_in; // @[RegFile.scala 66:20:@39170.4]
  wire  regs_351_io_reset; // @[RegFile.scala 66:20:@39170.4]
  wire [63:0] regs_351_io_out; // @[RegFile.scala 66:20:@39170.4]
  wire  regs_351_io_enable; // @[RegFile.scala 66:20:@39170.4]
  wire  regs_352_clock; // @[RegFile.scala 66:20:@39184.4]
  wire  regs_352_reset; // @[RegFile.scala 66:20:@39184.4]
  wire [63:0] regs_352_io_in; // @[RegFile.scala 66:20:@39184.4]
  wire  regs_352_io_reset; // @[RegFile.scala 66:20:@39184.4]
  wire [63:0] regs_352_io_out; // @[RegFile.scala 66:20:@39184.4]
  wire  regs_352_io_enable; // @[RegFile.scala 66:20:@39184.4]
  wire  regs_353_clock; // @[RegFile.scala 66:20:@39198.4]
  wire  regs_353_reset; // @[RegFile.scala 66:20:@39198.4]
  wire [63:0] regs_353_io_in; // @[RegFile.scala 66:20:@39198.4]
  wire  regs_353_io_reset; // @[RegFile.scala 66:20:@39198.4]
  wire [63:0] regs_353_io_out; // @[RegFile.scala 66:20:@39198.4]
  wire  regs_353_io_enable; // @[RegFile.scala 66:20:@39198.4]
  wire  regs_354_clock; // @[RegFile.scala 66:20:@39212.4]
  wire  regs_354_reset; // @[RegFile.scala 66:20:@39212.4]
  wire [63:0] regs_354_io_in; // @[RegFile.scala 66:20:@39212.4]
  wire  regs_354_io_reset; // @[RegFile.scala 66:20:@39212.4]
  wire [63:0] regs_354_io_out; // @[RegFile.scala 66:20:@39212.4]
  wire  regs_354_io_enable; // @[RegFile.scala 66:20:@39212.4]
  wire  regs_355_clock; // @[RegFile.scala 66:20:@39226.4]
  wire  regs_355_reset; // @[RegFile.scala 66:20:@39226.4]
  wire [63:0] regs_355_io_in; // @[RegFile.scala 66:20:@39226.4]
  wire  regs_355_io_reset; // @[RegFile.scala 66:20:@39226.4]
  wire [63:0] regs_355_io_out; // @[RegFile.scala 66:20:@39226.4]
  wire  regs_355_io_enable; // @[RegFile.scala 66:20:@39226.4]
  wire  regs_356_clock; // @[RegFile.scala 66:20:@39240.4]
  wire  regs_356_reset; // @[RegFile.scala 66:20:@39240.4]
  wire [63:0] regs_356_io_in; // @[RegFile.scala 66:20:@39240.4]
  wire  regs_356_io_reset; // @[RegFile.scala 66:20:@39240.4]
  wire [63:0] regs_356_io_out; // @[RegFile.scala 66:20:@39240.4]
  wire  regs_356_io_enable; // @[RegFile.scala 66:20:@39240.4]
  wire  regs_357_clock; // @[RegFile.scala 66:20:@39254.4]
  wire  regs_357_reset; // @[RegFile.scala 66:20:@39254.4]
  wire [63:0] regs_357_io_in; // @[RegFile.scala 66:20:@39254.4]
  wire  regs_357_io_reset; // @[RegFile.scala 66:20:@39254.4]
  wire [63:0] regs_357_io_out; // @[RegFile.scala 66:20:@39254.4]
  wire  regs_357_io_enable; // @[RegFile.scala 66:20:@39254.4]
  wire  regs_358_clock; // @[RegFile.scala 66:20:@39268.4]
  wire  regs_358_reset; // @[RegFile.scala 66:20:@39268.4]
  wire [63:0] regs_358_io_in; // @[RegFile.scala 66:20:@39268.4]
  wire  regs_358_io_reset; // @[RegFile.scala 66:20:@39268.4]
  wire [63:0] regs_358_io_out; // @[RegFile.scala 66:20:@39268.4]
  wire  regs_358_io_enable; // @[RegFile.scala 66:20:@39268.4]
  wire  regs_359_clock; // @[RegFile.scala 66:20:@39282.4]
  wire  regs_359_reset; // @[RegFile.scala 66:20:@39282.4]
  wire [63:0] regs_359_io_in; // @[RegFile.scala 66:20:@39282.4]
  wire  regs_359_io_reset; // @[RegFile.scala 66:20:@39282.4]
  wire [63:0] regs_359_io_out; // @[RegFile.scala 66:20:@39282.4]
  wire  regs_359_io_enable; // @[RegFile.scala 66:20:@39282.4]
  wire  regs_360_clock; // @[RegFile.scala 66:20:@39296.4]
  wire  regs_360_reset; // @[RegFile.scala 66:20:@39296.4]
  wire [63:0] regs_360_io_in; // @[RegFile.scala 66:20:@39296.4]
  wire  regs_360_io_reset; // @[RegFile.scala 66:20:@39296.4]
  wire [63:0] regs_360_io_out; // @[RegFile.scala 66:20:@39296.4]
  wire  regs_360_io_enable; // @[RegFile.scala 66:20:@39296.4]
  wire  regs_361_clock; // @[RegFile.scala 66:20:@39310.4]
  wire  regs_361_reset; // @[RegFile.scala 66:20:@39310.4]
  wire [63:0] regs_361_io_in; // @[RegFile.scala 66:20:@39310.4]
  wire  regs_361_io_reset; // @[RegFile.scala 66:20:@39310.4]
  wire [63:0] regs_361_io_out; // @[RegFile.scala 66:20:@39310.4]
  wire  regs_361_io_enable; // @[RegFile.scala 66:20:@39310.4]
  wire  regs_362_clock; // @[RegFile.scala 66:20:@39324.4]
  wire  regs_362_reset; // @[RegFile.scala 66:20:@39324.4]
  wire [63:0] regs_362_io_in; // @[RegFile.scala 66:20:@39324.4]
  wire  regs_362_io_reset; // @[RegFile.scala 66:20:@39324.4]
  wire [63:0] regs_362_io_out; // @[RegFile.scala 66:20:@39324.4]
  wire  regs_362_io_enable; // @[RegFile.scala 66:20:@39324.4]
  wire  regs_363_clock; // @[RegFile.scala 66:20:@39338.4]
  wire  regs_363_reset; // @[RegFile.scala 66:20:@39338.4]
  wire [63:0] regs_363_io_in; // @[RegFile.scala 66:20:@39338.4]
  wire  regs_363_io_reset; // @[RegFile.scala 66:20:@39338.4]
  wire [63:0] regs_363_io_out; // @[RegFile.scala 66:20:@39338.4]
  wire  regs_363_io_enable; // @[RegFile.scala 66:20:@39338.4]
  wire  regs_364_clock; // @[RegFile.scala 66:20:@39352.4]
  wire  regs_364_reset; // @[RegFile.scala 66:20:@39352.4]
  wire [63:0] regs_364_io_in; // @[RegFile.scala 66:20:@39352.4]
  wire  regs_364_io_reset; // @[RegFile.scala 66:20:@39352.4]
  wire [63:0] regs_364_io_out; // @[RegFile.scala 66:20:@39352.4]
  wire  regs_364_io_enable; // @[RegFile.scala 66:20:@39352.4]
  wire  regs_365_clock; // @[RegFile.scala 66:20:@39366.4]
  wire  regs_365_reset; // @[RegFile.scala 66:20:@39366.4]
  wire [63:0] regs_365_io_in; // @[RegFile.scala 66:20:@39366.4]
  wire  regs_365_io_reset; // @[RegFile.scala 66:20:@39366.4]
  wire [63:0] regs_365_io_out; // @[RegFile.scala 66:20:@39366.4]
  wire  regs_365_io_enable; // @[RegFile.scala 66:20:@39366.4]
  wire  regs_366_clock; // @[RegFile.scala 66:20:@39380.4]
  wire  regs_366_reset; // @[RegFile.scala 66:20:@39380.4]
  wire [63:0] regs_366_io_in; // @[RegFile.scala 66:20:@39380.4]
  wire  regs_366_io_reset; // @[RegFile.scala 66:20:@39380.4]
  wire [63:0] regs_366_io_out; // @[RegFile.scala 66:20:@39380.4]
  wire  regs_366_io_enable; // @[RegFile.scala 66:20:@39380.4]
  wire  regs_367_clock; // @[RegFile.scala 66:20:@39394.4]
  wire  regs_367_reset; // @[RegFile.scala 66:20:@39394.4]
  wire [63:0] regs_367_io_in; // @[RegFile.scala 66:20:@39394.4]
  wire  regs_367_io_reset; // @[RegFile.scala 66:20:@39394.4]
  wire [63:0] regs_367_io_out; // @[RegFile.scala 66:20:@39394.4]
  wire  regs_367_io_enable; // @[RegFile.scala 66:20:@39394.4]
  wire  regs_368_clock; // @[RegFile.scala 66:20:@39408.4]
  wire  regs_368_reset; // @[RegFile.scala 66:20:@39408.4]
  wire [63:0] regs_368_io_in; // @[RegFile.scala 66:20:@39408.4]
  wire  regs_368_io_reset; // @[RegFile.scala 66:20:@39408.4]
  wire [63:0] regs_368_io_out; // @[RegFile.scala 66:20:@39408.4]
  wire  regs_368_io_enable; // @[RegFile.scala 66:20:@39408.4]
  wire  regs_369_clock; // @[RegFile.scala 66:20:@39422.4]
  wire  regs_369_reset; // @[RegFile.scala 66:20:@39422.4]
  wire [63:0] regs_369_io_in; // @[RegFile.scala 66:20:@39422.4]
  wire  regs_369_io_reset; // @[RegFile.scala 66:20:@39422.4]
  wire [63:0] regs_369_io_out; // @[RegFile.scala 66:20:@39422.4]
  wire  regs_369_io_enable; // @[RegFile.scala 66:20:@39422.4]
  wire  regs_370_clock; // @[RegFile.scala 66:20:@39436.4]
  wire  regs_370_reset; // @[RegFile.scala 66:20:@39436.4]
  wire [63:0] regs_370_io_in; // @[RegFile.scala 66:20:@39436.4]
  wire  regs_370_io_reset; // @[RegFile.scala 66:20:@39436.4]
  wire [63:0] regs_370_io_out; // @[RegFile.scala 66:20:@39436.4]
  wire  regs_370_io_enable; // @[RegFile.scala 66:20:@39436.4]
  wire  regs_371_clock; // @[RegFile.scala 66:20:@39450.4]
  wire  regs_371_reset; // @[RegFile.scala 66:20:@39450.4]
  wire [63:0] regs_371_io_in; // @[RegFile.scala 66:20:@39450.4]
  wire  regs_371_io_reset; // @[RegFile.scala 66:20:@39450.4]
  wire [63:0] regs_371_io_out; // @[RegFile.scala 66:20:@39450.4]
  wire  regs_371_io_enable; // @[RegFile.scala 66:20:@39450.4]
  wire  regs_372_clock; // @[RegFile.scala 66:20:@39464.4]
  wire  regs_372_reset; // @[RegFile.scala 66:20:@39464.4]
  wire [63:0] regs_372_io_in; // @[RegFile.scala 66:20:@39464.4]
  wire  regs_372_io_reset; // @[RegFile.scala 66:20:@39464.4]
  wire [63:0] regs_372_io_out; // @[RegFile.scala 66:20:@39464.4]
  wire  regs_372_io_enable; // @[RegFile.scala 66:20:@39464.4]
  wire  regs_373_clock; // @[RegFile.scala 66:20:@39478.4]
  wire  regs_373_reset; // @[RegFile.scala 66:20:@39478.4]
  wire [63:0] regs_373_io_in; // @[RegFile.scala 66:20:@39478.4]
  wire  regs_373_io_reset; // @[RegFile.scala 66:20:@39478.4]
  wire [63:0] regs_373_io_out; // @[RegFile.scala 66:20:@39478.4]
  wire  regs_373_io_enable; // @[RegFile.scala 66:20:@39478.4]
  wire  regs_374_clock; // @[RegFile.scala 66:20:@39492.4]
  wire  regs_374_reset; // @[RegFile.scala 66:20:@39492.4]
  wire [63:0] regs_374_io_in; // @[RegFile.scala 66:20:@39492.4]
  wire  regs_374_io_reset; // @[RegFile.scala 66:20:@39492.4]
  wire [63:0] regs_374_io_out; // @[RegFile.scala 66:20:@39492.4]
  wire  regs_374_io_enable; // @[RegFile.scala 66:20:@39492.4]
  wire  regs_375_clock; // @[RegFile.scala 66:20:@39506.4]
  wire  regs_375_reset; // @[RegFile.scala 66:20:@39506.4]
  wire [63:0] regs_375_io_in; // @[RegFile.scala 66:20:@39506.4]
  wire  regs_375_io_reset; // @[RegFile.scala 66:20:@39506.4]
  wire [63:0] regs_375_io_out; // @[RegFile.scala 66:20:@39506.4]
  wire  regs_375_io_enable; // @[RegFile.scala 66:20:@39506.4]
  wire  regs_376_clock; // @[RegFile.scala 66:20:@39520.4]
  wire  regs_376_reset; // @[RegFile.scala 66:20:@39520.4]
  wire [63:0] regs_376_io_in; // @[RegFile.scala 66:20:@39520.4]
  wire  regs_376_io_reset; // @[RegFile.scala 66:20:@39520.4]
  wire [63:0] regs_376_io_out; // @[RegFile.scala 66:20:@39520.4]
  wire  regs_376_io_enable; // @[RegFile.scala 66:20:@39520.4]
  wire  regs_377_clock; // @[RegFile.scala 66:20:@39534.4]
  wire  regs_377_reset; // @[RegFile.scala 66:20:@39534.4]
  wire [63:0] regs_377_io_in; // @[RegFile.scala 66:20:@39534.4]
  wire  regs_377_io_reset; // @[RegFile.scala 66:20:@39534.4]
  wire [63:0] regs_377_io_out; // @[RegFile.scala 66:20:@39534.4]
  wire  regs_377_io_enable; // @[RegFile.scala 66:20:@39534.4]
  wire  regs_378_clock; // @[RegFile.scala 66:20:@39548.4]
  wire  regs_378_reset; // @[RegFile.scala 66:20:@39548.4]
  wire [63:0] regs_378_io_in; // @[RegFile.scala 66:20:@39548.4]
  wire  regs_378_io_reset; // @[RegFile.scala 66:20:@39548.4]
  wire [63:0] regs_378_io_out; // @[RegFile.scala 66:20:@39548.4]
  wire  regs_378_io_enable; // @[RegFile.scala 66:20:@39548.4]
  wire  regs_379_clock; // @[RegFile.scala 66:20:@39562.4]
  wire  regs_379_reset; // @[RegFile.scala 66:20:@39562.4]
  wire [63:0] regs_379_io_in; // @[RegFile.scala 66:20:@39562.4]
  wire  regs_379_io_reset; // @[RegFile.scala 66:20:@39562.4]
  wire [63:0] regs_379_io_out; // @[RegFile.scala 66:20:@39562.4]
  wire  regs_379_io_enable; // @[RegFile.scala 66:20:@39562.4]
  wire  regs_380_clock; // @[RegFile.scala 66:20:@39576.4]
  wire  regs_380_reset; // @[RegFile.scala 66:20:@39576.4]
  wire [63:0] regs_380_io_in; // @[RegFile.scala 66:20:@39576.4]
  wire  regs_380_io_reset; // @[RegFile.scala 66:20:@39576.4]
  wire [63:0] regs_380_io_out; // @[RegFile.scala 66:20:@39576.4]
  wire  regs_380_io_enable; // @[RegFile.scala 66:20:@39576.4]
  wire  regs_381_clock; // @[RegFile.scala 66:20:@39590.4]
  wire  regs_381_reset; // @[RegFile.scala 66:20:@39590.4]
  wire [63:0] regs_381_io_in; // @[RegFile.scala 66:20:@39590.4]
  wire  regs_381_io_reset; // @[RegFile.scala 66:20:@39590.4]
  wire [63:0] regs_381_io_out; // @[RegFile.scala 66:20:@39590.4]
  wire  regs_381_io_enable; // @[RegFile.scala 66:20:@39590.4]
  wire  regs_382_clock; // @[RegFile.scala 66:20:@39604.4]
  wire  regs_382_reset; // @[RegFile.scala 66:20:@39604.4]
  wire [63:0] regs_382_io_in; // @[RegFile.scala 66:20:@39604.4]
  wire  regs_382_io_reset; // @[RegFile.scala 66:20:@39604.4]
  wire [63:0] regs_382_io_out; // @[RegFile.scala 66:20:@39604.4]
  wire  regs_382_io_enable; // @[RegFile.scala 66:20:@39604.4]
  wire  regs_383_clock; // @[RegFile.scala 66:20:@39618.4]
  wire  regs_383_reset; // @[RegFile.scala 66:20:@39618.4]
  wire [63:0] regs_383_io_in; // @[RegFile.scala 66:20:@39618.4]
  wire  regs_383_io_reset; // @[RegFile.scala 66:20:@39618.4]
  wire [63:0] regs_383_io_out; // @[RegFile.scala 66:20:@39618.4]
  wire  regs_383_io_enable; // @[RegFile.scala 66:20:@39618.4]
  wire  regs_384_clock; // @[RegFile.scala 66:20:@39632.4]
  wire  regs_384_reset; // @[RegFile.scala 66:20:@39632.4]
  wire [63:0] regs_384_io_in; // @[RegFile.scala 66:20:@39632.4]
  wire  regs_384_io_reset; // @[RegFile.scala 66:20:@39632.4]
  wire [63:0] regs_384_io_out; // @[RegFile.scala 66:20:@39632.4]
  wire  regs_384_io_enable; // @[RegFile.scala 66:20:@39632.4]
  wire  regs_385_clock; // @[RegFile.scala 66:20:@39646.4]
  wire  regs_385_reset; // @[RegFile.scala 66:20:@39646.4]
  wire [63:0] regs_385_io_in; // @[RegFile.scala 66:20:@39646.4]
  wire  regs_385_io_reset; // @[RegFile.scala 66:20:@39646.4]
  wire [63:0] regs_385_io_out; // @[RegFile.scala 66:20:@39646.4]
  wire  regs_385_io_enable; // @[RegFile.scala 66:20:@39646.4]
  wire  regs_386_clock; // @[RegFile.scala 66:20:@39660.4]
  wire  regs_386_reset; // @[RegFile.scala 66:20:@39660.4]
  wire [63:0] regs_386_io_in; // @[RegFile.scala 66:20:@39660.4]
  wire  regs_386_io_reset; // @[RegFile.scala 66:20:@39660.4]
  wire [63:0] regs_386_io_out; // @[RegFile.scala 66:20:@39660.4]
  wire  regs_386_io_enable; // @[RegFile.scala 66:20:@39660.4]
  wire  regs_387_clock; // @[RegFile.scala 66:20:@39674.4]
  wire  regs_387_reset; // @[RegFile.scala 66:20:@39674.4]
  wire [63:0] regs_387_io_in; // @[RegFile.scala 66:20:@39674.4]
  wire  regs_387_io_reset; // @[RegFile.scala 66:20:@39674.4]
  wire [63:0] regs_387_io_out; // @[RegFile.scala 66:20:@39674.4]
  wire  regs_387_io_enable; // @[RegFile.scala 66:20:@39674.4]
  wire  regs_388_clock; // @[RegFile.scala 66:20:@39688.4]
  wire  regs_388_reset; // @[RegFile.scala 66:20:@39688.4]
  wire [63:0] regs_388_io_in; // @[RegFile.scala 66:20:@39688.4]
  wire  regs_388_io_reset; // @[RegFile.scala 66:20:@39688.4]
  wire [63:0] regs_388_io_out; // @[RegFile.scala 66:20:@39688.4]
  wire  regs_388_io_enable; // @[RegFile.scala 66:20:@39688.4]
  wire  regs_389_clock; // @[RegFile.scala 66:20:@39702.4]
  wire  regs_389_reset; // @[RegFile.scala 66:20:@39702.4]
  wire [63:0] regs_389_io_in; // @[RegFile.scala 66:20:@39702.4]
  wire  regs_389_io_reset; // @[RegFile.scala 66:20:@39702.4]
  wire [63:0] regs_389_io_out; // @[RegFile.scala 66:20:@39702.4]
  wire  regs_389_io_enable; // @[RegFile.scala 66:20:@39702.4]
  wire  regs_390_clock; // @[RegFile.scala 66:20:@39716.4]
  wire  regs_390_reset; // @[RegFile.scala 66:20:@39716.4]
  wire [63:0] regs_390_io_in; // @[RegFile.scala 66:20:@39716.4]
  wire  regs_390_io_reset; // @[RegFile.scala 66:20:@39716.4]
  wire [63:0] regs_390_io_out; // @[RegFile.scala 66:20:@39716.4]
  wire  regs_390_io_enable; // @[RegFile.scala 66:20:@39716.4]
  wire  regs_391_clock; // @[RegFile.scala 66:20:@39730.4]
  wire  regs_391_reset; // @[RegFile.scala 66:20:@39730.4]
  wire [63:0] regs_391_io_in; // @[RegFile.scala 66:20:@39730.4]
  wire  regs_391_io_reset; // @[RegFile.scala 66:20:@39730.4]
  wire [63:0] regs_391_io_out; // @[RegFile.scala 66:20:@39730.4]
  wire  regs_391_io_enable; // @[RegFile.scala 66:20:@39730.4]
  wire  regs_392_clock; // @[RegFile.scala 66:20:@39744.4]
  wire  regs_392_reset; // @[RegFile.scala 66:20:@39744.4]
  wire [63:0] regs_392_io_in; // @[RegFile.scala 66:20:@39744.4]
  wire  regs_392_io_reset; // @[RegFile.scala 66:20:@39744.4]
  wire [63:0] regs_392_io_out; // @[RegFile.scala 66:20:@39744.4]
  wire  regs_392_io_enable; // @[RegFile.scala 66:20:@39744.4]
  wire  regs_393_clock; // @[RegFile.scala 66:20:@39758.4]
  wire  regs_393_reset; // @[RegFile.scala 66:20:@39758.4]
  wire [63:0] regs_393_io_in; // @[RegFile.scala 66:20:@39758.4]
  wire  regs_393_io_reset; // @[RegFile.scala 66:20:@39758.4]
  wire [63:0] regs_393_io_out; // @[RegFile.scala 66:20:@39758.4]
  wire  regs_393_io_enable; // @[RegFile.scala 66:20:@39758.4]
  wire  regs_394_clock; // @[RegFile.scala 66:20:@39772.4]
  wire  regs_394_reset; // @[RegFile.scala 66:20:@39772.4]
  wire [63:0] regs_394_io_in; // @[RegFile.scala 66:20:@39772.4]
  wire  regs_394_io_reset; // @[RegFile.scala 66:20:@39772.4]
  wire [63:0] regs_394_io_out; // @[RegFile.scala 66:20:@39772.4]
  wire  regs_394_io_enable; // @[RegFile.scala 66:20:@39772.4]
  wire  regs_395_clock; // @[RegFile.scala 66:20:@39786.4]
  wire  regs_395_reset; // @[RegFile.scala 66:20:@39786.4]
  wire [63:0] regs_395_io_in; // @[RegFile.scala 66:20:@39786.4]
  wire  regs_395_io_reset; // @[RegFile.scala 66:20:@39786.4]
  wire [63:0] regs_395_io_out; // @[RegFile.scala 66:20:@39786.4]
  wire  regs_395_io_enable; // @[RegFile.scala 66:20:@39786.4]
  wire  regs_396_clock; // @[RegFile.scala 66:20:@39800.4]
  wire  regs_396_reset; // @[RegFile.scala 66:20:@39800.4]
  wire [63:0] regs_396_io_in; // @[RegFile.scala 66:20:@39800.4]
  wire  regs_396_io_reset; // @[RegFile.scala 66:20:@39800.4]
  wire [63:0] regs_396_io_out; // @[RegFile.scala 66:20:@39800.4]
  wire  regs_396_io_enable; // @[RegFile.scala 66:20:@39800.4]
  wire  regs_397_clock; // @[RegFile.scala 66:20:@39814.4]
  wire  regs_397_reset; // @[RegFile.scala 66:20:@39814.4]
  wire [63:0] regs_397_io_in; // @[RegFile.scala 66:20:@39814.4]
  wire  regs_397_io_reset; // @[RegFile.scala 66:20:@39814.4]
  wire [63:0] regs_397_io_out; // @[RegFile.scala 66:20:@39814.4]
  wire  regs_397_io_enable; // @[RegFile.scala 66:20:@39814.4]
  wire  regs_398_clock; // @[RegFile.scala 66:20:@39828.4]
  wire  regs_398_reset; // @[RegFile.scala 66:20:@39828.4]
  wire [63:0] regs_398_io_in; // @[RegFile.scala 66:20:@39828.4]
  wire  regs_398_io_reset; // @[RegFile.scala 66:20:@39828.4]
  wire [63:0] regs_398_io_out; // @[RegFile.scala 66:20:@39828.4]
  wire  regs_398_io_enable; // @[RegFile.scala 66:20:@39828.4]
  wire  regs_399_clock; // @[RegFile.scala 66:20:@39842.4]
  wire  regs_399_reset; // @[RegFile.scala 66:20:@39842.4]
  wire [63:0] regs_399_io_in; // @[RegFile.scala 66:20:@39842.4]
  wire  regs_399_io_reset; // @[RegFile.scala 66:20:@39842.4]
  wire [63:0] regs_399_io_out; // @[RegFile.scala 66:20:@39842.4]
  wire  regs_399_io_enable; // @[RegFile.scala 66:20:@39842.4]
  wire  regs_400_clock; // @[RegFile.scala 66:20:@39856.4]
  wire  regs_400_reset; // @[RegFile.scala 66:20:@39856.4]
  wire [63:0] regs_400_io_in; // @[RegFile.scala 66:20:@39856.4]
  wire  regs_400_io_reset; // @[RegFile.scala 66:20:@39856.4]
  wire [63:0] regs_400_io_out; // @[RegFile.scala 66:20:@39856.4]
  wire  regs_400_io_enable; // @[RegFile.scala 66:20:@39856.4]
  wire  regs_401_clock; // @[RegFile.scala 66:20:@39870.4]
  wire  regs_401_reset; // @[RegFile.scala 66:20:@39870.4]
  wire [63:0] regs_401_io_in; // @[RegFile.scala 66:20:@39870.4]
  wire  regs_401_io_reset; // @[RegFile.scala 66:20:@39870.4]
  wire [63:0] regs_401_io_out; // @[RegFile.scala 66:20:@39870.4]
  wire  regs_401_io_enable; // @[RegFile.scala 66:20:@39870.4]
  wire  regs_402_clock; // @[RegFile.scala 66:20:@39884.4]
  wire  regs_402_reset; // @[RegFile.scala 66:20:@39884.4]
  wire [63:0] regs_402_io_in; // @[RegFile.scala 66:20:@39884.4]
  wire  regs_402_io_reset; // @[RegFile.scala 66:20:@39884.4]
  wire [63:0] regs_402_io_out; // @[RegFile.scala 66:20:@39884.4]
  wire  regs_402_io_enable; // @[RegFile.scala 66:20:@39884.4]
  wire  regs_403_clock; // @[RegFile.scala 66:20:@39898.4]
  wire  regs_403_reset; // @[RegFile.scala 66:20:@39898.4]
  wire [63:0] regs_403_io_in; // @[RegFile.scala 66:20:@39898.4]
  wire  regs_403_io_reset; // @[RegFile.scala 66:20:@39898.4]
  wire [63:0] regs_403_io_out; // @[RegFile.scala 66:20:@39898.4]
  wire  regs_403_io_enable; // @[RegFile.scala 66:20:@39898.4]
  wire  regs_404_clock; // @[RegFile.scala 66:20:@39912.4]
  wire  regs_404_reset; // @[RegFile.scala 66:20:@39912.4]
  wire [63:0] regs_404_io_in; // @[RegFile.scala 66:20:@39912.4]
  wire  regs_404_io_reset; // @[RegFile.scala 66:20:@39912.4]
  wire [63:0] regs_404_io_out; // @[RegFile.scala 66:20:@39912.4]
  wire  regs_404_io_enable; // @[RegFile.scala 66:20:@39912.4]
  wire  regs_405_clock; // @[RegFile.scala 66:20:@39926.4]
  wire  regs_405_reset; // @[RegFile.scala 66:20:@39926.4]
  wire [63:0] regs_405_io_in; // @[RegFile.scala 66:20:@39926.4]
  wire  regs_405_io_reset; // @[RegFile.scala 66:20:@39926.4]
  wire [63:0] regs_405_io_out; // @[RegFile.scala 66:20:@39926.4]
  wire  regs_405_io_enable; // @[RegFile.scala 66:20:@39926.4]
  wire  regs_406_clock; // @[RegFile.scala 66:20:@39940.4]
  wire  regs_406_reset; // @[RegFile.scala 66:20:@39940.4]
  wire [63:0] regs_406_io_in; // @[RegFile.scala 66:20:@39940.4]
  wire  regs_406_io_reset; // @[RegFile.scala 66:20:@39940.4]
  wire [63:0] regs_406_io_out; // @[RegFile.scala 66:20:@39940.4]
  wire  regs_406_io_enable; // @[RegFile.scala 66:20:@39940.4]
  wire  regs_407_clock; // @[RegFile.scala 66:20:@39954.4]
  wire  regs_407_reset; // @[RegFile.scala 66:20:@39954.4]
  wire [63:0] regs_407_io_in; // @[RegFile.scala 66:20:@39954.4]
  wire  regs_407_io_reset; // @[RegFile.scala 66:20:@39954.4]
  wire [63:0] regs_407_io_out; // @[RegFile.scala 66:20:@39954.4]
  wire  regs_407_io_enable; // @[RegFile.scala 66:20:@39954.4]
  wire  regs_408_clock; // @[RegFile.scala 66:20:@39968.4]
  wire  regs_408_reset; // @[RegFile.scala 66:20:@39968.4]
  wire [63:0] regs_408_io_in; // @[RegFile.scala 66:20:@39968.4]
  wire  regs_408_io_reset; // @[RegFile.scala 66:20:@39968.4]
  wire [63:0] regs_408_io_out; // @[RegFile.scala 66:20:@39968.4]
  wire  regs_408_io_enable; // @[RegFile.scala 66:20:@39968.4]
  wire  regs_409_clock; // @[RegFile.scala 66:20:@39982.4]
  wire  regs_409_reset; // @[RegFile.scala 66:20:@39982.4]
  wire [63:0] regs_409_io_in; // @[RegFile.scala 66:20:@39982.4]
  wire  regs_409_io_reset; // @[RegFile.scala 66:20:@39982.4]
  wire [63:0] regs_409_io_out; // @[RegFile.scala 66:20:@39982.4]
  wire  regs_409_io_enable; // @[RegFile.scala 66:20:@39982.4]
  wire  regs_410_clock; // @[RegFile.scala 66:20:@39996.4]
  wire  regs_410_reset; // @[RegFile.scala 66:20:@39996.4]
  wire [63:0] regs_410_io_in; // @[RegFile.scala 66:20:@39996.4]
  wire  regs_410_io_reset; // @[RegFile.scala 66:20:@39996.4]
  wire [63:0] regs_410_io_out; // @[RegFile.scala 66:20:@39996.4]
  wire  regs_410_io_enable; // @[RegFile.scala 66:20:@39996.4]
  wire  regs_411_clock; // @[RegFile.scala 66:20:@40010.4]
  wire  regs_411_reset; // @[RegFile.scala 66:20:@40010.4]
  wire [63:0] regs_411_io_in; // @[RegFile.scala 66:20:@40010.4]
  wire  regs_411_io_reset; // @[RegFile.scala 66:20:@40010.4]
  wire [63:0] regs_411_io_out; // @[RegFile.scala 66:20:@40010.4]
  wire  regs_411_io_enable; // @[RegFile.scala 66:20:@40010.4]
  wire  regs_412_clock; // @[RegFile.scala 66:20:@40024.4]
  wire  regs_412_reset; // @[RegFile.scala 66:20:@40024.4]
  wire [63:0] regs_412_io_in; // @[RegFile.scala 66:20:@40024.4]
  wire  regs_412_io_reset; // @[RegFile.scala 66:20:@40024.4]
  wire [63:0] regs_412_io_out; // @[RegFile.scala 66:20:@40024.4]
  wire  regs_412_io_enable; // @[RegFile.scala 66:20:@40024.4]
  wire  regs_413_clock; // @[RegFile.scala 66:20:@40038.4]
  wire  regs_413_reset; // @[RegFile.scala 66:20:@40038.4]
  wire [63:0] regs_413_io_in; // @[RegFile.scala 66:20:@40038.4]
  wire  regs_413_io_reset; // @[RegFile.scala 66:20:@40038.4]
  wire [63:0] regs_413_io_out; // @[RegFile.scala 66:20:@40038.4]
  wire  regs_413_io_enable; // @[RegFile.scala 66:20:@40038.4]
  wire  regs_414_clock; // @[RegFile.scala 66:20:@40052.4]
  wire  regs_414_reset; // @[RegFile.scala 66:20:@40052.4]
  wire [63:0] regs_414_io_in; // @[RegFile.scala 66:20:@40052.4]
  wire  regs_414_io_reset; // @[RegFile.scala 66:20:@40052.4]
  wire [63:0] regs_414_io_out; // @[RegFile.scala 66:20:@40052.4]
  wire  regs_414_io_enable; // @[RegFile.scala 66:20:@40052.4]
  wire  regs_415_clock; // @[RegFile.scala 66:20:@40066.4]
  wire  regs_415_reset; // @[RegFile.scala 66:20:@40066.4]
  wire [63:0] regs_415_io_in; // @[RegFile.scala 66:20:@40066.4]
  wire  regs_415_io_reset; // @[RegFile.scala 66:20:@40066.4]
  wire [63:0] regs_415_io_out; // @[RegFile.scala 66:20:@40066.4]
  wire  regs_415_io_enable; // @[RegFile.scala 66:20:@40066.4]
  wire  regs_416_clock; // @[RegFile.scala 66:20:@40080.4]
  wire  regs_416_reset; // @[RegFile.scala 66:20:@40080.4]
  wire [63:0] regs_416_io_in; // @[RegFile.scala 66:20:@40080.4]
  wire  regs_416_io_reset; // @[RegFile.scala 66:20:@40080.4]
  wire [63:0] regs_416_io_out; // @[RegFile.scala 66:20:@40080.4]
  wire  regs_416_io_enable; // @[RegFile.scala 66:20:@40080.4]
  wire  regs_417_clock; // @[RegFile.scala 66:20:@40094.4]
  wire  regs_417_reset; // @[RegFile.scala 66:20:@40094.4]
  wire [63:0] regs_417_io_in; // @[RegFile.scala 66:20:@40094.4]
  wire  regs_417_io_reset; // @[RegFile.scala 66:20:@40094.4]
  wire [63:0] regs_417_io_out; // @[RegFile.scala 66:20:@40094.4]
  wire  regs_417_io_enable; // @[RegFile.scala 66:20:@40094.4]
  wire  regs_418_clock; // @[RegFile.scala 66:20:@40108.4]
  wire  regs_418_reset; // @[RegFile.scala 66:20:@40108.4]
  wire [63:0] regs_418_io_in; // @[RegFile.scala 66:20:@40108.4]
  wire  regs_418_io_reset; // @[RegFile.scala 66:20:@40108.4]
  wire [63:0] regs_418_io_out; // @[RegFile.scala 66:20:@40108.4]
  wire  regs_418_io_enable; // @[RegFile.scala 66:20:@40108.4]
  wire  regs_419_clock; // @[RegFile.scala 66:20:@40122.4]
  wire  regs_419_reset; // @[RegFile.scala 66:20:@40122.4]
  wire [63:0] regs_419_io_in; // @[RegFile.scala 66:20:@40122.4]
  wire  regs_419_io_reset; // @[RegFile.scala 66:20:@40122.4]
  wire [63:0] regs_419_io_out; // @[RegFile.scala 66:20:@40122.4]
  wire  regs_419_io_enable; // @[RegFile.scala 66:20:@40122.4]
  wire  regs_420_clock; // @[RegFile.scala 66:20:@40136.4]
  wire  regs_420_reset; // @[RegFile.scala 66:20:@40136.4]
  wire [63:0] regs_420_io_in; // @[RegFile.scala 66:20:@40136.4]
  wire  regs_420_io_reset; // @[RegFile.scala 66:20:@40136.4]
  wire [63:0] regs_420_io_out; // @[RegFile.scala 66:20:@40136.4]
  wire  regs_420_io_enable; // @[RegFile.scala 66:20:@40136.4]
  wire  regs_421_clock; // @[RegFile.scala 66:20:@40150.4]
  wire  regs_421_reset; // @[RegFile.scala 66:20:@40150.4]
  wire [63:0] regs_421_io_in; // @[RegFile.scala 66:20:@40150.4]
  wire  regs_421_io_reset; // @[RegFile.scala 66:20:@40150.4]
  wire [63:0] regs_421_io_out; // @[RegFile.scala 66:20:@40150.4]
  wire  regs_421_io_enable; // @[RegFile.scala 66:20:@40150.4]
  wire  regs_422_clock; // @[RegFile.scala 66:20:@40164.4]
  wire  regs_422_reset; // @[RegFile.scala 66:20:@40164.4]
  wire [63:0] regs_422_io_in; // @[RegFile.scala 66:20:@40164.4]
  wire  regs_422_io_reset; // @[RegFile.scala 66:20:@40164.4]
  wire [63:0] regs_422_io_out; // @[RegFile.scala 66:20:@40164.4]
  wire  regs_422_io_enable; // @[RegFile.scala 66:20:@40164.4]
  wire  regs_423_clock; // @[RegFile.scala 66:20:@40178.4]
  wire  regs_423_reset; // @[RegFile.scala 66:20:@40178.4]
  wire [63:0] regs_423_io_in; // @[RegFile.scala 66:20:@40178.4]
  wire  regs_423_io_reset; // @[RegFile.scala 66:20:@40178.4]
  wire [63:0] regs_423_io_out; // @[RegFile.scala 66:20:@40178.4]
  wire  regs_423_io_enable; // @[RegFile.scala 66:20:@40178.4]
  wire  regs_424_clock; // @[RegFile.scala 66:20:@40192.4]
  wire  regs_424_reset; // @[RegFile.scala 66:20:@40192.4]
  wire [63:0] regs_424_io_in; // @[RegFile.scala 66:20:@40192.4]
  wire  regs_424_io_reset; // @[RegFile.scala 66:20:@40192.4]
  wire [63:0] regs_424_io_out; // @[RegFile.scala 66:20:@40192.4]
  wire  regs_424_io_enable; // @[RegFile.scala 66:20:@40192.4]
  wire  regs_425_clock; // @[RegFile.scala 66:20:@40206.4]
  wire  regs_425_reset; // @[RegFile.scala 66:20:@40206.4]
  wire [63:0] regs_425_io_in; // @[RegFile.scala 66:20:@40206.4]
  wire  regs_425_io_reset; // @[RegFile.scala 66:20:@40206.4]
  wire [63:0] regs_425_io_out; // @[RegFile.scala 66:20:@40206.4]
  wire  regs_425_io_enable; // @[RegFile.scala 66:20:@40206.4]
  wire  regs_426_clock; // @[RegFile.scala 66:20:@40220.4]
  wire  regs_426_reset; // @[RegFile.scala 66:20:@40220.4]
  wire [63:0] regs_426_io_in; // @[RegFile.scala 66:20:@40220.4]
  wire  regs_426_io_reset; // @[RegFile.scala 66:20:@40220.4]
  wire [63:0] regs_426_io_out; // @[RegFile.scala 66:20:@40220.4]
  wire  regs_426_io_enable; // @[RegFile.scala 66:20:@40220.4]
  wire  regs_427_clock; // @[RegFile.scala 66:20:@40234.4]
  wire  regs_427_reset; // @[RegFile.scala 66:20:@40234.4]
  wire [63:0] regs_427_io_in; // @[RegFile.scala 66:20:@40234.4]
  wire  regs_427_io_reset; // @[RegFile.scala 66:20:@40234.4]
  wire [63:0] regs_427_io_out; // @[RegFile.scala 66:20:@40234.4]
  wire  regs_427_io_enable; // @[RegFile.scala 66:20:@40234.4]
  wire  regs_428_clock; // @[RegFile.scala 66:20:@40248.4]
  wire  regs_428_reset; // @[RegFile.scala 66:20:@40248.4]
  wire [63:0] regs_428_io_in; // @[RegFile.scala 66:20:@40248.4]
  wire  regs_428_io_reset; // @[RegFile.scala 66:20:@40248.4]
  wire [63:0] regs_428_io_out; // @[RegFile.scala 66:20:@40248.4]
  wire  regs_428_io_enable; // @[RegFile.scala 66:20:@40248.4]
  wire  regs_429_clock; // @[RegFile.scala 66:20:@40262.4]
  wire  regs_429_reset; // @[RegFile.scala 66:20:@40262.4]
  wire [63:0] regs_429_io_in; // @[RegFile.scala 66:20:@40262.4]
  wire  regs_429_io_reset; // @[RegFile.scala 66:20:@40262.4]
  wire [63:0] regs_429_io_out; // @[RegFile.scala 66:20:@40262.4]
  wire  regs_429_io_enable; // @[RegFile.scala 66:20:@40262.4]
  wire  regs_430_clock; // @[RegFile.scala 66:20:@40276.4]
  wire  regs_430_reset; // @[RegFile.scala 66:20:@40276.4]
  wire [63:0] regs_430_io_in; // @[RegFile.scala 66:20:@40276.4]
  wire  regs_430_io_reset; // @[RegFile.scala 66:20:@40276.4]
  wire [63:0] regs_430_io_out; // @[RegFile.scala 66:20:@40276.4]
  wire  regs_430_io_enable; // @[RegFile.scala 66:20:@40276.4]
  wire  regs_431_clock; // @[RegFile.scala 66:20:@40290.4]
  wire  regs_431_reset; // @[RegFile.scala 66:20:@40290.4]
  wire [63:0] regs_431_io_in; // @[RegFile.scala 66:20:@40290.4]
  wire  regs_431_io_reset; // @[RegFile.scala 66:20:@40290.4]
  wire [63:0] regs_431_io_out; // @[RegFile.scala 66:20:@40290.4]
  wire  regs_431_io_enable; // @[RegFile.scala 66:20:@40290.4]
  wire  regs_432_clock; // @[RegFile.scala 66:20:@40304.4]
  wire  regs_432_reset; // @[RegFile.scala 66:20:@40304.4]
  wire [63:0] regs_432_io_in; // @[RegFile.scala 66:20:@40304.4]
  wire  regs_432_io_reset; // @[RegFile.scala 66:20:@40304.4]
  wire [63:0] regs_432_io_out; // @[RegFile.scala 66:20:@40304.4]
  wire  regs_432_io_enable; // @[RegFile.scala 66:20:@40304.4]
  wire  regs_433_clock; // @[RegFile.scala 66:20:@40318.4]
  wire  regs_433_reset; // @[RegFile.scala 66:20:@40318.4]
  wire [63:0] regs_433_io_in; // @[RegFile.scala 66:20:@40318.4]
  wire  regs_433_io_reset; // @[RegFile.scala 66:20:@40318.4]
  wire [63:0] regs_433_io_out; // @[RegFile.scala 66:20:@40318.4]
  wire  regs_433_io_enable; // @[RegFile.scala 66:20:@40318.4]
  wire  regs_434_clock; // @[RegFile.scala 66:20:@40332.4]
  wire  regs_434_reset; // @[RegFile.scala 66:20:@40332.4]
  wire [63:0] regs_434_io_in; // @[RegFile.scala 66:20:@40332.4]
  wire  regs_434_io_reset; // @[RegFile.scala 66:20:@40332.4]
  wire [63:0] regs_434_io_out; // @[RegFile.scala 66:20:@40332.4]
  wire  regs_434_io_enable; // @[RegFile.scala 66:20:@40332.4]
  wire  regs_435_clock; // @[RegFile.scala 66:20:@40346.4]
  wire  regs_435_reset; // @[RegFile.scala 66:20:@40346.4]
  wire [63:0] regs_435_io_in; // @[RegFile.scala 66:20:@40346.4]
  wire  regs_435_io_reset; // @[RegFile.scala 66:20:@40346.4]
  wire [63:0] regs_435_io_out; // @[RegFile.scala 66:20:@40346.4]
  wire  regs_435_io_enable; // @[RegFile.scala 66:20:@40346.4]
  wire  regs_436_clock; // @[RegFile.scala 66:20:@40360.4]
  wire  regs_436_reset; // @[RegFile.scala 66:20:@40360.4]
  wire [63:0] regs_436_io_in; // @[RegFile.scala 66:20:@40360.4]
  wire  regs_436_io_reset; // @[RegFile.scala 66:20:@40360.4]
  wire [63:0] regs_436_io_out; // @[RegFile.scala 66:20:@40360.4]
  wire  regs_436_io_enable; // @[RegFile.scala 66:20:@40360.4]
  wire  regs_437_clock; // @[RegFile.scala 66:20:@40374.4]
  wire  regs_437_reset; // @[RegFile.scala 66:20:@40374.4]
  wire [63:0] regs_437_io_in; // @[RegFile.scala 66:20:@40374.4]
  wire  regs_437_io_reset; // @[RegFile.scala 66:20:@40374.4]
  wire [63:0] regs_437_io_out; // @[RegFile.scala 66:20:@40374.4]
  wire  regs_437_io_enable; // @[RegFile.scala 66:20:@40374.4]
  wire  regs_438_clock; // @[RegFile.scala 66:20:@40388.4]
  wire  regs_438_reset; // @[RegFile.scala 66:20:@40388.4]
  wire [63:0] regs_438_io_in; // @[RegFile.scala 66:20:@40388.4]
  wire  regs_438_io_reset; // @[RegFile.scala 66:20:@40388.4]
  wire [63:0] regs_438_io_out; // @[RegFile.scala 66:20:@40388.4]
  wire  regs_438_io_enable; // @[RegFile.scala 66:20:@40388.4]
  wire  regs_439_clock; // @[RegFile.scala 66:20:@40402.4]
  wire  regs_439_reset; // @[RegFile.scala 66:20:@40402.4]
  wire [63:0] regs_439_io_in; // @[RegFile.scala 66:20:@40402.4]
  wire  regs_439_io_reset; // @[RegFile.scala 66:20:@40402.4]
  wire [63:0] regs_439_io_out; // @[RegFile.scala 66:20:@40402.4]
  wire  regs_439_io_enable; // @[RegFile.scala 66:20:@40402.4]
  wire  regs_440_clock; // @[RegFile.scala 66:20:@40416.4]
  wire  regs_440_reset; // @[RegFile.scala 66:20:@40416.4]
  wire [63:0] regs_440_io_in; // @[RegFile.scala 66:20:@40416.4]
  wire  regs_440_io_reset; // @[RegFile.scala 66:20:@40416.4]
  wire [63:0] regs_440_io_out; // @[RegFile.scala 66:20:@40416.4]
  wire  regs_440_io_enable; // @[RegFile.scala 66:20:@40416.4]
  wire  regs_441_clock; // @[RegFile.scala 66:20:@40430.4]
  wire  regs_441_reset; // @[RegFile.scala 66:20:@40430.4]
  wire [63:0] regs_441_io_in; // @[RegFile.scala 66:20:@40430.4]
  wire  regs_441_io_reset; // @[RegFile.scala 66:20:@40430.4]
  wire [63:0] regs_441_io_out; // @[RegFile.scala 66:20:@40430.4]
  wire  regs_441_io_enable; // @[RegFile.scala 66:20:@40430.4]
  wire  regs_442_clock; // @[RegFile.scala 66:20:@40444.4]
  wire  regs_442_reset; // @[RegFile.scala 66:20:@40444.4]
  wire [63:0] regs_442_io_in; // @[RegFile.scala 66:20:@40444.4]
  wire  regs_442_io_reset; // @[RegFile.scala 66:20:@40444.4]
  wire [63:0] regs_442_io_out; // @[RegFile.scala 66:20:@40444.4]
  wire  regs_442_io_enable; // @[RegFile.scala 66:20:@40444.4]
  wire  regs_443_clock; // @[RegFile.scala 66:20:@40458.4]
  wire  regs_443_reset; // @[RegFile.scala 66:20:@40458.4]
  wire [63:0] regs_443_io_in; // @[RegFile.scala 66:20:@40458.4]
  wire  regs_443_io_reset; // @[RegFile.scala 66:20:@40458.4]
  wire [63:0] regs_443_io_out; // @[RegFile.scala 66:20:@40458.4]
  wire  regs_443_io_enable; // @[RegFile.scala 66:20:@40458.4]
  wire  regs_444_clock; // @[RegFile.scala 66:20:@40472.4]
  wire  regs_444_reset; // @[RegFile.scala 66:20:@40472.4]
  wire [63:0] regs_444_io_in; // @[RegFile.scala 66:20:@40472.4]
  wire  regs_444_io_reset; // @[RegFile.scala 66:20:@40472.4]
  wire [63:0] regs_444_io_out; // @[RegFile.scala 66:20:@40472.4]
  wire  regs_444_io_enable; // @[RegFile.scala 66:20:@40472.4]
  wire  regs_445_clock; // @[RegFile.scala 66:20:@40486.4]
  wire  regs_445_reset; // @[RegFile.scala 66:20:@40486.4]
  wire [63:0] regs_445_io_in; // @[RegFile.scala 66:20:@40486.4]
  wire  regs_445_io_reset; // @[RegFile.scala 66:20:@40486.4]
  wire [63:0] regs_445_io_out; // @[RegFile.scala 66:20:@40486.4]
  wire  regs_445_io_enable; // @[RegFile.scala 66:20:@40486.4]
  wire  regs_446_clock; // @[RegFile.scala 66:20:@40500.4]
  wire  regs_446_reset; // @[RegFile.scala 66:20:@40500.4]
  wire [63:0] regs_446_io_in; // @[RegFile.scala 66:20:@40500.4]
  wire  regs_446_io_reset; // @[RegFile.scala 66:20:@40500.4]
  wire [63:0] regs_446_io_out; // @[RegFile.scala 66:20:@40500.4]
  wire  regs_446_io_enable; // @[RegFile.scala 66:20:@40500.4]
  wire  regs_447_clock; // @[RegFile.scala 66:20:@40514.4]
  wire  regs_447_reset; // @[RegFile.scala 66:20:@40514.4]
  wire [63:0] regs_447_io_in; // @[RegFile.scala 66:20:@40514.4]
  wire  regs_447_io_reset; // @[RegFile.scala 66:20:@40514.4]
  wire [63:0] regs_447_io_out; // @[RegFile.scala 66:20:@40514.4]
  wire  regs_447_io_enable; // @[RegFile.scala 66:20:@40514.4]
  wire  regs_448_clock; // @[RegFile.scala 66:20:@40528.4]
  wire  regs_448_reset; // @[RegFile.scala 66:20:@40528.4]
  wire [63:0] regs_448_io_in; // @[RegFile.scala 66:20:@40528.4]
  wire  regs_448_io_reset; // @[RegFile.scala 66:20:@40528.4]
  wire [63:0] regs_448_io_out; // @[RegFile.scala 66:20:@40528.4]
  wire  regs_448_io_enable; // @[RegFile.scala 66:20:@40528.4]
  wire  regs_449_clock; // @[RegFile.scala 66:20:@40542.4]
  wire  regs_449_reset; // @[RegFile.scala 66:20:@40542.4]
  wire [63:0] regs_449_io_in; // @[RegFile.scala 66:20:@40542.4]
  wire  regs_449_io_reset; // @[RegFile.scala 66:20:@40542.4]
  wire [63:0] regs_449_io_out; // @[RegFile.scala 66:20:@40542.4]
  wire  regs_449_io_enable; // @[RegFile.scala 66:20:@40542.4]
  wire  regs_450_clock; // @[RegFile.scala 66:20:@40556.4]
  wire  regs_450_reset; // @[RegFile.scala 66:20:@40556.4]
  wire [63:0] regs_450_io_in; // @[RegFile.scala 66:20:@40556.4]
  wire  regs_450_io_reset; // @[RegFile.scala 66:20:@40556.4]
  wire [63:0] regs_450_io_out; // @[RegFile.scala 66:20:@40556.4]
  wire  regs_450_io_enable; // @[RegFile.scala 66:20:@40556.4]
  wire  regs_451_clock; // @[RegFile.scala 66:20:@40570.4]
  wire  regs_451_reset; // @[RegFile.scala 66:20:@40570.4]
  wire [63:0] regs_451_io_in; // @[RegFile.scala 66:20:@40570.4]
  wire  regs_451_io_reset; // @[RegFile.scala 66:20:@40570.4]
  wire [63:0] regs_451_io_out; // @[RegFile.scala 66:20:@40570.4]
  wire  regs_451_io_enable; // @[RegFile.scala 66:20:@40570.4]
  wire  regs_452_clock; // @[RegFile.scala 66:20:@40584.4]
  wire  regs_452_reset; // @[RegFile.scala 66:20:@40584.4]
  wire [63:0] regs_452_io_in; // @[RegFile.scala 66:20:@40584.4]
  wire  regs_452_io_reset; // @[RegFile.scala 66:20:@40584.4]
  wire [63:0] regs_452_io_out; // @[RegFile.scala 66:20:@40584.4]
  wire  regs_452_io_enable; // @[RegFile.scala 66:20:@40584.4]
  wire  regs_453_clock; // @[RegFile.scala 66:20:@40598.4]
  wire  regs_453_reset; // @[RegFile.scala 66:20:@40598.4]
  wire [63:0] regs_453_io_in; // @[RegFile.scala 66:20:@40598.4]
  wire  regs_453_io_reset; // @[RegFile.scala 66:20:@40598.4]
  wire [63:0] regs_453_io_out; // @[RegFile.scala 66:20:@40598.4]
  wire  regs_453_io_enable; // @[RegFile.scala 66:20:@40598.4]
  wire  regs_454_clock; // @[RegFile.scala 66:20:@40612.4]
  wire  regs_454_reset; // @[RegFile.scala 66:20:@40612.4]
  wire [63:0] regs_454_io_in; // @[RegFile.scala 66:20:@40612.4]
  wire  regs_454_io_reset; // @[RegFile.scala 66:20:@40612.4]
  wire [63:0] regs_454_io_out; // @[RegFile.scala 66:20:@40612.4]
  wire  regs_454_io_enable; // @[RegFile.scala 66:20:@40612.4]
  wire  regs_455_clock; // @[RegFile.scala 66:20:@40626.4]
  wire  regs_455_reset; // @[RegFile.scala 66:20:@40626.4]
  wire [63:0] regs_455_io_in; // @[RegFile.scala 66:20:@40626.4]
  wire  regs_455_io_reset; // @[RegFile.scala 66:20:@40626.4]
  wire [63:0] regs_455_io_out; // @[RegFile.scala 66:20:@40626.4]
  wire  regs_455_io_enable; // @[RegFile.scala 66:20:@40626.4]
  wire  regs_456_clock; // @[RegFile.scala 66:20:@40640.4]
  wire  regs_456_reset; // @[RegFile.scala 66:20:@40640.4]
  wire [63:0] regs_456_io_in; // @[RegFile.scala 66:20:@40640.4]
  wire  regs_456_io_reset; // @[RegFile.scala 66:20:@40640.4]
  wire [63:0] regs_456_io_out; // @[RegFile.scala 66:20:@40640.4]
  wire  regs_456_io_enable; // @[RegFile.scala 66:20:@40640.4]
  wire  regs_457_clock; // @[RegFile.scala 66:20:@40654.4]
  wire  regs_457_reset; // @[RegFile.scala 66:20:@40654.4]
  wire [63:0] regs_457_io_in; // @[RegFile.scala 66:20:@40654.4]
  wire  regs_457_io_reset; // @[RegFile.scala 66:20:@40654.4]
  wire [63:0] regs_457_io_out; // @[RegFile.scala 66:20:@40654.4]
  wire  regs_457_io_enable; // @[RegFile.scala 66:20:@40654.4]
  wire  regs_458_clock; // @[RegFile.scala 66:20:@40668.4]
  wire  regs_458_reset; // @[RegFile.scala 66:20:@40668.4]
  wire [63:0] regs_458_io_in; // @[RegFile.scala 66:20:@40668.4]
  wire  regs_458_io_reset; // @[RegFile.scala 66:20:@40668.4]
  wire [63:0] regs_458_io_out; // @[RegFile.scala 66:20:@40668.4]
  wire  regs_458_io_enable; // @[RegFile.scala 66:20:@40668.4]
  wire  regs_459_clock; // @[RegFile.scala 66:20:@40682.4]
  wire  regs_459_reset; // @[RegFile.scala 66:20:@40682.4]
  wire [63:0] regs_459_io_in; // @[RegFile.scala 66:20:@40682.4]
  wire  regs_459_io_reset; // @[RegFile.scala 66:20:@40682.4]
  wire [63:0] regs_459_io_out; // @[RegFile.scala 66:20:@40682.4]
  wire  regs_459_io_enable; // @[RegFile.scala 66:20:@40682.4]
  wire  regs_460_clock; // @[RegFile.scala 66:20:@40696.4]
  wire  regs_460_reset; // @[RegFile.scala 66:20:@40696.4]
  wire [63:0] regs_460_io_in; // @[RegFile.scala 66:20:@40696.4]
  wire  regs_460_io_reset; // @[RegFile.scala 66:20:@40696.4]
  wire [63:0] regs_460_io_out; // @[RegFile.scala 66:20:@40696.4]
  wire  regs_460_io_enable; // @[RegFile.scala 66:20:@40696.4]
  wire  regs_461_clock; // @[RegFile.scala 66:20:@40710.4]
  wire  regs_461_reset; // @[RegFile.scala 66:20:@40710.4]
  wire [63:0] regs_461_io_in; // @[RegFile.scala 66:20:@40710.4]
  wire  regs_461_io_reset; // @[RegFile.scala 66:20:@40710.4]
  wire [63:0] regs_461_io_out; // @[RegFile.scala 66:20:@40710.4]
  wire  regs_461_io_enable; // @[RegFile.scala 66:20:@40710.4]
  wire  regs_462_clock; // @[RegFile.scala 66:20:@40724.4]
  wire  regs_462_reset; // @[RegFile.scala 66:20:@40724.4]
  wire [63:0] regs_462_io_in; // @[RegFile.scala 66:20:@40724.4]
  wire  regs_462_io_reset; // @[RegFile.scala 66:20:@40724.4]
  wire [63:0] regs_462_io_out; // @[RegFile.scala 66:20:@40724.4]
  wire  regs_462_io_enable; // @[RegFile.scala 66:20:@40724.4]
  wire  regs_463_clock; // @[RegFile.scala 66:20:@40738.4]
  wire  regs_463_reset; // @[RegFile.scala 66:20:@40738.4]
  wire [63:0] regs_463_io_in; // @[RegFile.scala 66:20:@40738.4]
  wire  regs_463_io_reset; // @[RegFile.scala 66:20:@40738.4]
  wire [63:0] regs_463_io_out; // @[RegFile.scala 66:20:@40738.4]
  wire  regs_463_io_enable; // @[RegFile.scala 66:20:@40738.4]
  wire  regs_464_clock; // @[RegFile.scala 66:20:@40752.4]
  wire  regs_464_reset; // @[RegFile.scala 66:20:@40752.4]
  wire [63:0] regs_464_io_in; // @[RegFile.scala 66:20:@40752.4]
  wire  regs_464_io_reset; // @[RegFile.scala 66:20:@40752.4]
  wire [63:0] regs_464_io_out; // @[RegFile.scala 66:20:@40752.4]
  wire  regs_464_io_enable; // @[RegFile.scala 66:20:@40752.4]
  wire  regs_465_clock; // @[RegFile.scala 66:20:@40766.4]
  wire  regs_465_reset; // @[RegFile.scala 66:20:@40766.4]
  wire [63:0] regs_465_io_in; // @[RegFile.scala 66:20:@40766.4]
  wire  regs_465_io_reset; // @[RegFile.scala 66:20:@40766.4]
  wire [63:0] regs_465_io_out; // @[RegFile.scala 66:20:@40766.4]
  wire  regs_465_io_enable; // @[RegFile.scala 66:20:@40766.4]
  wire  regs_466_clock; // @[RegFile.scala 66:20:@40780.4]
  wire  regs_466_reset; // @[RegFile.scala 66:20:@40780.4]
  wire [63:0] regs_466_io_in; // @[RegFile.scala 66:20:@40780.4]
  wire  regs_466_io_reset; // @[RegFile.scala 66:20:@40780.4]
  wire [63:0] regs_466_io_out; // @[RegFile.scala 66:20:@40780.4]
  wire  regs_466_io_enable; // @[RegFile.scala 66:20:@40780.4]
  wire  regs_467_clock; // @[RegFile.scala 66:20:@40794.4]
  wire  regs_467_reset; // @[RegFile.scala 66:20:@40794.4]
  wire [63:0] regs_467_io_in; // @[RegFile.scala 66:20:@40794.4]
  wire  regs_467_io_reset; // @[RegFile.scala 66:20:@40794.4]
  wire [63:0] regs_467_io_out; // @[RegFile.scala 66:20:@40794.4]
  wire  regs_467_io_enable; // @[RegFile.scala 66:20:@40794.4]
  wire  regs_468_clock; // @[RegFile.scala 66:20:@40808.4]
  wire  regs_468_reset; // @[RegFile.scala 66:20:@40808.4]
  wire [63:0] regs_468_io_in; // @[RegFile.scala 66:20:@40808.4]
  wire  regs_468_io_reset; // @[RegFile.scala 66:20:@40808.4]
  wire [63:0] regs_468_io_out; // @[RegFile.scala 66:20:@40808.4]
  wire  regs_468_io_enable; // @[RegFile.scala 66:20:@40808.4]
  wire  regs_469_clock; // @[RegFile.scala 66:20:@40822.4]
  wire  regs_469_reset; // @[RegFile.scala 66:20:@40822.4]
  wire [63:0] regs_469_io_in; // @[RegFile.scala 66:20:@40822.4]
  wire  regs_469_io_reset; // @[RegFile.scala 66:20:@40822.4]
  wire [63:0] regs_469_io_out; // @[RegFile.scala 66:20:@40822.4]
  wire  regs_469_io_enable; // @[RegFile.scala 66:20:@40822.4]
  wire  regs_470_clock; // @[RegFile.scala 66:20:@40836.4]
  wire  regs_470_reset; // @[RegFile.scala 66:20:@40836.4]
  wire [63:0] regs_470_io_in; // @[RegFile.scala 66:20:@40836.4]
  wire  regs_470_io_reset; // @[RegFile.scala 66:20:@40836.4]
  wire [63:0] regs_470_io_out; // @[RegFile.scala 66:20:@40836.4]
  wire  regs_470_io_enable; // @[RegFile.scala 66:20:@40836.4]
  wire  regs_471_clock; // @[RegFile.scala 66:20:@40850.4]
  wire  regs_471_reset; // @[RegFile.scala 66:20:@40850.4]
  wire [63:0] regs_471_io_in; // @[RegFile.scala 66:20:@40850.4]
  wire  regs_471_io_reset; // @[RegFile.scala 66:20:@40850.4]
  wire [63:0] regs_471_io_out; // @[RegFile.scala 66:20:@40850.4]
  wire  regs_471_io_enable; // @[RegFile.scala 66:20:@40850.4]
  wire  regs_472_clock; // @[RegFile.scala 66:20:@40864.4]
  wire  regs_472_reset; // @[RegFile.scala 66:20:@40864.4]
  wire [63:0] regs_472_io_in; // @[RegFile.scala 66:20:@40864.4]
  wire  regs_472_io_reset; // @[RegFile.scala 66:20:@40864.4]
  wire [63:0] regs_472_io_out; // @[RegFile.scala 66:20:@40864.4]
  wire  regs_472_io_enable; // @[RegFile.scala 66:20:@40864.4]
  wire  regs_473_clock; // @[RegFile.scala 66:20:@40878.4]
  wire  regs_473_reset; // @[RegFile.scala 66:20:@40878.4]
  wire [63:0] regs_473_io_in; // @[RegFile.scala 66:20:@40878.4]
  wire  regs_473_io_reset; // @[RegFile.scala 66:20:@40878.4]
  wire [63:0] regs_473_io_out; // @[RegFile.scala 66:20:@40878.4]
  wire  regs_473_io_enable; // @[RegFile.scala 66:20:@40878.4]
  wire  regs_474_clock; // @[RegFile.scala 66:20:@40892.4]
  wire  regs_474_reset; // @[RegFile.scala 66:20:@40892.4]
  wire [63:0] regs_474_io_in; // @[RegFile.scala 66:20:@40892.4]
  wire  regs_474_io_reset; // @[RegFile.scala 66:20:@40892.4]
  wire [63:0] regs_474_io_out; // @[RegFile.scala 66:20:@40892.4]
  wire  regs_474_io_enable; // @[RegFile.scala 66:20:@40892.4]
  wire  regs_475_clock; // @[RegFile.scala 66:20:@40906.4]
  wire  regs_475_reset; // @[RegFile.scala 66:20:@40906.4]
  wire [63:0] regs_475_io_in; // @[RegFile.scala 66:20:@40906.4]
  wire  regs_475_io_reset; // @[RegFile.scala 66:20:@40906.4]
  wire [63:0] regs_475_io_out; // @[RegFile.scala 66:20:@40906.4]
  wire  regs_475_io_enable; // @[RegFile.scala 66:20:@40906.4]
  wire  regs_476_clock; // @[RegFile.scala 66:20:@40920.4]
  wire  regs_476_reset; // @[RegFile.scala 66:20:@40920.4]
  wire [63:0] regs_476_io_in; // @[RegFile.scala 66:20:@40920.4]
  wire  regs_476_io_reset; // @[RegFile.scala 66:20:@40920.4]
  wire [63:0] regs_476_io_out; // @[RegFile.scala 66:20:@40920.4]
  wire  regs_476_io_enable; // @[RegFile.scala 66:20:@40920.4]
  wire  regs_477_clock; // @[RegFile.scala 66:20:@40934.4]
  wire  regs_477_reset; // @[RegFile.scala 66:20:@40934.4]
  wire [63:0] regs_477_io_in; // @[RegFile.scala 66:20:@40934.4]
  wire  regs_477_io_reset; // @[RegFile.scala 66:20:@40934.4]
  wire [63:0] regs_477_io_out; // @[RegFile.scala 66:20:@40934.4]
  wire  regs_477_io_enable; // @[RegFile.scala 66:20:@40934.4]
  wire  regs_478_clock; // @[RegFile.scala 66:20:@40948.4]
  wire  regs_478_reset; // @[RegFile.scala 66:20:@40948.4]
  wire [63:0] regs_478_io_in; // @[RegFile.scala 66:20:@40948.4]
  wire  regs_478_io_reset; // @[RegFile.scala 66:20:@40948.4]
  wire [63:0] regs_478_io_out; // @[RegFile.scala 66:20:@40948.4]
  wire  regs_478_io_enable; // @[RegFile.scala 66:20:@40948.4]
  wire  regs_479_clock; // @[RegFile.scala 66:20:@40962.4]
  wire  regs_479_reset; // @[RegFile.scala 66:20:@40962.4]
  wire [63:0] regs_479_io_in; // @[RegFile.scala 66:20:@40962.4]
  wire  regs_479_io_reset; // @[RegFile.scala 66:20:@40962.4]
  wire [63:0] regs_479_io_out; // @[RegFile.scala 66:20:@40962.4]
  wire  regs_479_io_enable; // @[RegFile.scala 66:20:@40962.4]
  wire  regs_480_clock; // @[RegFile.scala 66:20:@40976.4]
  wire  regs_480_reset; // @[RegFile.scala 66:20:@40976.4]
  wire [63:0] regs_480_io_in; // @[RegFile.scala 66:20:@40976.4]
  wire  regs_480_io_reset; // @[RegFile.scala 66:20:@40976.4]
  wire [63:0] regs_480_io_out; // @[RegFile.scala 66:20:@40976.4]
  wire  regs_480_io_enable; // @[RegFile.scala 66:20:@40976.4]
  wire  regs_481_clock; // @[RegFile.scala 66:20:@40990.4]
  wire  regs_481_reset; // @[RegFile.scala 66:20:@40990.4]
  wire [63:0] regs_481_io_in; // @[RegFile.scala 66:20:@40990.4]
  wire  regs_481_io_reset; // @[RegFile.scala 66:20:@40990.4]
  wire [63:0] regs_481_io_out; // @[RegFile.scala 66:20:@40990.4]
  wire  regs_481_io_enable; // @[RegFile.scala 66:20:@40990.4]
  wire  regs_482_clock; // @[RegFile.scala 66:20:@41004.4]
  wire  regs_482_reset; // @[RegFile.scala 66:20:@41004.4]
  wire [63:0] regs_482_io_in; // @[RegFile.scala 66:20:@41004.4]
  wire  regs_482_io_reset; // @[RegFile.scala 66:20:@41004.4]
  wire [63:0] regs_482_io_out; // @[RegFile.scala 66:20:@41004.4]
  wire  regs_482_io_enable; // @[RegFile.scala 66:20:@41004.4]
  wire  regs_483_clock; // @[RegFile.scala 66:20:@41018.4]
  wire  regs_483_reset; // @[RegFile.scala 66:20:@41018.4]
  wire [63:0] regs_483_io_in; // @[RegFile.scala 66:20:@41018.4]
  wire  regs_483_io_reset; // @[RegFile.scala 66:20:@41018.4]
  wire [63:0] regs_483_io_out; // @[RegFile.scala 66:20:@41018.4]
  wire  regs_483_io_enable; // @[RegFile.scala 66:20:@41018.4]
  wire  regs_484_clock; // @[RegFile.scala 66:20:@41032.4]
  wire  regs_484_reset; // @[RegFile.scala 66:20:@41032.4]
  wire [63:0] regs_484_io_in; // @[RegFile.scala 66:20:@41032.4]
  wire  regs_484_io_reset; // @[RegFile.scala 66:20:@41032.4]
  wire [63:0] regs_484_io_out; // @[RegFile.scala 66:20:@41032.4]
  wire  regs_484_io_enable; // @[RegFile.scala 66:20:@41032.4]
  wire  regs_485_clock; // @[RegFile.scala 66:20:@41046.4]
  wire  regs_485_reset; // @[RegFile.scala 66:20:@41046.4]
  wire [63:0] regs_485_io_in; // @[RegFile.scala 66:20:@41046.4]
  wire  regs_485_io_reset; // @[RegFile.scala 66:20:@41046.4]
  wire [63:0] regs_485_io_out; // @[RegFile.scala 66:20:@41046.4]
  wire  regs_485_io_enable; // @[RegFile.scala 66:20:@41046.4]
  wire  regs_486_clock; // @[RegFile.scala 66:20:@41060.4]
  wire  regs_486_reset; // @[RegFile.scala 66:20:@41060.4]
  wire [63:0] regs_486_io_in; // @[RegFile.scala 66:20:@41060.4]
  wire  regs_486_io_reset; // @[RegFile.scala 66:20:@41060.4]
  wire [63:0] regs_486_io_out; // @[RegFile.scala 66:20:@41060.4]
  wire  regs_486_io_enable; // @[RegFile.scala 66:20:@41060.4]
  wire  regs_487_clock; // @[RegFile.scala 66:20:@41074.4]
  wire  regs_487_reset; // @[RegFile.scala 66:20:@41074.4]
  wire [63:0] regs_487_io_in; // @[RegFile.scala 66:20:@41074.4]
  wire  regs_487_io_reset; // @[RegFile.scala 66:20:@41074.4]
  wire [63:0] regs_487_io_out; // @[RegFile.scala 66:20:@41074.4]
  wire  regs_487_io_enable; // @[RegFile.scala 66:20:@41074.4]
  wire  regs_488_clock; // @[RegFile.scala 66:20:@41088.4]
  wire  regs_488_reset; // @[RegFile.scala 66:20:@41088.4]
  wire [63:0] regs_488_io_in; // @[RegFile.scala 66:20:@41088.4]
  wire  regs_488_io_reset; // @[RegFile.scala 66:20:@41088.4]
  wire [63:0] regs_488_io_out; // @[RegFile.scala 66:20:@41088.4]
  wire  regs_488_io_enable; // @[RegFile.scala 66:20:@41088.4]
  wire  regs_489_clock; // @[RegFile.scala 66:20:@41102.4]
  wire  regs_489_reset; // @[RegFile.scala 66:20:@41102.4]
  wire [63:0] regs_489_io_in; // @[RegFile.scala 66:20:@41102.4]
  wire  regs_489_io_reset; // @[RegFile.scala 66:20:@41102.4]
  wire [63:0] regs_489_io_out; // @[RegFile.scala 66:20:@41102.4]
  wire  regs_489_io_enable; // @[RegFile.scala 66:20:@41102.4]
  wire  regs_490_clock; // @[RegFile.scala 66:20:@41116.4]
  wire  regs_490_reset; // @[RegFile.scala 66:20:@41116.4]
  wire [63:0] regs_490_io_in; // @[RegFile.scala 66:20:@41116.4]
  wire  regs_490_io_reset; // @[RegFile.scala 66:20:@41116.4]
  wire [63:0] regs_490_io_out; // @[RegFile.scala 66:20:@41116.4]
  wire  regs_490_io_enable; // @[RegFile.scala 66:20:@41116.4]
  wire  regs_491_clock; // @[RegFile.scala 66:20:@41130.4]
  wire  regs_491_reset; // @[RegFile.scala 66:20:@41130.4]
  wire [63:0] regs_491_io_in; // @[RegFile.scala 66:20:@41130.4]
  wire  regs_491_io_reset; // @[RegFile.scala 66:20:@41130.4]
  wire [63:0] regs_491_io_out; // @[RegFile.scala 66:20:@41130.4]
  wire  regs_491_io_enable; // @[RegFile.scala 66:20:@41130.4]
  wire  regs_492_clock; // @[RegFile.scala 66:20:@41144.4]
  wire  regs_492_reset; // @[RegFile.scala 66:20:@41144.4]
  wire [63:0] regs_492_io_in; // @[RegFile.scala 66:20:@41144.4]
  wire  regs_492_io_reset; // @[RegFile.scala 66:20:@41144.4]
  wire [63:0] regs_492_io_out; // @[RegFile.scala 66:20:@41144.4]
  wire  regs_492_io_enable; // @[RegFile.scala 66:20:@41144.4]
  wire  regs_493_clock; // @[RegFile.scala 66:20:@41158.4]
  wire  regs_493_reset; // @[RegFile.scala 66:20:@41158.4]
  wire [63:0] regs_493_io_in; // @[RegFile.scala 66:20:@41158.4]
  wire  regs_493_io_reset; // @[RegFile.scala 66:20:@41158.4]
  wire [63:0] regs_493_io_out; // @[RegFile.scala 66:20:@41158.4]
  wire  regs_493_io_enable; // @[RegFile.scala 66:20:@41158.4]
  wire  regs_494_clock; // @[RegFile.scala 66:20:@41172.4]
  wire  regs_494_reset; // @[RegFile.scala 66:20:@41172.4]
  wire [63:0] regs_494_io_in; // @[RegFile.scala 66:20:@41172.4]
  wire  regs_494_io_reset; // @[RegFile.scala 66:20:@41172.4]
  wire [63:0] regs_494_io_out; // @[RegFile.scala 66:20:@41172.4]
  wire  regs_494_io_enable; // @[RegFile.scala 66:20:@41172.4]
  wire  regs_495_clock; // @[RegFile.scala 66:20:@41186.4]
  wire  regs_495_reset; // @[RegFile.scala 66:20:@41186.4]
  wire [63:0] regs_495_io_in; // @[RegFile.scala 66:20:@41186.4]
  wire  regs_495_io_reset; // @[RegFile.scala 66:20:@41186.4]
  wire [63:0] regs_495_io_out; // @[RegFile.scala 66:20:@41186.4]
  wire  regs_495_io_enable; // @[RegFile.scala 66:20:@41186.4]
  wire  regs_496_clock; // @[RegFile.scala 66:20:@41200.4]
  wire  regs_496_reset; // @[RegFile.scala 66:20:@41200.4]
  wire [63:0] regs_496_io_in; // @[RegFile.scala 66:20:@41200.4]
  wire  regs_496_io_reset; // @[RegFile.scala 66:20:@41200.4]
  wire [63:0] regs_496_io_out; // @[RegFile.scala 66:20:@41200.4]
  wire  regs_496_io_enable; // @[RegFile.scala 66:20:@41200.4]
  wire  regs_497_clock; // @[RegFile.scala 66:20:@41214.4]
  wire  regs_497_reset; // @[RegFile.scala 66:20:@41214.4]
  wire [63:0] regs_497_io_in; // @[RegFile.scala 66:20:@41214.4]
  wire  regs_497_io_reset; // @[RegFile.scala 66:20:@41214.4]
  wire [63:0] regs_497_io_out; // @[RegFile.scala 66:20:@41214.4]
  wire  regs_497_io_enable; // @[RegFile.scala 66:20:@41214.4]
  wire  regs_498_clock; // @[RegFile.scala 66:20:@41228.4]
  wire  regs_498_reset; // @[RegFile.scala 66:20:@41228.4]
  wire [63:0] regs_498_io_in; // @[RegFile.scala 66:20:@41228.4]
  wire  regs_498_io_reset; // @[RegFile.scala 66:20:@41228.4]
  wire [63:0] regs_498_io_out; // @[RegFile.scala 66:20:@41228.4]
  wire  regs_498_io_enable; // @[RegFile.scala 66:20:@41228.4]
  wire  regs_499_clock; // @[RegFile.scala 66:20:@41242.4]
  wire  regs_499_reset; // @[RegFile.scala 66:20:@41242.4]
  wire [63:0] regs_499_io_in; // @[RegFile.scala 66:20:@41242.4]
  wire  regs_499_io_reset; // @[RegFile.scala 66:20:@41242.4]
  wire [63:0] regs_499_io_out; // @[RegFile.scala 66:20:@41242.4]
  wire  regs_499_io_enable; // @[RegFile.scala 66:20:@41242.4]
  wire  regs_500_clock; // @[RegFile.scala 66:20:@41256.4]
  wire  regs_500_reset; // @[RegFile.scala 66:20:@41256.4]
  wire [63:0] regs_500_io_in; // @[RegFile.scala 66:20:@41256.4]
  wire  regs_500_io_reset; // @[RegFile.scala 66:20:@41256.4]
  wire [63:0] regs_500_io_out; // @[RegFile.scala 66:20:@41256.4]
  wire  regs_500_io_enable; // @[RegFile.scala 66:20:@41256.4]
  wire  regs_501_clock; // @[RegFile.scala 66:20:@41270.4]
  wire  regs_501_reset; // @[RegFile.scala 66:20:@41270.4]
  wire [63:0] regs_501_io_in; // @[RegFile.scala 66:20:@41270.4]
  wire  regs_501_io_reset; // @[RegFile.scala 66:20:@41270.4]
  wire [63:0] regs_501_io_out; // @[RegFile.scala 66:20:@41270.4]
  wire  regs_501_io_enable; // @[RegFile.scala 66:20:@41270.4]
  wire  regs_502_clock; // @[RegFile.scala 66:20:@41284.4]
  wire  regs_502_reset; // @[RegFile.scala 66:20:@41284.4]
  wire [63:0] regs_502_io_in; // @[RegFile.scala 66:20:@41284.4]
  wire  regs_502_io_reset; // @[RegFile.scala 66:20:@41284.4]
  wire [63:0] regs_502_io_out; // @[RegFile.scala 66:20:@41284.4]
  wire  regs_502_io_enable; // @[RegFile.scala 66:20:@41284.4]
  wire [63:0] rport_io_ins_0; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_1; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_2; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_3; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_4; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_5; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_6; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_7; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_8; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_9; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_10; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_11; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_12; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_13; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_14; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_15; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_16; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_17; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_18; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_19; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_20; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_21; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_22; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_23; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_24; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_25; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_26; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_27; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_28; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_29; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_30; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_31; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_32; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_33; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_34; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_35; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_36; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_37; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_38; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_39; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_40; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_41; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_42; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_43; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_44; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_45; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_46; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_47; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_48; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_49; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_50; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_51; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_52; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_53; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_54; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_55; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_56; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_57; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_58; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_59; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_60; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_61; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_62; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_63; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_64; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_65; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_66; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_67; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_68; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_69; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_70; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_71; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_72; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_73; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_74; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_75; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_76; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_77; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_78; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_79; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_80; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_81; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_82; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_83; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_84; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_85; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_86; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_87; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_88; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_89; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_90; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_91; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_92; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_93; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_94; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_95; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_96; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_97; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_98; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_99; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_100; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_101; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_102; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_103; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_104; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_105; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_106; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_107; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_108; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_109; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_110; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_111; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_112; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_113; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_114; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_115; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_116; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_117; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_118; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_119; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_120; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_121; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_122; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_123; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_124; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_125; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_126; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_127; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_128; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_129; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_130; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_131; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_132; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_133; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_134; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_135; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_136; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_137; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_138; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_139; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_140; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_141; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_142; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_143; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_144; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_145; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_146; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_147; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_148; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_149; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_150; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_151; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_152; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_153; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_154; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_155; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_156; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_157; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_158; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_159; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_160; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_161; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_162; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_163; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_164; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_165; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_166; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_167; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_168; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_169; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_170; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_171; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_172; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_173; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_174; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_175; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_176; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_177; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_178; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_179; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_180; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_181; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_182; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_183; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_184; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_185; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_186; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_187; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_188; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_189; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_190; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_191; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_192; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_193; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_194; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_195; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_196; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_197; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_198; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_199; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_200; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_201; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_202; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_203; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_204; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_205; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_206; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_207; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_208; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_209; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_210; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_211; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_212; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_213; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_214; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_215; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_216; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_217; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_218; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_219; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_220; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_221; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_222; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_223; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_224; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_225; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_226; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_227; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_228; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_229; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_230; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_231; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_232; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_233; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_234; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_235; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_236; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_237; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_238; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_239; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_240; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_241; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_242; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_243; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_244; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_245; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_246; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_247; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_248; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_249; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_250; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_251; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_252; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_253; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_254; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_255; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_256; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_257; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_258; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_259; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_260; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_261; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_262; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_263; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_264; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_265; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_266; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_267; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_268; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_269; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_270; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_271; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_272; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_273; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_274; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_275; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_276; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_277; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_278; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_279; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_280; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_281; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_282; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_283; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_284; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_285; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_286; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_287; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_288; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_289; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_290; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_291; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_292; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_293; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_294; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_295; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_296; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_297; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_298; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_299; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_300; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_301; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_302; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_303; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_304; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_305; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_306; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_307; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_308; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_309; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_310; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_311; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_312; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_313; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_314; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_315; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_316; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_317; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_318; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_319; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_320; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_321; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_322; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_323; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_324; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_325; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_326; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_327; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_328; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_329; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_330; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_331; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_332; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_333; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_334; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_335; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_336; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_337; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_338; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_339; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_340; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_341; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_342; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_343; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_344; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_345; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_346; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_347; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_348; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_349; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_350; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_351; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_352; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_353; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_354; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_355; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_356; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_357; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_358; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_359; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_360; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_361; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_362; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_363; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_364; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_365; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_366; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_367; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_368; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_369; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_370; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_371; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_372; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_373; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_374; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_375; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_376; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_377; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_378; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_379; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_380; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_381; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_382; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_383; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_384; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_385; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_386; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_387; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_388; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_389; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_390; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_391; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_392; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_393; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_394; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_395; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_396; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_397; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_398; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_399; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_400; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_401; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_402; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_403; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_404; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_405; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_406; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_407; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_408; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_409; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_410; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_411; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_412; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_413; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_414; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_415; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_416; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_417; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_418; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_419; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_420; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_421; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_422; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_423; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_424; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_425; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_426; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_427; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_428; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_429; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_430; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_431; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_432; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_433; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_434; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_435; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_436; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_437; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_438; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_439; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_440; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_441; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_442; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_443; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_444; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_445; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_446; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_447; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_448; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_449; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_450; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_451; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_452; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_453; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_454; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_455; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_456; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_457; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_458; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_459; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_460; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_461; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_462; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_463; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_464; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_465; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_466; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_467; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_468; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_469; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_470; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_471; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_472; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_473; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_474; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_475; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_476; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_477; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_478; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_479; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_480; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_481; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_482; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_483; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_484; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_485; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_486; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_487; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_488; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_489; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_490; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_491; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_492; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_493; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_494; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_495; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_496; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_497; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_498; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_499; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_500; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_501; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_ins_502; // @[RegFile.scala 95:21:@41298.4]
  wire [8:0] rport_io_sel; // @[RegFile.scala 95:21:@41298.4]
  wire [63:0] rport_io_out; // @[RegFile.scala 95:21:@41298.4]
  wire  _T_3076; // @[RegFile.scala 80:42:@34258.4]
  wire  _T_3082; // @[RegFile.scala 68:46:@34270.4]
  wire  _T_3083; // @[RegFile.scala 68:34:@34271.4]
  wire  _T_3096; // @[RegFile.scala 80:42:@34289.4]
  wire  _T_3102; // @[RegFile.scala 74:80:@34301.4]
  wire  _T_3103; // @[RegFile.scala 74:68:@34302.4]
  FringeFF regs_0 ( // @[RegFile.scala 66:20:@34255.4]
    .clock(regs_0_clock),
    .reset(regs_0_reset),
    .io_in(regs_0_io_in),
    .io_reset(regs_0_io_reset),
    .io_out(regs_0_io_out),
    .io_enable(regs_0_io_enable)
  );
  FringeFF regs_1 ( // @[RegFile.scala 66:20:@34267.4]
    .clock(regs_1_clock),
    .reset(regs_1_reset),
    .io_in(regs_1_io_in),
    .io_reset(regs_1_io_reset),
    .io_out(regs_1_io_out),
    .io_enable(regs_1_io_enable)
  );
  FringeFF regs_2 ( // @[RegFile.scala 66:20:@34286.4]
    .clock(regs_2_clock),
    .reset(regs_2_reset),
    .io_in(regs_2_io_in),
    .io_reset(regs_2_io_reset),
    .io_out(regs_2_io_out),
    .io_enable(regs_2_io_enable)
  );
  FringeFF regs_3 ( // @[RegFile.scala 66:20:@34298.4]
    .clock(regs_3_clock),
    .reset(regs_3_reset),
    .io_in(regs_3_io_in),
    .io_reset(regs_3_io_reset),
    .io_out(regs_3_io_out),
    .io_enable(regs_3_io_enable)
  );
  FringeFF regs_4 ( // @[RegFile.scala 66:20:@34312.4]
    .clock(regs_4_clock),
    .reset(regs_4_reset),
    .io_in(regs_4_io_in),
    .io_reset(regs_4_io_reset),
    .io_out(regs_4_io_out),
    .io_enable(regs_4_io_enable)
  );
  FringeFF regs_5 ( // @[RegFile.scala 66:20:@34326.4]
    .clock(regs_5_clock),
    .reset(regs_5_reset),
    .io_in(regs_5_io_in),
    .io_reset(regs_5_io_reset),
    .io_out(regs_5_io_out),
    .io_enable(regs_5_io_enable)
  );
  FringeFF regs_6 ( // @[RegFile.scala 66:20:@34340.4]
    .clock(regs_6_clock),
    .reset(regs_6_reset),
    .io_in(regs_6_io_in),
    .io_reset(regs_6_io_reset),
    .io_out(regs_6_io_out),
    .io_enable(regs_6_io_enable)
  );
  FringeFF regs_7 ( // @[RegFile.scala 66:20:@34354.4]
    .clock(regs_7_clock),
    .reset(regs_7_reset),
    .io_in(regs_7_io_in),
    .io_reset(regs_7_io_reset),
    .io_out(regs_7_io_out),
    .io_enable(regs_7_io_enable)
  );
  FringeFF regs_8 ( // @[RegFile.scala 66:20:@34368.4]
    .clock(regs_8_clock),
    .reset(regs_8_reset),
    .io_in(regs_8_io_in),
    .io_reset(regs_8_io_reset),
    .io_out(regs_8_io_out),
    .io_enable(regs_8_io_enable)
  );
  FringeFF regs_9 ( // @[RegFile.scala 66:20:@34382.4]
    .clock(regs_9_clock),
    .reset(regs_9_reset),
    .io_in(regs_9_io_in),
    .io_reset(regs_9_io_reset),
    .io_out(regs_9_io_out),
    .io_enable(regs_9_io_enable)
  );
  FringeFF regs_10 ( // @[RegFile.scala 66:20:@34396.4]
    .clock(regs_10_clock),
    .reset(regs_10_reset),
    .io_in(regs_10_io_in),
    .io_reset(regs_10_io_reset),
    .io_out(regs_10_io_out),
    .io_enable(regs_10_io_enable)
  );
  FringeFF regs_11 ( // @[RegFile.scala 66:20:@34410.4]
    .clock(regs_11_clock),
    .reset(regs_11_reset),
    .io_in(regs_11_io_in),
    .io_reset(regs_11_io_reset),
    .io_out(regs_11_io_out),
    .io_enable(regs_11_io_enable)
  );
  FringeFF regs_12 ( // @[RegFile.scala 66:20:@34424.4]
    .clock(regs_12_clock),
    .reset(regs_12_reset),
    .io_in(regs_12_io_in),
    .io_reset(regs_12_io_reset),
    .io_out(regs_12_io_out),
    .io_enable(regs_12_io_enable)
  );
  FringeFF regs_13 ( // @[RegFile.scala 66:20:@34438.4]
    .clock(regs_13_clock),
    .reset(regs_13_reset),
    .io_in(regs_13_io_in),
    .io_reset(regs_13_io_reset),
    .io_out(regs_13_io_out),
    .io_enable(regs_13_io_enable)
  );
  FringeFF regs_14 ( // @[RegFile.scala 66:20:@34452.4]
    .clock(regs_14_clock),
    .reset(regs_14_reset),
    .io_in(regs_14_io_in),
    .io_reset(regs_14_io_reset),
    .io_out(regs_14_io_out),
    .io_enable(regs_14_io_enable)
  );
  FringeFF regs_15 ( // @[RegFile.scala 66:20:@34466.4]
    .clock(regs_15_clock),
    .reset(regs_15_reset),
    .io_in(regs_15_io_in),
    .io_reset(regs_15_io_reset),
    .io_out(regs_15_io_out),
    .io_enable(regs_15_io_enable)
  );
  FringeFF regs_16 ( // @[RegFile.scala 66:20:@34480.4]
    .clock(regs_16_clock),
    .reset(regs_16_reset),
    .io_in(regs_16_io_in),
    .io_reset(regs_16_io_reset),
    .io_out(regs_16_io_out),
    .io_enable(regs_16_io_enable)
  );
  FringeFF regs_17 ( // @[RegFile.scala 66:20:@34494.4]
    .clock(regs_17_clock),
    .reset(regs_17_reset),
    .io_in(regs_17_io_in),
    .io_reset(regs_17_io_reset),
    .io_out(regs_17_io_out),
    .io_enable(regs_17_io_enable)
  );
  FringeFF regs_18 ( // @[RegFile.scala 66:20:@34508.4]
    .clock(regs_18_clock),
    .reset(regs_18_reset),
    .io_in(regs_18_io_in),
    .io_reset(regs_18_io_reset),
    .io_out(regs_18_io_out),
    .io_enable(regs_18_io_enable)
  );
  FringeFF regs_19 ( // @[RegFile.scala 66:20:@34522.4]
    .clock(regs_19_clock),
    .reset(regs_19_reset),
    .io_in(regs_19_io_in),
    .io_reset(regs_19_io_reset),
    .io_out(regs_19_io_out),
    .io_enable(regs_19_io_enable)
  );
  FringeFF regs_20 ( // @[RegFile.scala 66:20:@34536.4]
    .clock(regs_20_clock),
    .reset(regs_20_reset),
    .io_in(regs_20_io_in),
    .io_reset(regs_20_io_reset),
    .io_out(regs_20_io_out),
    .io_enable(regs_20_io_enable)
  );
  FringeFF regs_21 ( // @[RegFile.scala 66:20:@34550.4]
    .clock(regs_21_clock),
    .reset(regs_21_reset),
    .io_in(regs_21_io_in),
    .io_reset(regs_21_io_reset),
    .io_out(regs_21_io_out),
    .io_enable(regs_21_io_enable)
  );
  FringeFF regs_22 ( // @[RegFile.scala 66:20:@34564.4]
    .clock(regs_22_clock),
    .reset(regs_22_reset),
    .io_in(regs_22_io_in),
    .io_reset(regs_22_io_reset),
    .io_out(regs_22_io_out),
    .io_enable(regs_22_io_enable)
  );
  FringeFF regs_23 ( // @[RegFile.scala 66:20:@34578.4]
    .clock(regs_23_clock),
    .reset(regs_23_reset),
    .io_in(regs_23_io_in),
    .io_reset(regs_23_io_reset),
    .io_out(regs_23_io_out),
    .io_enable(regs_23_io_enable)
  );
  FringeFF regs_24 ( // @[RegFile.scala 66:20:@34592.4]
    .clock(regs_24_clock),
    .reset(regs_24_reset),
    .io_in(regs_24_io_in),
    .io_reset(regs_24_io_reset),
    .io_out(regs_24_io_out),
    .io_enable(regs_24_io_enable)
  );
  FringeFF regs_25 ( // @[RegFile.scala 66:20:@34606.4]
    .clock(regs_25_clock),
    .reset(regs_25_reset),
    .io_in(regs_25_io_in),
    .io_reset(regs_25_io_reset),
    .io_out(regs_25_io_out),
    .io_enable(regs_25_io_enable)
  );
  FringeFF regs_26 ( // @[RegFile.scala 66:20:@34620.4]
    .clock(regs_26_clock),
    .reset(regs_26_reset),
    .io_in(regs_26_io_in),
    .io_reset(regs_26_io_reset),
    .io_out(regs_26_io_out),
    .io_enable(regs_26_io_enable)
  );
  FringeFF regs_27 ( // @[RegFile.scala 66:20:@34634.4]
    .clock(regs_27_clock),
    .reset(regs_27_reset),
    .io_in(regs_27_io_in),
    .io_reset(regs_27_io_reset),
    .io_out(regs_27_io_out),
    .io_enable(regs_27_io_enable)
  );
  FringeFF regs_28 ( // @[RegFile.scala 66:20:@34648.4]
    .clock(regs_28_clock),
    .reset(regs_28_reset),
    .io_in(regs_28_io_in),
    .io_reset(regs_28_io_reset),
    .io_out(regs_28_io_out),
    .io_enable(regs_28_io_enable)
  );
  FringeFF regs_29 ( // @[RegFile.scala 66:20:@34662.4]
    .clock(regs_29_clock),
    .reset(regs_29_reset),
    .io_in(regs_29_io_in),
    .io_reset(regs_29_io_reset),
    .io_out(regs_29_io_out),
    .io_enable(regs_29_io_enable)
  );
  FringeFF regs_30 ( // @[RegFile.scala 66:20:@34676.4]
    .clock(regs_30_clock),
    .reset(regs_30_reset),
    .io_in(regs_30_io_in),
    .io_reset(regs_30_io_reset),
    .io_out(regs_30_io_out),
    .io_enable(regs_30_io_enable)
  );
  FringeFF regs_31 ( // @[RegFile.scala 66:20:@34690.4]
    .clock(regs_31_clock),
    .reset(regs_31_reset),
    .io_in(regs_31_io_in),
    .io_reset(regs_31_io_reset),
    .io_out(regs_31_io_out),
    .io_enable(regs_31_io_enable)
  );
  FringeFF regs_32 ( // @[RegFile.scala 66:20:@34704.4]
    .clock(regs_32_clock),
    .reset(regs_32_reset),
    .io_in(regs_32_io_in),
    .io_reset(regs_32_io_reset),
    .io_out(regs_32_io_out),
    .io_enable(regs_32_io_enable)
  );
  FringeFF regs_33 ( // @[RegFile.scala 66:20:@34718.4]
    .clock(regs_33_clock),
    .reset(regs_33_reset),
    .io_in(regs_33_io_in),
    .io_reset(regs_33_io_reset),
    .io_out(regs_33_io_out),
    .io_enable(regs_33_io_enable)
  );
  FringeFF regs_34 ( // @[RegFile.scala 66:20:@34732.4]
    .clock(regs_34_clock),
    .reset(regs_34_reset),
    .io_in(regs_34_io_in),
    .io_reset(regs_34_io_reset),
    .io_out(regs_34_io_out),
    .io_enable(regs_34_io_enable)
  );
  FringeFF regs_35 ( // @[RegFile.scala 66:20:@34746.4]
    .clock(regs_35_clock),
    .reset(regs_35_reset),
    .io_in(regs_35_io_in),
    .io_reset(regs_35_io_reset),
    .io_out(regs_35_io_out),
    .io_enable(regs_35_io_enable)
  );
  FringeFF regs_36 ( // @[RegFile.scala 66:20:@34760.4]
    .clock(regs_36_clock),
    .reset(regs_36_reset),
    .io_in(regs_36_io_in),
    .io_reset(regs_36_io_reset),
    .io_out(regs_36_io_out),
    .io_enable(regs_36_io_enable)
  );
  FringeFF regs_37 ( // @[RegFile.scala 66:20:@34774.4]
    .clock(regs_37_clock),
    .reset(regs_37_reset),
    .io_in(regs_37_io_in),
    .io_reset(regs_37_io_reset),
    .io_out(regs_37_io_out),
    .io_enable(regs_37_io_enable)
  );
  FringeFF regs_38 ( // @[RegFile.scala 66:20:@34788.4]
    .clock(regs_38_clock),
    .reset(regs_38_reset),
    .io_in(regs_38_io_in),
    .io_reset(regs_38_io_reset),
    .io_out(regs_38_io_out),
    .io_enable(regs_38_io_enable)
  );
  FringeFF regs_39 ( // @[RegFile.scala 66:20:@34802.4]
    .clock(regs_39_clock),
    .reset(regs_39_reset),
    .io_in(regs_39_io_in),
    .io_reset(regs_39_io_reset),
    .io_out(regs_39_io_out),
    .io_enable(regs_39_io_enable)
  );
  FringeFF regs_40 ( // @[RegFile.scala 66:20:@34816.4]
    .clock(regs_40_clock),
    .reset(regs_40_reset),
    .io_in(regs_40_io_in),
    .io_reset(regs_40_io_reset),
    .io_out(regs_40_io_out),
    .io_enable(regs_40_io_enable)
  );
  FringeFF regs_41 ( // @[RegFile.scala 66:20:@34830.4]
    .clock(regs_41_clock),
    .reset(regs_41_reset),
    .io_in(regs_41_io_in),
    .io_reset(regs_41_io_reset),
    .io_out(regs_41_io_out),
    .io_enable(regs_41_io_enable)
  );
  FringeFF regs_42 ( // @[RegFile.scala 66:20:@34844.4]
    .clock(regs_42_clock),
    .reset(regs_42_reset),
    .io_in(regs_42_io_in),
    .io_reset(regs_42_io_reset),
    .io_out(regs_42_io_out),
    .io_enable(regs_42_io_enable)
  );
  FringeFF regs_43 ( // @[RegFile.scala 66:20:@34858.4]
    .clock(regs_43_clock),
    .reset(regs_43_reset),
    .io_in(regs_43_io_in),
    .io_reset(regs_43_io_reset),
    .io_out(regs_43_io_out),
    .io_enable(regs_43_io_enable)
  );
  FringeFF regs_44 ( // @[RegFile.scala 66:20:@34872.4]
    .clock(regs_44_clock),
    .reset(regs_44_reset),
    .io_in(regs_44_io_in),
    .io_reset(regs_44_io_reset),
    .io_out(regs_44_io_out),
    .io_enable(regs_44_io_enable)
  );
  FringeFF regs_45 ( // @[RegFile.scala 66:20:@34886.4]
    .clock(regs_45_clock),
    .reset(regs_45_reset),
    .io_in(regs_45_io_in),
    .io_reset(regs_45_io_reset),
    .io_out(regs_45_io_out),
    .io_enable(regs_45_io_enable)
  );
  FringeFF regs_46 ( // @[RegFile.scala 66:20:@34900.4]
    .clock(regs_46_clock),
    .reset(regs_46_reset),
    .io_in(regs_46_io_in),
    .io_reset(regs_46_io_reset),
    .io_out(regs_46_io_out),
    .io_enable(regs_46_io_enable)
  );
  FringeFF regs_47 ( // @[RegFile.scala 66:20:@34914.4]
    .clock(regs_47_clock),
    .reset(regs_47_reset),
    .io_in(regs_47_io_in),
    .io_reset(regs_47_io_reset),
    .io_out(regs_47_io_out),
    .io_enable(regs_47_io_enable)
  );
  FringeFF regs_48 ( // @[RegFile.scala 66:20:@34928.4]
    .clock(regs_48_clock),
    .reset(regs_48_reset),
    .io_in(regs_48_io_in),
    .io_reset(regs_48_io_reset),
    .io_out(regs_48_io_out),
    .io_enable(regs_48_io_enable)
  );
  FringeFF regs_49 ( // @[RegFile.scala 66:20:@34942.4]
    .clock(regs_49_clock),
    .reset(regs_49_reset),
    .io_in(regs_49_io_in),
    .io_reset(regs_49_io_reset),
    .io_out(regs_49_io_out),
    .io_enable(regs_49_io_enable)
  );
  FringeFF regs_50 ( // @[RegFile.scala 66:20:@34956.4]
    .clock(regs_50_clock),
    .reset(regs_50_reset),
    .io_in(regs_50_io_in),
    .io_reset(regs_50_io_reset),
    .io_out(regs_50_io_out),
    .io_enable(regs_50_io_enable)
  );
  FringeFF regs_51 ( // @[RegFile.scala 66:20:@34970.4]
    .clock(regs_51_clock),
    .reset(regs_51_reset),
    .io_in(regs_51_io_in),
    .io_reset(regs_51_io_reset),
    .io_out(regs_51_io_out),
    .io_enable(regs_51_io_enable)
  );
  FringeFF regs_52 ( // @[RegFile.scala 66:20:@34984.4]
    .clock(regs_52_clock),
    .reset(regs_52_reset),
    .io_in(regs_52_io_in),
    .io_reset(regs_52_io_reset),
    .io_out(regs_52_io_out),
    .io_enable(regs_52_io_enable)
  );
  FringeFF regs_53 ( // @[RegFile.scala 66:20:@34998.4]
    .clock(regs_53_clock),
    .reset(regs_53_reset),
    .io_in(regs_53_io_in),
    .io_reset(regs_53_io_reset),
    .io_out(regs_53_io_out),
    .io_enable(regs_53_io_enable)
  );
  FringeFF regs_54 ( // @[RegFile.scala 66:20:@35012.4]
    .clock(regs_54_clock),
    .reset(regs_54_reset),
    .io_in(regs_54_io_in),
    .io_reset(regs_54_io_reset),
    .io_out(regs_54_io_out),
    .io_enable(regs_54_io_enable)
  );
  FringeFF regs_55 ( // @[RegFile.scala 66:20:@35026.4]
    .clock(regs_55_clock),
    .reset(regs_55_reset),
    .io_in(regs_55_io_in),
    .io_reset(regs_55_io_reset),
    .io_out(regs_55_io_out),
    .io_enable(regs_55_io_enable)
  );
  FringeFF regs_56 ( // @[RegFile.scala 66:20:@35040.4]
    .clock(regs_56_clock),
    .reset(regs_56_reset),
    .io_in(regs_56_io_in),
    .io_reset(regs_56_io_reset),
    .io_out(regs_56_io_out),
    .io_enable(regs_56_io_enable)
  );
  FringeFF regs_57 ( // @[RegFile.scala 66:20:@35054.4]
    .clock(regs_57_clock),
    .reset(regs_57_reset),
    .io_in(regs_57_io_in),
    .io_reset(regs_57_io_reset),
    .io_out(regs_57_io_out),
    .io_enable(regs_57_io_enable)
  );
  FringeFF regs_58 ( // @[RegFile.scala 66:20:@35068.4]
    .clock(regs_58_clock),
    .reset(regs_58_reset),
    .io_in(regs_58_io_in),
    .io_reset(regs_58_io_reset),
    .io_out(regs_58_io_out),
    .io_enable(regs_58_io_enable)
  );
  FringeFF regs_59 ( // @[RegFile.scala 66:20:@35082.4]
    .clock(regs_59_clock),
    .reset(regs_59_reset),
    .io_in(regs_59_io_in),
    .io_reset(regs_59_io_reset),
    .io_out(regs_59_io_out),
    .io_enable(regs_59_io_enable)
  );
  FringeFF regs_60 ( // @[RegFile.scala 66:20:@35096.4]
    .clock(regs_60_clock),
    .reset(regs_60_reset),
    .io_in(regs_60_io_in),
    .io_reset(regs_60_io_reset),
    .io_out(regs_60_io_out),
    .io_enable(regs_60_io_enable)
  );
  FringeFF regs_61 ( // @[RegFile.scala 66:20:@35110.4]
    .clock(regs_61_clock),
    .reset(regs_61_reset),
    .io_in(regs_61_io_in),
    .io_reset(regs_61_io_reset),
    .io_out(regs_61_io_out),
    .io_enable(regs_61_io_enable)
  );
  FringeFF regs_62 ( // @[RegFile.scala 66:20:@35124.4]
    .clock(regs_62_clock),
    .reset(regs_62_reset),
    .io_in(regs_62_io_in),
    .io_reset(regs_62_io_reset),
    .io_out(regs_62_io_out),
    .io_enable(regs_62_io_enable)
  );
  FringeFF regs_63 ( // @[RegFile.scala 66:20:@35138.4]
    .clock(regs_63_clock),
    .reset(regs_63_reset),
    .io_in(regs_63_io_in),
    .io_reset(regs_63_io_reset),
    .io_out(regs_63_io_out),
    .io_enable(regs_63_io_enable)
  );
  FringeFF regs_64 ( // @[RegFile.scala 66:20:@35152.4]
    .clock(regs_64_clock),
    .reset(regs_64_reset),
    .io_in(regs_64_io_in),
    .io_reset(regs_64_io_reset),
    .io_out(regs_64_io_out),
    .io_enable(regs_64_io_enable)
  );
  FringeFF regs_65 ( // @[RegFile.scala 66:20:@35166.4]
    .clock(regs_65_clock),
    .reset(regs_65_reset),
    .io_in(regs_65_io_in),
    .io_reset(regs_65_io_reset),
    .io_out(regs_65_io_out),
    .io_enable(regs_65_io_enable)
  );
  FringeFF regs_66 ( // @[RegFile.scala 66:20:@35180.4]
    .clock(regs_66_clock),
    .reset(regs_66_reset),
    .io_in(regs_66_io_in),
    .io_reset(regs_66_io_reset),
    .io_out(regs_66_io_out),
    .io_enable(regs_66_io_enable)
  );
  FringeFF regs_67 ( // @[RegFile.scala 66:20:@35194.4]
    .clock(regs_67_clock),
    .reset(regs_67_reset),
    .io_in(regs_67_io_in),
    .io_reset(regs_67_io_reset),
    .io_out(regs_67_io_out),
    .io_enable(regs_67_io_enable)
  );
  FringeFF regs_68 ( // @[RegFile.scala 66:20:@35208.4]
    .clock(regs_68_clock),
    .reset(regs_68_reset),
    .io_in(regs_68_io_in),
    .io_reset(regs_68_io_reset),
    .io_out(regs_68_io_out),
    .io_enable(regs_68_io_enable)
  );
  FringeFF regs_69 ( // @[RegFile.scala 66:20:@35222.4]
    .clock(regs_69_clock),
    .reset(regs_69_reset),
    .io_in(regs_69_io_in),
    .io_reset(regs_69_io_reset),
    .io_out(regs_69_io_out),
    .io_enable(regs_69_io_enable)
  );
  FringeFF regs_70 ( // @[RegFile.scala 66:20:@35236.4]
    .clock(regs_70_clock),
    .reset(regs_70_reset),
    .io_in(regs_70_io_in),
    .io_reset(regs_70_io_reset),
    .io_out(regs_70_io_out),
    .io_enable(regs_70_io_enable)
  );
  FringeFF regs_71 ( // @[RegFile.scala 66:20:@35250.4]
    .clock(regs_71_clock),
    .reset(regs_71_reset),
    .io_in(regs_71_io_in),
    .io_reset(regs_71_io_reset),
    .io_out(regs_71_io_out),
    .io_enable(regs_71_io_enable)
  );
  FringeFF regs_72 ( // @[RegFile.scala 66:20:@35264.4]
    .clock(regs_72_clock),
    .reset(regs_72_reset),
    .io_in(regs_72_io_in),
    .io_reset(regs_72_io_reset),
    .io_out(regs_72_io_out),
    .io_enable(regs_72_io_enable)
  );
  FringeFF regs_73 ( // @[RegFile.scala 66:20:@35278.4]
    .clock(regs_73_clock),
    .reset(regs_73_reset),
    .io_in(regs_73_io_in),
    .io_reset(regs_73_io_reset),
    .io_out(regs_73_io_out),
    .io_enable(regs_73_io_enable)
  );
  FringeFF regs_74 ( // @[RegFile.scala 66:20:@35292.4]
    .clock(regs_74_clock),
    .reset(regs_74_reset),
    .io_in(regs_74_io_in),
    .io_reset(regs_74_io_reset),
    .io_out(regs_74_io_out),
    .io_enable(regs_74_io_enable)
  );
  FringeFF regs_75 ( // @[RegFile.scala 66:20:@35306.4]
    .clock(regs_75_clock),
    .reset(regs_75_reset),
    .io_in(regs_75_io_in),
    .io_reset(regs_75_io_reset),
    .io_out(regs_75_io_out),
    .io_enable(regs_75_io_enable)
  );
  FringeFF regs_76 ( // @[RegFile.scala 66:20:@35320.4]
    .clock(regs_76_clock),
    .reset(regs_76_reset),
    .io_in(regs_76_io_in),
    .io_reset(regs_76_io_reset),
    .io_out(regs_76_io_out),
    .io_enable(regs_76_io_enable)
  );
  FringeFF regs_77 ( // @[RegFile.scala 66:20:@35334.4]
    .clock(regs_77_clock),
    .reset(regs_77_reset),
    .io_in(regs_77_io_in),
    .io_reset(regs_77_io_reset),
    .io_out(regs_77_io_out),
    .io_enable(regs_77_io_enable)
  );
  FringeFF regs_78 ( // @[RegFile.scala 66:20:@35348.4]
    .clock(regs_78_clock),
    .reset(regs_78_reset),
    .io_in(regs_78_io_in),
    .io_reset(regs_78_io_reset),
    .io_out(regs_78_io_out),
    .io_enable(regs_78_io_enable)
  );
  FringeFF regs_79 ( // @[RegFile.scala 66:20:@35362.4]
    .clock(regs_79_clock),
    .reset(regs_79_reset),
    .io_in(regs_79_io_in),
    .io_reset(regs_79_io_reset),
    .io_out(regs_79_io_out),
    .io_enable(regs_79_io_enable)
  );
  FringeFF regs_80 ( // @[RegFile.scala 66:20:@35376.4]
    .clock(regs_80_clock),
    .reset(regs_80_reset),
    .io_in(regs_80_io_in),
    .io_reset(regs_80_io_reset),
    .io_out(regs_80_io_out),
    .io_enable(regs_80_io_enable)
  );
  FringeFF regs_81 ( // @[RegFile.scala 66:20:@35390.4]
    .clock(regs_81_clock),
    .reset(regs_81_reset),
    .io_in(regs_81_io_in),
    .io_reset(regs_81_io_reset),
    .io_out(regs_81_io_out),
    .io_enable(regs_81_io_enable)
  );
  FringeFF regs_82 ( // @[RegFile.scala 66:20:@35404.4]
    .clock(regs_82_clock),
    .reset(regs_82_reset),
    .io_in(regs_82_io_in),
    .io_reset(regs_82_io_reset),
    .io_out(regs_82_io_out),
    .io_enable(regs_82_io_enable)
  );
  FringeFF regs_83 ( // @[RegFile.scala 66:20:@35418.4]
    .clock(regs_83_clock),
    .reset(regs_83_reset),
    .io_in(regs_83_io_in),
    .io_reset(regs_83_io_reset),
    .io_out(regs_83_io_out),
    .io_enable(regs_83_io_enable)
  );
  FringeFF regs_84 ( // @[RegFile.scala 66:20:@35432.4]
    .clock(regs_84_clock),
    .reset(regs_84_reset),
    .io_in(regs_84_io_in),
    .io_reset(regs_84_io_reset),
    .io_out(regs_84_io_out),
    .io_enable(regs_84_io_enable)
  );
  FringeFF regs_85 ( // @[RegFile.scala 66:20:@35446.4]
    .clock(regs_85_clock),
    .reset(regs_85_reset),
    .io_in(regs_85_io_in),
    .io_reset(regs_85_io_reset),
    .io_out(regs_85_io_out),
    .io_enable(regs_85_io_enable)
  );
  FringeFF regs_86 ( // @[RegFile.scala 66:20:@35460.4]
    .clock(regs_86_clock),
    .reset(regs_86_reset),
    .io_in(regs_86_io_in),
    .io_reset(regs_86_io_reset),
    .io_out(regs_86_io_out),
    .io_enable(regs_86_io_enable)
  );
  FringeFF regs_87 ( // @[RegFile.scala 66:20:@35474.4]
    .clock(regs_87_clock),
    .reset(regs_87_reset),
    .io_in(regs_87_io_in),
    .io_reset(regs_87_io_reset),
    .io_out(regs_87_io_out),
    .io_enable(regs_87_io_enable)
  );
  FringeFF regs_88 ( // @[RegFile.scala 66:20:@35488.4]
    .clock(regs_88_clock),
    .reset(regs_88_reset),
    .io_in(regs_88_io_in),
    .io_reset(regs_88_io_reset),
    .io_out(regs_88_io_out),
    .io_enable(regs_88_io_enable)
  );
  FringeFF regs_89 ( // @[RegFile.scala 66:20:@35502.4]
    .clock(regs_89_clock),
    .reset(regs_89_reset),
    .io_in(regs_89_io_in),
    .io_reset(regs_89_io_reset),
    .io_out(regs_89_io_out),
    .io_enable(regs_89_io_enable)
  );
  FringeFF regs_90 ( // @[RegFile.scala 66:20:@35516.4]
    .clock(regs_90_clock),
    .reset(regs_90_reset),
    .io_in(regs_90_io_in),
    .io_reset(regs_90_io_reset),
    .io_out(regs_90_io_out),
    .io_enable(regs_90_io_enable)
  );
  FringeFF regs_91 ( // @[RegFile.scala 66:20:@35530.4]
    .clock(regs_91_clock),
    .reset(regs_91_reset),
    .io_in(regs_91_io_in),
    .io_reset(regs_91_io_reset),
    .io_out(regs_91_io_out),
    .io_enable(regs_91_io_enable)
  );
  FringeFF regs_92 ( // @[RegFile.scala 66:20:@35544.4]
    .clock(regs_92_clock),
    .reset(regs_92_reset),
    .io_in(regs_92_io_in),
    .io_reset(regs_92_io_reset),
    .io_out(regs_92_io_out),
    .io_enable(regs_92_io_enable)
  );
  FringeFF regs_93 ( // @[RegFile.scala 66:20:@35558.4]
    .clock(regs_93_clock),
    .reset(regs_93_reset),
    .io_in(regs_93_io_in),
    .io_reset(regs_93_io_reset),
    .io_out(regs_93_io_out),
    .io_enable(regs_93_io_enable)
  );
  FringeFF regs_94 ( // @[RegFile.scala 66:20:@35572.4]
    .clock(regs_94_clock),
    .reset(regs_94_reset),
    .io_in(regs_94_io_in),
    .io_reset(regs_94_io_reset),
    .io_out(regs_94_io_out),
    .io_enable(regs_94_io_enable)
  );
  FringeFF regs_95 ( // @[RegFile.scala 66:20:@35586.4]
    .clock(regs_95_clock),
    .reset(regs_95_reset),
    .io_in(regs_95_io_in),
    .io_reset(regs_95_io_reset),
    .io_out(regs_95_io_out),
    .io_enable(regs_95_io_enable)
  );
  FringeFF regs_96 ( // @[RegFile.scala 66:20:@35600.4]
    .clock(regs_96_clock),
    .reset(regs_96_reset),
    .io_in(regs_96_io_in),
    .io_reset(regs_96_io_reset),
    .io_out(regs_96_io_out),
    .io_enable(regs_96_io_enable)
  );
  FringeFF regs_97 ( // @[RegFile.scala 66:20:@35614.4]
    .clock(regs_97_clock),
    .reset(regs_97_reset),
    .io_in(regs_97_io_in),
    .io_reset(regs_97_io_reset),
    .io_out(regs_97_io_out),
    .io_enable(regs_97_io_enable)
  );
  FringeFF regs_98 ( // @[RegFile.scala 66:20:@35628.4]
    .clock(regs_98_clock),
    .reset(regs_98_reset),
    .io_in(regs_98_io_in),
    .io_reset(regs_98_io_reset),
    .io_out(regs_98_io_out),
    .io_enable(regs_98_io_enable)
  );
  FringeFF regs_99 ( // @[RegFile.scala 66:20:@35642.4]
    .clock(regs_99_clock),
    .reset(regs_99_reset),
    .io_in(regs_99_io_in),
    .io_reset(regs_99_io_reset),
    .io_out(regs_99_io_out),
    .io_enable(regs_99_io_enable)
  );
  FringeFF regs_100 ( // @[RegFile.scala 66:20:@35656.4]
    .clock(regs_100_clock),
    .reset(regs_100_reset),
    .io_in(regs_100_io_in),
    .io_reset(regs_100_io_reset),
    .io_out(regs_100_io_out),
    .io_enable(regs_100_io_enable)
  );
  FringeFF regs_101 ( // @[RegFile.scala 66:20:@35670.4]
    .clock(regs_101_clock),
    .reset(regs_101_reset),
    .io_in(regs_101_io_in),
    .io_reset(regs_101_io_reset),
    .io_out(regs_101_io_out),
    .io_enable(regs_101_io_enable)
  );
  FringeFF regs_102 ( // @[RegFile.scala 66:20:@35684.4]
    .clock(regs_102_clock),
    .reset(regs_102_reset),
    .io_in(regs_102_io_in),
    .io_reset(regs_102_io_reset),
    .io_out(regs_102_io_out),
    .io_enable(regs_102_io_enable)
  );
  FringeFF regs_103 ( // @[RegFile.scala 66:20:@35698.4]
    .clock(regs_103_clock),
    .reset(regs_103_reset),
    .io_in(regs_103_io_in),
    .io_reset(regs_103_io_reset),
    .io_out(regs_103_io_out),
    .io_enable(regs_103_io_enable)
  );
  FringeFF regs_104 ( // @[RegFile.scala 66:20:@35712.4]
    .clock(regs_104_clock),
    .reset(regs_104_reset),
    .io_in(regs_104_io_in),
    .io_reset(regs_104_io_reset),
    .io_out(regs_104_io_out),
    .io_enable(regs_104_io_enable)
  );
  FringeFF regs_105 ( // @[RegFile.scala 66:20:@35726.4]
    .clock(regs_105_clock),
    .reset(regs_105_reset),
    .io_in(regs_105_io_in),
    .io_reset(regs_105_io_reset),
    .io_out(regs_105_io_out),
    .io_enable(regs_105_io_enable)
  );
  FringeFF regs_106 ( // @[RegFile.scala 66:20:@35740.4]
    .clock(regs_106_clock),
    .reset(regs_106_reset),
    .io_in(regs_106_io_in),
    .io_reset(regs_106_io_reset),
    .io_out(regs_106_io_out),
    .io_enable(regs_106_io_enable)
  );
  FringeFF regs_107 ( // @[RegFile.scala 66:20:@35754.4]
    .clock(regs_107_clock),
    .reset(regs_107_reset),
    .io_in(regs_107_io_in),
    .io_reset(regs_107_io_reset),
    .io_out(regs_107_io_out),
    .io_enable(regs_107_io_enable)
  );
  FringeFF regs_108 ( // @[RegFile.scala 66:20:@35768.4]
    .clock(regs_108_clock),
    .reset(regs_108_reset),
    .io_in(regs_108_io_in),
    .io_reset(regs_108_io_reset),
    .io_out(regs_108_io_out),
    .io_enable(regs_108_io_enable)
  );
  FringeFF regs_109 ( // @[RegFile.scala 66:20:@35782.4]
    .clock(regs_109_clock),
    .reset(regs_109_reset),
    .io_in(regs_109_io_in),
    .io_reset(regs_109_io_reset),
    .io_out(regs_109_io_out),
    .io_enable(regs_109_io_enable)
  );
  FringeFF regs_110 ( // @[RegFile.scala 66:20:@35796.4]
    .clock(regs_110_clock),
    .reset(regs_110_reset),
    .io_in(regs_110_io_in),
    .io_reset(regs_110_io_reset),
    .io_out(regs_110_io_out),
    .io_enable(regs_110_io_enable)
  );
  FringeFF regs_111 ( // @[RegFile.scala 66:20:@35810.4]
    .clock(regs_111_clock),
    .reset(regs_111_reset),
    .io_in(regs_111_io_in),
    .io_reset(regs_111_io_reset),
    .io_out(regs_111_io_out),
    .io_enable(regs_111_io_enable)
  );
  FringeFF regs_112 ( // @[RegFile.scala 66:20:@35824.4]
    .clock(regs_112_clock),
    .reset(regs_112_reset),
    .io_in(regs_112_io_in),
    .io_reset(regs_112_io_reset),
    .io_out(regs_112_io_out),
    .io_enable(regs_112_io_enable)
  );
  FringeFF regs_113 ( // @[RegFile.scala 66:20:@35838.4]
    .clock(regs_113_clock),
    .reset(regs_113_reset),
    .io_in(regs_113_io_in),
    .io_reset(regs_113_io_reset),
    .io_out(regs_113_io_out),
    .io_enable(regs_113_io_enable)
  );
  FringeFF regs_114 ( // @[RegFile.scala 66:20:@35852.4]
    .clock(regs_114_clock),
    .reset(regs_114_reset),
    .io_in(regs_114_io_in),
    .io_reset(regs_114_io_reset),
    .io_out(regs_114_io_out),
    .io_enable(regs_114_io_enable)
  );
  FringeFF regs_115 ( // @[RegFile.scala 66:20:@35866.4]
    .clock(regs_115_clock),
    .reset(regs_115_reset),
    .io_in(regs_115_io_in),
    .io_reset(regs_115_io_reset),
    .io_out(regs_115_io_out),
    .io_enable(regs_115_io_enable)
  );
  FringeFF regs_116 ( // @[RegFile.scala 66:20:@35880.4]
    .clock(regs_116_clock),
    .reset(regs_116_reset),
    .io_in(regs_116_io_in),
    .io_reset(regs_116_io_reset),
    .io_out(regs_116_io_out),
    .io_enable(regs_116_io_enable)
  );
  FringeFF regs_117 ( // @[RegFile.scala 66:20:@35894.4]
    .clock(regs_117_clock),
    .reset(regs_117_reset),
    .io_in(regs_117_io_in),
    .io_reset(regs_117_io_reset),
    .io_out(regs_117_io_out),
    .io_enable(regs_117_io_enable)
  );
  FringeFF regs_118 ( // @[RegFile.scala 66:20:@35908.4]
    .clock(regs_118_clock),
    .reset(regs_118_reset),
    .io_in(regs_118_io_in),
    .io_reset(regs_118_io_reset),
    .io_out(regs_118_io_out),
    .io_enable(regs_118_io_enable)
  );
  FringeFF regs_119 ( // @[RegFile.scala 66:20:@35922.4]
    .clock(regs_119_clock),
    .reset(regs_119_reset),
    .io_in(regs_119_io_in),
    .io_reset(regs_119_io_reset),
    .io_out(regs_119_io_out),
    .io_enable(regs_119_io_enable)
  );
  FringeFF regs_120 ( // @[RegFile.scala 66:20:@35936.4]
    .clock(regs_120_clock),
    .reset(regs_120_reset),
    .io_in(regs_120_io_in),
    .io_reset(regs_120_io_reset),
    .io_out(regs_120_io_out),
    .io_enable(regs_120_io_enable)
  );
  FringeFF regs_121 ( // @[RegFile.scala 66:20:@35950.4]
    .clock(regs_121_clock),
    .reset(regs_121_reset),
    .io_in(regs_121_io_in),
    .io_reset(regs_121_io_reset),
    .io_out(regs_121_io_out),
    .io_enable(regs_121_io_enable)
  );
  FringeFF regs_122 ( // @[RegFile.scala 66:20:@35964.4]
    .clock(regs_122_clock),
    .reset(regs_122_reset),
    .io_in(regs_122_io_in),
    .io_reset(regs_122_io_reset),
    .io_out(regs_122_io_out),
    .io_enable(regs_122_io_enable)
  );
  FringeFF regs_123 ( // @[RegFile.scala 66:20:@35978.4]
    .clock(regs_123_clock),
    .reset(regs_123_reset),
    .io_in(regs_123_io_in),
    .io_reset(regs_123_io_reset),
    .io_out(regs_123_io_out),
    .io_enable(regs_123_io_enable)
  );
  FringeFF regs_124 ( // @[RegFile.scala 66:20:@35992.4]
    .clock(regs_124_clock),
    .reset(regs_124_reset),
    .io_in(regs_124_io_in),
    .io_reset(regs_124_io_reset),
    .io_out(regs_124_io_out),
    .io_enable(regs_124_io_enable)
  );
  FringeFF regs_125 ( // @[RegFile.scala 66:20:@36006.4]
    .clock(regs_125_clock),
    .reset(regs_125_reset),
    .io_in(regs_125_io_in),
    .io_reset(regs_125_io_reset),
    .io_out(regs_125_io_out),
    .io_enable(regs_125_io_enable)
  );
  FringeFF regs_126 ( // @[RegFile.scala 66:20:@36020.4]
    .clock(regs_126_clock),
    .reset(regs_126_reset),
    .io_in(regs_126_io_in),
    .io_reset(regs_126_io_reset),
    .io_out(regs_126_io_out),
    .io_enable(regs_126_io_enable)
  );
  FringeFF regs_127 ( // @[RegFile.scala 66:20:@36034.4]
    .clock(regs_127_clock),
    .reset(regs_127_reset),
    .io_in(regs_127_io_in),
    .io_reset(regs_127_io_reset),
    .io_out(regs_127_io_out),
    .io_enable(regs_127_io_enable)
  );
  FringeFF regs_128 ( // @[RegFile.scala 66:20:@36048.4]
    .clock(regs_128_clock),
    .reset(regs_128_reset),
    .io_in(regs_128_io_in),
    .io_reset(regs_128_io_reset),
    .io_out(regs_128_io_out),
    .io_enable(regs_128_io_enable)
  );
  FringeFF regs_129 ( // @[RegFile.scala 66:20:@36062.4]
    .clock(regs_129_clock),
    .reset(regs_129_reset),
    .io_in(regs_129_io_in),
    .io_reset(regs_129_io_reset),
    .io_out(regs_129_io_out),
    .io_enable(regs_129_io_enable)
  );
  FringeFF regs_130 ( // @[RegFile.scala 66:20:@36076.4]
    .clock(regs_130_clock),
    .reset(regs_130_reset),
    .io_in(regs_130_io_in),
    .io_reset(regs_130_io_reset),
    .io_out(regs_130_io_out),
    .io_enable(regs_130_io_enable)
  );
  FringeFF regs_131 ( // @[RegFile.scala 66:20:@36090.4]
    .clock(regs_131_clock),
    .reset(regs_131_reset),
    .io_in(regs_131_io_in),
    .io_reset(regs_131_io_reset),
    .io_out(regs_131_io_out),
    .io_enable(regs_131_io_enable)
  );
  FringeFF regs_132 ( // @[RegFile.scala 66:20:@36104.4]
    .clock(regs_132_clock),
    .reset(regs_132_reset),
    .io_in(regs_132_io_in),
    .io_reset(regs_132_io_reset),
    .io_out(regs_132_io_out),
    .io_enable(regs_132_io_enable)
  );
  FringeFF regs_133 ( // @[RegFile.scala 66:20:@36118.4]
    .clock(regs_133_clock),
    .reset(regs_133_reset),
    .io_in(regs_133_io_in),
    .io_reset(regs_133_io_reset),
    .io_out(regs_133_io_out),
    .io_enable(regs_133_io_enable)
  );
  FringeFF regs_134 ( // @[RegFile.scala 66:20:@36132.4]
    .clock(regs_134_clock),
    .reset(regs_134_reset),
    .io_in(regs_134_io_in),
    .io_reset(regs_134_io_reset),
    .io_out(regs_134_io_out),
    .io_enable(regs_134_io_enable)
  );
  FringeFF regs_135 ( // @[RegFile.scala 66:20:@36146.4]
    .clock(regs_135_clock),
    .reset(regs_135_reset),
    .io_in(regs_135_io_in),
    .io_reset(regs_135_io_reset),
    .io_out(regs_135_io_out),
    .io_enable(regs_135_io_enable)
  );
  FringeFF regs_136 ( // @[RegFile.scala 66:20:@36160.4]
    .clock(regs_136_clock),
    .reset(regs_136_reset),
    .io_in(regs_136_io_in),
    .io_reset(regs_136_io_reset),
    .io_out(regs_136_io_out),
    .io_enable(regs_136_io_enable)
  );
  FringeFF regs_137 ( // @[RegFile.scala 66:20:@36174.4]
    .clock(regs_137_clock),
    .reset(regs_137_reset),
    .io_in(regs_137_io_in),
    .io_reset(regs_137_io_reset),
    .io_out(regs_137_io_out),
    .io_enable(regs_137_io_enable)
  );
  FringeFF regs_138 ( // @[RegFile.scala 66:20:@36188.4]
    .clock(regs_138_clock),
    .reset(regs_138_reset),
    .io_in(regs_138_io_in),
    .io_reset(regs_138_io_reset),
    .io_out(regs_138_io_out),
    .io_enable(regs_138_io_enable)
  );
  FringeFF regs_139 ( // @[RegFile.scala 66:20:@36202.4]
    .clock(regs_139_clock),
    .reset(regs_139_reset),
    .io_in(regs_139_io_in),
    .io_reset(regs_139_io_reset),
    .io_out(regs_139_io_out),
    .io_enable(regs_139_io_enable)
  );
  FringeFF regs_140 ( // @[RegFile.scala 66:20:@36216.4]
    .clock(regs_140_clock),
    .reset(regs_140_reset),
    .io_in(regs_140_io_in),
    .io_reset(regs_140_io_reset),
    .io_out(regs_140_io_out),
    .io_enable(regs_140_io_enable)
  );
  FringeFF regs_141 ( // @[RegFile.scala 66:20:@36230.4]
    .clock(regs_141_clock),
    .reset(regs_141_reset),
    .io_in(regs_141_io_in),
    .io_reset(regs_141_io_reset),
    .io_out(regs_141_io_out),
    .io_enable(regs_141_io_enable)
  );
  FringeFF regs_142 ( // @[RegFile.scala 66:20:@36244.4]
    .clock(regs_142_clock),
    .reset(regs_142_reset),
    .io_in(regs_142_io_in),
    .io_reset(regs_142_io_reset),
    .io_out(regs_142_io_out),
    .io_enable(regs_142_io_enable)
  );
  FringeFF regs_143 ( // @[RegFile.scala 66:20:@36258.4]
    .clock(regs_143_clock),
    .reset(regs_143_reset),
    .io_in(regs_143_io_in),
    .io_reset(regs_143_io_reset),
    .io_out(regs_143_io_out),
    .io_enable(regs_143_io_enable)
  );
  FringeFF regs_144 ( // @[RegFile.scala 66:20:@36272.4]
    .clock(regs_144_clock),
    .reset(regs_144_reset),
    .io_in(regs_144_io_in),
    .io_reset(regs_144_io_reset),
    .io_out(regs_144_io_out),
    .io_enable(regs_144_io_enable)
  );
  FringeFF regs_145 ( // @[RegFile.scala 66:20:@36286.4]
    .clock(regs_145_clock),
    .reset(regs_145_reset),
    .io_in(regs_145_io_in),
    .io_reset(regs_145_io_reset),
    .io_out(regs_145_io_out),
    .io_enable(regs_145_io_enable)
  );
  FringeFF regs_146 ( // @[RegFile.scala 66:20:@36300.4]
    .clock(regs_146_clock),
    .reset(regs_146_reset),
    .io_in(regs_146_io_in),
    .io_reset(regs_146_io_reset),
    .io_out(regs_146_io_out),
    .io_enable(regs_146_io_enable)
  );
  FringeFF regs_147 ( // @[RegFile.scala 66:20:@36314.4]
    .clock(regs_147_clock),
    .reset(regs_147_reset),
    .io_in(regs_147_io_in),
    .io_reset(regs_147_io_reset),
    .io_out(regs_147_io_out),
    .io_enable(regs_147_io_enable)
  );
  FringeFF regs_148 ( // @[RegFile.scala 66:20:@36328.4]
    .clock(regs_148_clock),
    .reset(regs_148_reset),
    .io_in(regs_148_io_in),
    .io_reset(regs_148_io_reset),
    .io_out(regs_148_io_out),
    .io_enable(regs_148_io_enable)
  );
  FringeFF regs_149 ( // @[RegFile.scala 66:20:@36342.4]
    .clock(regs_149_clock),
    .reset(regs_149_reset),
    .io_in(regs_149_io_in),
    .io_reset(regs_149_io_reset),
    .io_out(regs_149_io_out),
    .io_enable(regs_149_io_enable)
  );
  FringeFF regs_150 ( // @[RegFile.scala 66:20:@36356.4]
    .clock(regs_150_clock),
    .reset(regs_150_reset),
    .io_in(regs_150_io_in),
    .io_reset(regs_150_io_reset),
    .io_out(regs_150_io_out),
    .io_enable(regs_150_io_enable)
  );
  FringeFF regs_151 ( // @[RegFile.scala 66:20:@36370.4]
    .clock(regs_151_clock),
    .reset(regs_151_reset),
    .io_in(regs_151_io_in),
    .io_reset(regs_151_io_reset),
    .io_out(regs_151_io_out),
    .io_enable(regs_151_io_enable)
  );
  FringeFF regs_152 ( // @[RegFile.scala 66:20:@36384.4]
    .clock(regs_152_clock),
    .reset(regs_152_reset),
    .io_in(regs_152_io_in),
    .io_reset(regs_152_io_reset),
    .io_out(regs_152_io_out),
    .io_enable(regs_152_io_enable)
  );
  FringeFF regs_153 ( // @[RegFile.scala 66:20:@36398.4]
    .clock(regs_153_clock),
    .reset(regs_153_reset),
    .io_in(regs_153_io_in),
    .io_reset(regs_153_io_reset),
    .io_out(regs_153_io_out),
    .io_enable(regs_153_io_enable)
  );
  FringeFF regs_154 ( // @[RegFile.scala 66:20:@36412.4]
    .clock(regs_154_clock),
    .reset(regs_154_reset),
    .io_in(regs_154_io_in),
    .io_reset(regs_154_io_reset),
    .io_out(regs_154_io_out),
    .io_enable(regs_154_io_enable)
  );
  FringeFF regs_155 ( // @[RegFile.scala 66:20:@36426.4]
    .clock(regs_155_clock),
    .reset(regs_155_reset),
    .io_in(regs_155_io_in),
    .io_reset(regs_155_io_reset),
    .io_out(regs_155_io_out),
    .io_enable(regs_155_io_enable)
  );
  FringeFF regs_156 ( // @[RegFile.scala 66:20:@36440.4]
    .clock(regs_156_clock),
    .reset(regs_156_reset),
    .io_in(regs_156_io_in),
    .io_reset(regs_156_io_reset),
    .io_out(regs_156_io_out),
    .io_enable(regs_156_io_enable)
  );
  FringeFF regs_157 ( // @[RegFile.scala 66:20:@36454.4]
    .clock(regs_157_clock),
    .reset(regs_157_reset),
    .io_in(regs_157_io_in),
    .io_reset(regs_157_io_reset),
    .io_out(regs_157_io_out),
    .io_enable(regs_157_io_enable)
  );
  FringeFF regs_158 ( // @[RegFile.scala 66:20:@36468.4]
    .clock(regs_158_clock),
    .reset(regs_158_reset),
    .io_in(regs_158_io_in),
    .io_reset(regs_158_io_reset),
    .io_out(regs_158_io_out),
    .io_enable(regs_158_io_enable)
  );
  FringeFF regs_159 ( // @[RegFile.scala 66:20:@36482.4]
    .clock(regs_159_clock),
    .reset(regs_159_reset),
    .io_in(regs_159_io_in),
    .io_reset(regs_159_io_reset),
    .io_out(regs_159_io_out),
    .io_enable(regs_159_io_enable)
  );
  FringeFF regs_160 ( // @[RegFile.scala 66:20:@36496.4]
    .clock(regs_160_clock),
    .reset(regs_160_reset),
    .io_in(regs_160_io_in),
    .io_reset(regs_160_io_reset),
    .io_out(regs_160_io_out),
    .io_enable(regs_160_io_enable)
  );
  FringeFF regs_161 ( // @[RegFile.scala 66:20:@36510.4]
    .clock(regs_161_clock),
    .reset(regs_161_reset),
    .io_in(regs_161_io_in),
    .io_reset(regs_161_io_reset),
    .io_out(regs_161_io_out),
    .io_enable(regs_161_io_enable)
  );
  FringeFF regs_162 ( // @[RegFile.scala 66:20:@36524.4]
    .clock(regs_162_clock),
    .reset(regs_162_reset),
    .io_in(regs_162_io_in),
    .io_reset(regs_162_io_reset),
    .io_out(regs_162_io_out),
    .io_enable(regs_162_io_enable)
  );
  FringeFF regs_163 ( // @[RegFile.scala 66:20:@36538.4]
    .clock(regs_163_clock),
    .reset(regs_163_reset),
    .io_in(regs_163_io_in),
    .io_reset(regs_163_io_reset),
    .io_out(regs_163_io_out),
    .io_enable(regs_163_io_enable)
  );
  FringeFF regs_164 ( // @[RegFile.scala 66:20:@36552.4]
    .clock(regs_164_clock),
    .reset(regs_164_reset),
    .io_in(regs_164_io_in),
    .io_reset(regs_164_io_reset),
    .io_out(regs_164_io_out),
    .io_enable(regs_164_io_enable)
  );
  FringeFF regs_165 ( // @[RegFile.scala 66:20:@36566.4]
    .clock(regs_165_clock),
    .reset(regs_165_reset),
    .io_in(regs_165_io_in),
    .io_reset(regs_165_io_reset),
    .io_out(regs_165_io_out),
    .io_enable(regs_165_io_enable)
  );
  FringeFF regs_166 ( // @[RegFile.scala 66:20:@36580.4]
    .clock(regs_166_clock),
    .reset(regs_166_reset),
    .io_in(regs_166_io_in),
    .io_reset(regs_166_io_reset),
    .io_out(regs_166_io_out),
    .io_enable(regs_166_io_enable)
  );
  FringeFF regs_167 ( // @[RegFile.scala 66:20:@36594.4]
    .clock(regs_167_clock),
    .reset(regs_167_reset),
    .io_in(regs_167_io_in),
    .io_reset(regs_167_io_reset),
    .io_out(regs_167_io_out),
    .io_enable(regs_167_io_enable)
  );
  FringeFF regs_168 ( // @[RegFile.scala 66:20:@36608.4]
    .clock(regs_168_clock),
    .reset(regs_168_reset),
    .io_in(regs_168_io_in),
    .io_reset(regs_168_io_reset),
    .io_out(regs_168_io_out),
    .io_enable(regs_168_io_enable)
  );
  FringeFF regs_169 ( // @[RegFile.scala 66:20:@36622.4]
    .clock(regs_169_clock),
    .reset(regs_169_reset),
    .io_in(regs_169_io_in),
    .io_reset(regs_169_io_reset),
    .io_out(regs_169_io_out),
    .io_enable(regs_169_io_enable)
  );
  FringeFF regs_170 ( // @[RegFile.scala 66:20:@36636.4]
    .clock(regs_170_clock),
    .reset(regs_170_reset),
    .io_in(regs_170_io_in),
    .io_reset(regs_170_io_reset),
    .io_out(regs_170_io_out),
    .io_enable(regs_170_io_enable)
  );
  FringeFF regs_171 ( // @[RegFile.scala 66:20:@36650.4]
    .clock(regs_171_clock),
    .reset(regs_171_reset),
    .io_in(regs_171_io_in),
    .io_reset(regs_171_io_reset),
    .io_out(regs_171_io_out),
    .io_enable(regs_171_io_enable)
  );
  FringeFF regs_172 ( // @[RegFile.scala 66:20:@36664.4]
    .clock(regs_172_clock),
    .reset(regs_172_reset),
    .io_in(regs_172_io_in),
    .io_reset(regs_172_io_reset),
    .io_out(regs_172_io_out),
    .io_enable(regs_172_io_enable)
  );
  FringeFF regs_173 ( // @[RegFile.scala 66:20:@36678.4]
    .clock(regs_173_clock),
    .reset(regs_173_reset),
    .io_in(regs_173_io_in),
    .io_reset(regs_173_io_reset),
    .io_out(regs_173_io_out),
    .io_enable(regs_173_io_enable)
  );
  FringeFF regs_174 ( // @[RegFile.scala 66:20:@36692.4]
    .clock(regs_174_clock),
    .reset(regs_174_reset),
    .io_in(regs_174_io_in),
    .io_reset(regs_174_io_reset),
    .io_out(regs_174_io_out),
    .io_enable(regs_174_io_enable)
  );
  FringeFF regs_175 ( // @[RegFile.scala 66:20:@36706.4]
    .clock(regs_175_clock),
    .reset(regs_175_reset),
    .io_in(regs_175_io_in),
    .io_reset(regs_175_io_reset),
    .io_out(regs_175_io_out),
    .io_enable(regs_175_io_enable)
  );
  FringeFF regs_176 ( // @[RegFile.scala 66:20:@36720.4]
    .clock(regs_176_clock),
    .reset(regs_176_reset),
    .io_in(regs_176_io_in),
    .io_reset(regs_176_io_reset),
    .io_out(regs_176_io_out),
    .io_enable(regs_176_io_enable)
  );
  FringeFF regs_177 ( // @[RegFile.scala 66:20:@36734.4]
    .clock(regs_177_clock),
    .reset(regs_177_reset),
    .io_in(regs_177_io_in),
    .io_reset(regs_177_io_reset),
    .io_out(regs_177_io_out),
    .io_enable(regs_177_io_enable)
  );
  FringeFF regs_178 ( // @[RegFile.scala 66:20:@36748.4]
    .clock(regs_178_clock),
    .reset(regs_178_reset),
    .io_in(regs_178_io_in),
    .io_reset(regs_178_io_reset),
    .io_out(regs_178_io_out),
    .io_enable(regs_178_io_enable)
  );
  FringeFF regs_179 ( // @[RegFile.scala 66:20:@36762.4]
    .clock(regs_179_clock),
    .reset(regs_179_reset),
    .io_in(regs_179_io_in),
    .io_reset(regs_179_io_reset),
    .io_out(regs_179_io_out),
    .io_enable(regs_179_io_enable)
  );
  FringeFF regs_180 ( // @[RegFile.scala 66:20:@36776.4]
    .clock(regs_180_clock),
    .reset(regs_180_reset),
    .io_in(regs_180_io_in),
    .io_reset(regs_180_io_reset),
    .io_out(regs_180_io_out),
    .io_enable(regs_180_io_enable)
  );
  FringeFF regs_181 ( // @[RegFile.scala 66:20:@36790.4]
    .clock(regs_181_clock),
    .reset(regs_181_reset),
    .io_in(regs_181_io_in),
    .io_reset(regs_181_io_reset),
    .io_out(regs_181_io_out),
    .io_enable(regs_181_io_enable)
  );
  FringeFF regs_182 ( // @[RegFile.scala 66:20:@36804.4]
    .clock(regs_182_clock),
    .reset(regs_182_reset),
    .io_in(regs_182_io_in),
    .io_reset(regs_182_io_reset),
    .io_out(regs_182_io_out),
    .io_enable(regs_182_io_enable)
  );
  FringeFF regs_183 ( // @[RegFile.scala 66:20:@36818.4]
    .clock(regs_183_clock),
    .reset(regs_183_reset),
    .io_in(regs_183_io_in),
    .io_reset(regs_183_io_reset),
    .io_out(regs_183_io_out),
    .io_enable(regs_183_io_enable)
  );
  FringeFF regs_184 ( // @[RegFile.scala 66:20:@36832.4]
    .clock(regs_184_clock),
    .reset(regs_184_reset),
    .io_in(regs_184_io_in),
    .io_reset(regs_184_io_reset),
    .io_out(regs_184_io_out),
    .io_enable(regs_184_io_enable)
  );
  FringeFF regs_185 ( // @[RegFile.scala 66:20:@36846.4]
    .clock(regs_185_clock),
    .reset(regs_185_reset),
    .io_in(regs_185_io_in),
    .io_reset(regs_185_io_reset),
    .io_out(regs_185_io_out),
    .io_enable(regs_185_io_enable)
  );
  FringeFF regs_186 ( // @[RegFile.scala 66:20:@36860.4]
    .clock(regs_186_clock),
    .reset(regs_186_reset),
    .io_in(regs_186_io_in),
    .io_reset(regs_186_io_reset),
    .io_out(regs_186_io_out),
    .io_enable(regs_186_io_enable)
  );
  FringeFF regs_187 ( // @[RegFile.scala 66:20:@36874.4]
    .clock(regs_187_clock),
    .reset(regs_187_reset),
    .io_in(regs_187_io_in),
    .io_reset(regs_187_io_reset),
    .io_out(regs_187_io_out),
    .io_enable(regs_187_io_enable)
  );
  FringeFF regs_188 ( // @[RegFile.scala 66:20:@36888.4]
    .clock(regs_188_clock),
    .reset(regs_188_reset),
    .io_in(regs_188_io_in),
    .io_reset(regs_188_io_reset),
    .io_out(regs_188_io_out),
    .io_enable(regs_188_io_enable)
  );
  FringeFF regs_189 ( // @[RegFile.scala 66:20:@36902.4]
    .clock(regs_189_clock),
    .reset(regs_189_reset),
    .io_in(regs_189_io_in),
    .io_reset(regs_189_io_reset),
    .io_out(regs_189_io_out),
    .io_enable(regs_189_io_enable)
  );
  FringeFF regs_190 ( // @[RegFile.scala 66:20:@36916.4]
    .clock(regs_190_clock),
    .reset(regs_190_reset),
    .io_in(regs_190_io_in),
    .io_reset(regs_190_io_reset),
    .io_out(regs_190_io_out),
    .io_enable(regs_190_io_enable)
  );
  FringeFF regs_191 ( // @[RegFile.scala 66:20:@36930.4]
    .clock(regs_191_clock),
    .reset(regs_191_reset),
    .io_in(regs_191_io_in),
    .io_reset(regs_191_io_reset),
    .io_out(regs_191_io_out),
    .io_enable(regs_191_io_enable)
  );
  FringeFF regs_192 ( // @[RegFile.scala 66:20:@36944.4]
    .clock(regs_192_clock),
    .reset(regs_192_reset),
    .io_in(regs_192_io_in),
    .io_reset(regs_192_io_reset),
    .io_out(regs_192_io_out),
    .io_enable(regs_192_io_enable)
  );
  FringeFF regs_193 ( // @[RegFile.scala 66:20:@36958.4]
    .clock(regs_193_clock),
    .reset(regs_193_reset),
    .io_in(regs_193_io_in),
    .io_reset(regs_193_io_reset),
    .io_out(regs_193_io_out),
    .io_enable(regs_193_io_enable)
  );
  FringeFF regs_194 ( // @[RegFile.scala 66:20:@36972.4]
    .clock(regs_194_clock),
    .reset(regs_194_reset),
    .io_in(regs_194_io_in),
    .io_reset(regs_194_io_reset),
    .io_out(regs_194_io_out),
    .io_enable(regs_194_io_enable)
  );
  FringeFF regs_195 ( // @[RegFile.scala 66:20:@36986.4]
    .clock(regs_195_clock),
    .reset(regs_195_reset),
    .io_in(regs_195_io_in),
    .io_reset(regs_195_io_reset),
    .io_out(regs_195_io_out),
    .io_enable(regs_195_io_enable)
  );
  FringeFF regs_196 ( // @[RegFile.scala 66:20:@37000.4]
    .clock(regs_196_clock),
    .reset(regs_196_reset),
    .io_in(regs_196_io_in),
    .io_reset(regs_196_io_reset),
    .io_out(regs_196_io_out),
    .io_enable(regs_196_io_enable)
  );
  FringeFF regs_197 ( // @[RegFile.scala 66:20:@37014.4]
    .clock(regs_197_clock),
    .reset(regs_197_reset),
    .io_in(regs_197_io_in),
    .io_reset(regs_197_io_reset),
    .io_out(regs_197_io_out),
    .io_enable(regs_197_io_enable)
  );
  FringeFF regs_198 ( // @[RegFile.scala 66:20:@37028.4]
    .clock(regs_198_clock),
    .reset(regs_198_reset),
    .io_in(regs_198_io_in),
    .io_reset(regs_198_io_reset),
    .io_out(regs_198_io_out),
    .io_enable(regs_198_io_enable)
  );
  FringeFF regs_199 ( // @[RegFile.scala 66:20:@37042.4]
    .clock(regs_199_clock),
    .reset(regs_199_reset),
    .io_in(regs_199_io_in),
    .io_reset(regs_199_io_reset),
    .io_out(regs_199_io_out),
    .io_enable(regs_199_io_enable)
  );
  FringeFF regs_200 ( // @[RegFile.scala 66:20:@37056.4]
    .clock(regs_200_clock),
    .reset(regs_200_reset),
    .io_in(regs_200_io_in),
    .io_reset(regs_200_io_reset),
    .io_out(regs_200_io_out),
    .io_enable(regs_200_io_enable)
  );
  FringeFF regs_201 ( // @[RegFile.scala 66:20:@37070.4]
    .clock(regs_201_clock),
    .reset(regs_201_reset),
    .io_in(regs_201_io_in),
    .io_reset(regs_201_io_reset),
    .io_out(regs_201_io_out),
    .io_enable(regs_201_io_enable)
  );
  FringeFF regs_202 ( // @[RegFile.scala 66:20:@37084.4]
    .clock(regs_202_clock),
    .reset(regs_202_reset),
    .io_in(regs_202_io_in),
    .io_reset(regs_202_io_reset),
    .io_out(regs_202_io_out),
    .io_enable(regs_202_io_enable)
  );
  FringeFF regs_203 ( // @[RegFile.scala 66:20:@37098.4]
    .clock(regs_203_clock),
    .reset(regs_203_reset),
    .io_in(regs_203_io_in),
    .io_reset(regs_203_io_reset),
    .io_out(regs_203_io_out),
    .io_enable(regs_203_io_enable)
  );
  FringeFF regs_204 ( // @[RegFile.scala 66:20:@37112.4]
    .clock(regs_204_clock),
    .reset(regs_204_reset),
    .io_in(regs_204_io_in),
    .io_reset(regs_204_io_reset),
    .io_out(regs_204_io_out),
    .io_enable(regs_204_io_enable)
  );
  FringeFF regs_205 ( // @[RegFile.scala 66:20:@37126.4]
    .clock(regs_205_clock),
    .reset(regs_205_reset),
    .io_in(regs_205_io_in),
    .io_reset(regs_205_io_reset),
    .io_out(regs_205_io_out),
    .io_enable(regs_205_io_enable)
  );
  FringeFF regs_206 ( // @[RegFile.scala 66:20:@37140.4]
    .clock(regs_206_clock),
    .reset(regs_206_reset),
    .io_in(regs_206_io_in),
    .io_reset(regs_206_io_reset),
    .io_out(regs_206_io_out),
    .io_enable(regs_206_io_enable)
  );
  FringeFF regs_207 ( // @[RegFile.scala 66:20:@37154.4]
    .clock(regs_207_clock),
    .reset(regs_207_reset),
    .io_in(regs_207_io_in),
    .io_reset(regs_207_io_reset),
    .io_out(regs_207_io_out),
    .io_enable(regs_207_io_enable)
  );
  FringeFF regs_208 ( // @[RegFile.scala 66:20:@37168.4]
    .clock(regs_208_clock),
    .reset(regs_208_reset),
    .io_in(regs_208_io_in),
    .io_reset(regs_208_io_reset),
    .io_out(regs_208_io_out),
    .io_enable(regs_208_io_enable)
  );
  FringeFF regs_209 ( // @[RegFile.scala 66:20:@37182.4]
    .clock(regs_209_clock),
    .reset(regs_209_reset),
    .io_in(regs_209_io_in),
    .io_reset(regs_209_io_reset),
    .io_out(regs_209_io_out),
    .io_enable(regs_209_io_enable)
  );
  FringeFF regs_210 ( // @[RegFile.scala 66:20:@37196.4]
    .clock(regs_210_clock),
    .reset(regs_210_reset),
    .io_in(regs_210_io_in),
    .io_reset(regs_210_io_reset),
    .io_out(regs_210_io_out),
    .io_enable(regs_210_io_enable)
  );
  FringeFF regs_211 ( // @[RegFile.scala 66:20:@37210.4]
    .clock(regs_211_clock),
    .reset(regs_211_reset),
    .io_in(regs_211_io_in),
    .io_reset(regs_211_io_reset),
    .io_out(regs_211_io_out),
    .io_enable(regs_211_io_enable)
  );
  FringeFF regs_212 ( // @[RegFile.scala 66:20:@37224.4]
    .clock(regs_212_clock),
    .reset(regs_212_reset),
    .io_in(regs_212_io_in),
    .io_reset(regs_212_io_reset),
    .io_out(regs_212_io_out),
    .io_enable(regs_212_io_enable)
  );
  FringeFF regs_213 ( // @[RegFile.scala 66:20:@37238.4]
    .clock(regs_213_clock),
    .reset(regs_213_reset),
    .io_in(regs_213_io_in),
    .io_reset(regs_213_io_reset),
    .io_out(regs_213_io_out),
    .io_enable(regs_213_io_enable)
  );
  FringeFF regs_214 ( // @[RegFile.scala 66:20:@37252.4]
    .clock(regs_214_clock),
    .reset(regs_214_reset),
    .io_in(regs_214_io_in),
    .io_reset(regs_214_io_reset),
    .io_out(regs_214_io_out),
    .io_enable(regs_214_io_enable)
  );
  FringeFF regs_215 ( // @[RegFile.scala 66:20:@37266.4]
    .clock(regs_215_clock),
    .reset(regs_215_reset),
    .io_in(regs_215_io_in),
    .io_reset(regs_215_io_reset),
    .io_out(regs_215_io_out),
    .io_enable(regs_215_io_enable)
  );
  FringeFF regs_216 ( // @[RegFile.scala 66:20:@37280.4]
    .clock(regs_216_clock),
    .reset(regs_216_reset),
    .io_in(regs_216_io_in),
    .io_reset(regs_216_io_reset),
    .io_out(regs_216_io_out),
    .io_enable(regs_216_io_enable)
  );
  FringeFF regs_217 ( // @[RegFile.scala 66:20:@37294.4]
    .clock(regs_217_clock),
    .reset(regs_217_reset),
    .io_in(regs_217_io_in),
    .io_reset(regs_217_io_reset),
    .io_out(regs_217_io_out),
    .io_enable(regs_217_io_enable)
  );
  FringeFF regs_218 ( // @[RegFile.scala 66:20:@37308.4]
    .clock(regs_218_clock),
    .reset(regs_218_reset),
    .io_in(regs_218_io_in),
    .io_reset(regs_218_io_reset),
    .io_out(regs_218_io_out),
    .io_enable(regs_218_io_enable)
  );
  FringeFF regs_219 ( // @[RegFile.scala 66:20:@37322.4]
    .clock(regs_219_clock),
    .reset(regs_219_reset),
    .io_in(regs_219_io_in),
    .io_reset(regs_219_io_reset),
    .io_out(regs_219_io_out),
    .io_enable(regs_219_io_enable)
  );
  FringeFF regs_220 ( // @[RegFile.scala 66:20:@37336.4]
    .clock(regs_220_clock),
    .reset(regs_220_reset),
    .io_in(regs_220_io_in),
    .io_reset(regs_220_io_reset),
    .io_out(regs_220_io_out),
    .io_enable(regs_220_io_enable)
  );
  FringeFF regs_221 ( // @[RegFile.scala 66:20:@37350.4]
    .clock(regs_221_clock),
    .reset(regs_221_reset),
    .io_in(regs_221_io_in),
    .io_reset(regs_221_io_reset),
    .io_out(regs_221_io_out),
    .io_enable(regs_221_io_enable)
  );
  FringeFF regs_222 ( // @[RegFile.scala 66:20:@37364.4]
    .clock(regs_222_clock),
    .reset(regs_222_reset),
    .io_in(regs_222_io_in),
    .io_reset(regs_222_io_reset),
    .io_out(regs_222_io_out),
    .io_enable(regs_222_io_enable)
  );
  FringeFF regs_223 ( // @[RegFile.scala 66:20:@37378.4]
    .clock(regs_223_clock),
    .reset(regs_223_reset),
    .io_in(regs_223_io_in),
    .io_reset(regs_223_io_reset),
    .io_out(regs_223_io_out),
    .io_enable(regs_223_io_enable)
  );
  FringeFF regs_224 ( // @[RegFile.scala 66:20:@37392.4]
    .clock(regs_224_clock),
    .reset(regs_224_reset),
    .io_in(regs_224_io_in),
    .io_reset(regs_224_io_reset),
    .io_out(regs_224_io_out),
    .io_enable(regs_224_io_enable)
  );
  FringeFF regs_225 ( // @[RegFile.scala 66:20:@37406.4]
    .clock(regs_225_clock),
    .reset(regs_225_reset),
    .io_in(regs_225_io_in),
    .io_reset(regs_225_io_reset),
    .io_out(regs_225_io_out),
    .io_enable(regs_225_io_enable)
  );
  FringeFF regs_226 ( // @[RegFile.scala 66:20:@37420.4]
    .clock(regs_226_clock),
    .reset(regs_226_reset),
    .io_in(regs_226_io_in),
    .io_reset(regs_226_io_reset),
    .io_out(regs_226_io_out),
    .io_enable(regs_226_io_enable)
  );
  FringeFF regs_227 ( // @[RegFile.scala 66:20:@37434.4]
    .clock(regs_227_clock),
    .reset(regs_227_reset),
    .io_in(regs_227_io_in),
    .io_reset(regs_227_io_reset),
    .io_out(regs_227_io_out),
    .io_enable(regs_227_io_enable)
  );
  FringeFF regs_228 ( // @[RegFile.scala 66:20:@37448.4]
    .clock(regs_228_clock),
    .reset(regs_228_reset),
    .io_in(regs_228_io_in),
    .io_reset(regs_228_io_reset),
    .io_out(regs_228_io_out),
    .io_enable(regs_228_io_enable)
  );
  FringeFF regs_229 ( // @[RegFile.scala 66:20:@37462.4]
    .clock(regs_229_clock),
    .reset(regs_229_reset),
    .io_in(regs_229_io_in),
    .io_reset(regs_229_io_reset),
    .io_out(regs_229_io_out),
    .io_enable(regs_229_io_enable)
  );
  FringeFF regs_230 ( // @[RegFile.scala 66:20:@37476.4]
    .clock(regs_230_clock),
    .reset(regs_230_reset),
    .io_in(regs_230_io_in),
    .io_reset(regs_230_io_reset),
    .io_out(regs_230_io_out),
    .io_enable(regs_230_io_enable)
  );
  FringeFF regs_231 ( // @[RegFile.scala 66:20:@37490.4]
    .clock(regs_231_clock),
    .reset(regs_231_reset),
    .io_in(regs_231_io_in),
    .io_reset(regs_231_io_reset),
    .io_out(regs_231_io_out),
    .io_enable(regs_231_io_enable)
  );
  FringeFF regs_232 ( // @[RegFile.scala 66:20:@37504.4]
    .clock(regs_232_clock),
    .reset(regs_232_reset),
    .io_in(regs_232_io_in),
    .io_reset(regs_232_io_reset),
    .io_out(regs_232_io_out),
    .io_enable(regs_232_io_enable)
  );
  FringeFF regs_233 ( // @[RegFile.scala 66:20:@37518.4]
    .clock(regs_233_clock),
    .reset(regs_233_reset),
    .io_in(regs_233_io_in),
    .io_reset(regs_233_io_reset),
    .io_out(regs_233_io_out),
    .io_enable(regs_233_io_enable)
  );
  FringeFF regs_234 ( // @[RegFile.scala 66:20:@37532.4]
    .clock(regs_234_clock),
    .reset(regs_234_reset),
    .io_in(regs_234_io_in),
    .io_reset(regs_234_io_reset),
    .io_out(regs_234_io_out),
    .io_enable(regs_234_io_enable)
  );
  FringeFF regs_235 ( // @[RegFile.scala 66:20:@37546.4]
    .clock(regs_235_clock),
    .reset(regs_235_reset),
    .io_in(regs_235_io_in),
    .io_reset(regs_235_io_reset),
    .io_out(regs_235_io_out),
    .io_enable(regs_235_io_enable)
  );
  FringeFF regs_236 ( // @[RegFile.scala 66:20:@37560.4]
    .clock(regs_236_clock),
    .reset(regs_236_reset),
    .io_in(regs_236_io_in),
    .io_reset(regs_236_io_reset),
    .io_out(regs_236_io_out),
    .io_enable(regs_236_io_enable)
  );
  FringeFF regs_237 ( // @[RegFile.scala 66:20:@37574.4]
    .clock(regs_237_clock),
    .reset(regs_237_reset),
    .io_in(regs_237_io_in),
    .io_reset(regs_237_io_reset),
    .io_out(regs_237_io_out),
    .io_enable(regs_237_io_enable)
  );
  FringeFF regs_238 ( // @[RegFile.scala 66:20:@37588.4]
    .clock(regs_238_clock),
    .reset(regs_238_reset),
    .io_in(regs_238_io_in),
    .io_reset(regs_238_io_reset),
    .io_out(regs_238_io_out),
    .io_enable(regs_238_io_enable)
  );
  FringeFF regs_239 ( // @[RegFile.scala 66:20:@37602.4]
    .clock(regs_239_clock),
    .reset(regs_239_reset),
    .io_in(regs_239_io_in),
    .io_reset(regs_239_io_reset),
    .io_out(regs_239_io_out),
    .io_enable(regs_239_io_enable)
  );
  FringeFF regs_240 ( // @[RegFile.scala 66:20:@37616.4]
    .clock(regs_240_clock),
    .reset(regs_240_reset),
    .io_in(regs_240_io_in),
    .io_reset(regs_240_io_reset),
    .io_out(regs_240_io_out),
    .io_enable(regs_240_io_enable)
  );
  FringeFF regs_241 ( // @[RegFile.scala 66:20:@37630.4]
    .clock(regs_241_clock),
    .reset(regs_241_reset),
    .io_in(regs_241_io_in),
    .io_reset(regs_241_io_reset),
    .io_out(regs_241_io_out),
    .io_enable(regs_241_io_enable)
  );
  FringeFF regs_242 ( // @[RegFile.scala 66:20:@37644.4]
    .clock(regs_242_clock),
    .reset(regs_242_reset),
    .io_in(regs_242_io_in),
    .io_reset(regs_242_io_reset),
    .io_out(regs_242_io_out),
    .io_enable(regs_242_io_enable)
  );
  FringeFF regs_243 ( // @[RegFile.scala 66:20:@37658.4]
    .clock(regs_243_clock),
    .reset(regs_243_reset),
    .io_in(regs_243_io_in),
    .io_reset(regs_243_io_reset),
    .io_out(regs_243_io_out),
    .io_enable(regs_243_io_enable)
  );
  FringeFF regs_244 ( // @[RegFile.scala 66:20:@37672.4]
    .clock(regs_244_clock),
    .reset(regs_244_reset),
    .io_in(regs_244_io_in),
    .io_reset(regs_244_io_reset),
    .io_out(regs_244_io_out),
    .io_enable(regs_244_io_enable)
  );
  FringeFF regs_245 ( // @[RegFile.scala 66:20:@37686.4]
    .clock(regs_245_clock),
    .reset(regs_245_reset),
    .io_in(regs_245_io_in),
    .io_reset(regs_245_io_reset),
    .io_out(regs_245_io_out),
    .io_enable(regs_245_io_enable)
  );
  FringeFF regs_246 ( // @[RegFile.scala 66:20:@37700.4]
    .clock(regs_246_clock),
    .reset(regs_246_reset),
    .io_in(regs_246_io_in),
    .io_reset(regs_246_io_reset),
    .io_out(regs_246_io_out),
    .io_enable(regs_246_io_enable)
  );
  FringeFF regs_247 ( // @[RegFile.scala 66:20:@37714.4]
    .clock(regs_247_clock),
    .reset(regs_247_reset),
    .io_in(regs_247_io_in),
    .io_reset(regs_247_io_reset),
    .io_out(regs_247_io_out),
    .io_enable(regs_247_io_enable)
  );
  FringeFF regs_248 ( // @[RegFile.scala 66:20:@37728.4]
    .clock(regs_248_clock),
    .reset(regs_248_reset),
    .io_in(regs_248_io_in),
    .io_reset(regs_248_io_reset),
    .io_out(regs_248_io_out),
    .io_enable(regs_248_io_enable)
  );
  FringeFF regs_249 ( // @[RegFile.scala 66:20:@37742.4]
    .clock(regs_249_clock),
    .reset(regs_249_reset),
    .io_in(regs_249_io_in),
    .io_reset(regs_249_io_reset),
    .io_out(regs_249_io_out),
    .io_enable(regs_249_io_enable)
  );
  FringeFF regs_250 ( // @[RegFile.scala 66:20:@37756.4]
    .clock(regs_250_clock),
    .reset(regs_250_reset),
    .io_in(regs_250_io_in),
    .io_reset(regs_250_io_reset),
    .io_out(regs_250_io_out),
    .io_enable(regs_250_io_enable)
  );
  FringeFF regs_251 ( // @[RegFile.scala 66:20:@37770.4]
    .clock(regs_251_clock),
    .reset(regs_251_reset),
    .io_in(regs_251_io_in),
    .io_reset(regs_251_io_reset),
    .io_out(regs_251_io_out),
    .io_enable(regs_251_io_enable)
  );
  FringeFF regs_252 ( // @[RegFile.scala 66:20:@37784.4]
    .clock(regs_252_clock),
    .reset(regs_252_reset),
    .io_in(regs_252_io_in),
    .io_reset(regs_252_io_reset),
    .io_out(regs_252_io_out),
    .io_enable(regs_252_io_enable)
  );
  FringeFF regs_253 ( // @[RegFile.scala 66:20:@37798.4]
    .clock(regs_253_clock),
    .reset(regs_253_reset),
    .io_in(regs_253_io_in),
    .io_reset(regs_253_io_reset),
    .io_out(regs_253_io_out),
    .io_enable(regs_253_io_enable)
  );
  FringeFF regs_254 ( // @[RegFile.scala 66:20:@37812.4]
    .clock(regs_254_clock),
    .reset(regs_254_reset),
    .io_in(regs_254_io_in),
    .io_reset(regs_254_io_reset),
    .io_out(regs_254_io_out),
    .io_enable(regs_254_io_enable)
  );
  FringeFF regs_255 ( // @[RegFile.scala 66:20:@37826.4]
    .clock(regs_255_clock),
    .reset(regs_255_reset),
    .io_in(regs_255_io_in),
    .io_reset(regs_255_io_reset),
    .io_out(regs_255_io_out),
    .io_enable(regs_255_io_enable)
  );
  FringeFF regs_256 ( // @[RegFile.scala 66:20:@37840.4]
    .clock(regs_256_clock),
    .reset(regs_256_reset),
    .io_in(regs_256_io_in),
    .io_reset(regs_256_io_reset),
    .io_out(regs_256_io_out),
    .io_enable(regs_256_io_enable)
  );
  FringeFF regs_257 ( // @[RegFile.scala 66:20:@37854.4]
    .clock(regs_257_clock),
    .reset(regs_257_reset),
    .io_in(regs_257_io_in),
    .io_reset(regs_257_io_reset),
    .io_out(regs_257_io_out),
    .io_enable(regs_257_io_enable)
  );
  FringeFF regs_258 ( // @[RegFile.scala 66:20:@37868.4]
    .clock(regs_258_clock),
    .reset(regs_258_reset),
    .io_in(regs_258_io_in),
    .io_reset(regs_258_io_reset),
    .io_out(regs_258_io_out),
    .io_enable(regs_258_io_enable)
  );
  FringeFF regs_259 ( // @[RegFile.scala 66:20:@37882.4]
    .clock(regs_259_clock),
    .reset(regs_259_reset),
    .io_in(regs_259_io_in),
    .io_reset(regs_259_io_reset),
    .io_out(regs_259_io_out),
    .io_enable(regs_259_io_enable)
  );
  FringeFF regs_260 ( // @[RegFile.scala 66:20:@37896.4]
    .clock(regs_260_clock),
    .reset(regs_260_reset),
    .io_in(regs_260_io_in),
    .io_reset(regs_260_io_reset),
    .io_out(regs_260_io_out),
    .io_enable(regs_260_io_enable)
  );
  FringeFF regs_261 ( // @[RegFile.scala 66:20:@37910.4]
    .clock(regs_261_clock),
    .reset(regs_261_reset),
    .io_in(regs_261_io_in),
    .io_reset(regs_261_io_reset),
    .io_out(regs_261_io_out),
    .io_enable(regs_261_io_enable)
  );
  FringeFF regs_262 ( // @[RegFile.scala 66:20:@37924.4]
    .clock(regs_262_clock),
    .reset(regs_262_reset),
    .io_in(regs_262_io_in),
    .io_reset(regs_262_io_reset),
    .io_out(regs_262_io_out),
    .io_enable(regs_262_io_enable)
  );
  FringeFF regs_263 ( // @[RegFile.scala 66:20:@37938.4]
    .clock(regs_263_clock),
    .reset(regs_263_reset),
    .io_in(regs_263_io_in),
    .io_reset(regs_263_io_reset),
    .io_out(regs_263_io_out),
    .io_enable(regs_263_io_enable)
  );
  FringeFF regs_264 ( // @[RegFile.scala 66:20:@37952.4]
    .clock(regs_264_clock),
    .reset(regs_264_reset),
    .io_in(regs_264_io_in),
    .io_reset(regs_264_io_reset),
    .io_out(regs_264_io_out),
    .io_enable(regs_264_io_enable)
  );
  FringeFF regs_265 ( // @[RegFile.scala 66:20:@37966.4]
    .clock(regs_265_clock),
    .reset(regs_265_reset),
    .io_in(regs_265_io_in),
    .io_reset(regs_265_io_reset),
    .io_out(regs_265_io_out),
    .io_enable(regs_265_io_enable)
  );
  FringeFF regs_266 ( // @[RegFile.scala 66:20:@37980.4]
    .clock(regs_266_clock),
    .reset(regs_266_reset),
    .io_in(regs_266_io_in),
    .io_reset(regs_266_io_reset),
    .io_out(regs_266_io_out),
    .io_enable(regs_266_io_enable)
  );
  FringeFF regs_267 ( // @[RegFile.scala 66:20:@37994.4]
    .clock(regs_267_clock),
    .reset(regs_267_reset),
    .io_in(regs_267_io_in),
    .io_reset(regs_267_io_reset),
    .io_out(regs_267_io_out),
    .io_enable(regs_267_io_enable)
  );
  FringeFF regs_268 ( // @[RegFile.scala 66:20:@38008.4]
    .clock(regs_268_clock),
    .reset(regs_268_reset),
    .io_in(regs_268_io_in),
    .io_reset(regs_268_io_reset),
    .io_out(regs_268_io_out),
    .io_enable(regs_268_io_enable)
  );
  FringeFF regs_269 ( // @[RegFile.scala 66:20:@38022.4]
    .clock(regs_269_clock),
    .reset(regs_269_reset),
    .io_in(regs_269_io_in),
    .io_reset(regs_269_io_reset),
    .io_out(regs_269_io_out),
    .io_enable(regs_269_io_enable)
  );
  FringeFF regs_270 ( // @[RegFile.scala 66:20:@38036.4]
    .clock(regs_270_clock),
    .reset(regs_270_reset),
    .io_in(regs_270_io_in),
    .io_reset(regs_270_io_reset),
    .io_out(regs_270_io_out),
    .io_enable(regs_270_io_enable)
  );
  FringeFF regs_271 ( // @[RegFile.scala 66:20:@38050.4]
    .clock(regs_271_clock),
    .reset(regs_271_reset),
    .io_in(regs_271_io_in),
    .io_reset(regs_271_io_reset),
    .io_out(regs_271_io_out),
    .io_enable(regs_271_io_enable)
  );
  FringeFF regs_272 ( // @[RegFile.scala 66:20:@38064.4]
    .clock(regs_272_clock),
    .reset(regs_272_reset),
    .io_in(regs_272_io_in),
    .io_reset(regs_272_io_reset),
    .io_out(regs_272_io_out),
    .io_enable(regs_272_io_enable)
  );
  FringeFF regs_273 ( // @[RegFile.scala 66:20:@38078.4]
    .clock(regs_273_clock),
    .reset(regs_273_reset),
    .io_in(regs_273_io_in),
    .io_reset(regs_273_io_reset),
    .io_out(regs_273_io_out),
    .io_enable(regs_273_io_enable)
  );
  FringeFF regs_274 ( // @[RegFile.scala 66:20:@38092.4]
    .clock(regs_274_clock),
    .reset(regs_274_reset),
    .io_in(regs_274_io_in),
    .io_reset(regs_274_io_reset),
    .io_out(regs_274_io_out),
    .io_enable(regs_274_io_enable)
  );
  FringeFF regs_275 ( // @[RegFile.scala 66:20:@38106.4]
    .clock(regs_275_clock),
    .reset(regs_275_reset),
    .io_in(regs_275_io_in),
    .io_reset(regs_275_io_reset),
    .io_out(regs_275_io_out),
    .io_enable(regs_275_io_enable)
  );
  FringeFF regs_276 ( // @[RegFile.scala 66:20:@38120.4]
    .clock(regs_276_clock),
    .reset(regs_276_reset),
    .io_in(regs_276_io_in),
    .io_reset(regs_276_io_reset),
    .io_out(regs_276_io_out),
    .io_enable(regs_276_io_enable)
  );
  FringeFF regs_277 ( // @[RegFile.scala 66:20:@38134.4]
    .clock(regs_277_clock),
    .reset(regs_277_reset),
    .io_in(regs_277_io_in),
    .io_reset(regs_277_io_reset),
    .io_out(regs_277_io_out),
    .io_enable(regs_277_io_enable)
  );
  FringeFF regs_278 ( // @[RegFile.scala 66:20:@38148.4]
    .clock(regs_278_clock),
    .reset(regs_278_reset),
    .io_in(regs_278_io_in),
    .io_reset(regs_278_io_reset),
    .io_out(regs_278_io_out),
    .io_enable(regs_278_io_enable)
  );
  FringeFF regs_279 ( // @[RegFile.scala 66:20:@38162.4]
    .clock(regs_279_clock),
    .reset(regs_279_reset),
    .io_in(regs_279_io_in),
    .io_reset(regs_279_io_reset),
    .io_out(regs_279_io_out),
    .io_enable(regs_279_io_enable)
  );
  FringeFF regs_280 ( // @[RegFile.scala 66:20:@38176.4]
    .clock(regs_280_clock),
    .reset(regs_280_reset),
    .io_in(regs_280_io_in),
    .io_reset(regs_280_io_reset),
    .io_out(regs_280_io_out),
    .io_enable(regs_280_io_enable)
  );
  FringeFF regs_281 ( // @[RegFile.scala 66:20:@38190.4]
    .clock(regs_281_clock),
    .reset(regs_281_reset),
    .io_in(regs_281_io_in),
    .io_reset(regs_281_io_reset),
    .io_out(regs_281_io_out),
    .io_enable(regs_281_io_enable)
  );
  FringeFF regs_282 ( // @[RegFile.scala 66:20:@38204.4]
    .clock(regs_282_clock),
    .reset(regs_282_reset),
    .io_in(regs_282_io_in),
    .io_reset(regs_282_io_reset),
    .io_out(regs_282_io_out),
    .io_enable(regs_282_io_enable)
  );
  FringeFF regs_283 ( // @[RegFile.scala 66:20:@38218.4]
    .clock(regs_283_clock),
    .reset(regs_283_reset),
    .io_in(regs_283_io_in),
    .io_reset(regs_283_io_reset),
    .io_out(regs_283_io_out),
    .io_enable(regs_283_io_enable)
  );
  FringeFF regs_284 ( // @[RegFile.scala 66:20:@38232.4]
    .clock(regs_284_clock),
    .reset(regs_284_reset),
    .io_in(regs_284_io_in),
    .io_reset(regs_284_io_reset),
    .io_out(regs_284_io_out),
    .io_enable(regs_284_io_enable)
  );
  FringeFF regs_285 ( // @[RegFile.scala 66:20:@38246.4]
    .clock(regs_285_clock),
    .reset(regs_285_reset),
    .io_in(regs_285_io_in),
    .io_reset(regs_285_io_reset),
    .io_out(regs_285_io_out),
    .io_enable(regs_285_io_enable)
  );
  FringeFF regs_286 ( // @[RegFile.scala 66:20:@38260.4]
    .clock(regs_286_clock),
    .reset(regs_286_reset),
    .io_in(regs_286_io_in),
    .io_reset(regs_286_io_reset),
    .io_out(regs_286_io_out),
    .io_enable(regs_286_io_enable)
  );
  FringeFF regs_287 ( // @[RegFile.scala 66:20:@38274.4]
    .clock(regs_287_clock),
    .reset(regs_287_reset),
    .io_in(regs_287_io_in),
    .io_reset(regs_287_io_reset),
    .io_out(regs_287_io_out),
    .io_enable(regs_287_io_enable)
  );
  FringeFF regs_288 ( // @[RegFile.scala 66:20:@38288.4]
    .clock(regs_288_clock),
    .reset(regs_288_reset),
    .io_in(regs_288_io_in),
    .io_reset(regs_288_io_reset),
    .io_out(regs_288_io_out),
    .io_enable(regs_288_io_enable)
  );
  FringeFF regs_289 ( // @[RegFile.scala 66:20:@38302.4]
    .clock(regs_289_clock),
    .reset(regs_289_reset),
    .io_in(regs_289_io_in),
    .io_reset(regs_289_io_reset),
    .io_out(regs_289_io_out),
    .io_enable(regs_289_io_enable)
  );
  FringeFF regs_290 ( // @[RegFile.scala 66:20:@38316.4]
    .clock(regs_290_clock),
    .reset(regs_290_reset),
    .io_in(regs_290_io_in),
    .io_reset(regs_290_io_reset),
    .io_out(regs_290_io_out),
    .io_enable(regs_290_io_enable)
  );
  FringeFF regs_291 ( // @[RegFile.scala 66:20:@38330.4]
    .clock(regs_291_clock),
    .reset(regs_291_reset),
    .io_in(regs_291_io_in),
    .io_reset(regs_291_io_reset),
    .io_out(regs_291_io_out),
    .io_enable(regs_291_io_enable)
  );
  FringeFF regs_292 ( // @[RegFile.scala 66:20:@38344.4]
    .clock(regs_292_clock),
    .reset(regs_292_reset),
    .io_in(regs_292_io_in),
    .io_reset(regs_292_io_reset),
    .io_out(regs_292_io_out),
    .io_enable(regs_292_io_enable)
  );
  FringeFF regs_293 ( // @[RegFile.scala 66:20:@38358.4]
    .clock(regs_293_clock),
    .reset(regs_293_reset),
    .io_in(regs_293_io_in),
    .io_reset(regs_293_io_reset),
    .io_out(regs_293_io_out),
    .io_enable(regs_293_io_enable)
  );
  FringeFF regs_294 ( // @[RegFile.scala 66:20:@38372.4]
    .clock(regs_294_clock),
    .reset(regs_294_reset),
    .io_in(regs_294_io_in),
    .io_reset(regs_294_io_reset),
    .io_out(regs_294_io_out),
    .io_enable(regs_294_io_enable)
  );
  FringeFF regs_295 ( // @[RegFile.scala 66:20:@38386.4]
    .clock(regs_295_clock),
    .reset(regs_295_reset),
    .io_in(regs_295_io_in),
    .io_reset(regs_295_io_reset),
    .io_out(regs_295_io_out),
    .io_enable(regs_295_io_enable)
  );
  FringeFF regs_296 ( // @[RegFile.scala 66:20:@38400.4]
    .clock(regs_296_clock),
    .reset(regs_296_reset),
    .io_in(regs_296_io_in),
    .io_reset(regs_296_io_reset),
    .io_out(regs_296_io_out),
    .io_enable(regs_296_io_enable)
  );
  FringeFF regs_297 ( // @[RegFile.scala 66:20:@38414.4]
    .clock(regs_297_clock),
    .reset(regs_297_reset),
    .io_in(regs_297_io_in),
    .io_reset(regs_297_io_reset),
    .io_out(regs_297_io_out),
    .io_enable(regs_297_io_enable)
  );
  FringeFF regs_298 ( // @[RegFile.scala 66:20:@38428.4]
    .clock(regs_298_clock),
    .reset(regs_298_reset),
    .io_in(regs_298_io_in),
    .io_reset(regs_298_io_reset),
    .io_out(regs_298_io_out),
    .io_enable(regs_298_io_enable)
  );
  FringeFF regs_299 ( // @[RegFile.scala 66:20:@38442.4]
    .clock(regs_299_clock),
    .reset(regs_299_reset),
    .io_in(regs_299_io_in),
    .io_reset(regs_299_io_reset),
    .io_out(regs_299_io_out),
    .io_enable(regs_299_io_enable)
  );
  FringeFF regs_300 ( // @[RegFile.scala 66:20:@38456.4]
    .clock(regs_300_clock),
    .reset(regs_300_reset),
    .io_in(regs_300_io_in),
    .io_reset(regs_300_io_reset),
    .io_out(regs_300_io_out),
    .io_enable(regs_300_io_enable)
  );
  FringeFF regs_301 ( // @[RegFile.scala 66:20:@38470.4]
    .clock(regs_301_clock),
    .reset(regs_301_reset),
    .io_in(regs_301_io_in),
    .io_reset(regs_301_io_reset),
    .io_out(regs_301_io_out),
    .io_enable(regs_301_io_enable)
  );
  FringeFF regs_302 ( // @[RegFile.scala 66:20:@38484.4]
    .clock(regs_302_clock),
    .reset(regs_302_reset),
    .io_in(regs_302_io_in),
    .io_reset(regs_302_io_reset),
    .io_out(regs_302_io_out),
    .io_enable(regs_302_io_enable)
  );
  FringeFF regs_303 ( // @[RegFile.scala 66:20:@38498.4]
    .clock(regs_303_clock),
    .reset(regs_303_reset),
    .io_in(regs_303_io_in),
    .io_reset(regs_303_io_reset),
    .io_out(regs_303_io_out),
    .io_enable(regs_303_io_enable)
  );
  FringeFF regs_304 ( // @[RegFile.scala 66:20:@38512.4]
    .clock(regs_304_clock),
    .reset(regs_304_reset),
    .io_in(regs_304_io_in),
    .io_reset(regs_304_io_reset),
    .io_out(regs_304_io_out),
    .io_enable(regs_304_io_enable)
  );
  FringeFF regs_305 ( // @[RegFile.scala 66:20:@38526.4]
    .clock(regs_305_clock),
    .reset(regs_305_reset),
    .io_in(regs_305_io_in),
    .io_reset(regs_305_io_reset),
    .io_out(regs_305_io_out),
    .io_enable(regs_305_io_enable)
  );
  FringeFF regs_306 ( // @[RegFile.scala 66:20:@38540.4]
    .clock(regs_306_clock),
    .reset(regs_306_reset),
    .io_in(regs_306_io_in),
    .io_reset(regs_306_io_reset),
    .io_out(regs_306_io_out),
    .io_enable(regs_306_io_enable)
  );
  FringeFF regs_307 ( // @[RegFile.scala 66:20:@38554.4]
    .clock(regs_307_clock),
    .reset(regs_307_reset),
    .io_in(regs_307_io_in),
    .io_reset(regs_307_io_reset),
    .io_out(regs_307_io_out),
    .io_enable(regs_307_io_enable)
  );
  FringeFF regs_308 ( // @[RegFile.scala 66:20:@38568.4]
    .clock(regs_308_clock),
    .reset(regs_308_reset),
    .io_in(regs_308_io_in),
    .io_reset(regs_308_io_reset),
    .io_out(regs_308_io_out),
    .io_enable(regs_308_io_enable)
  );
  FringeFF regs_309 ( // @[RegFile.scala 66:20:@38582.4]
    .clock(regs_309_clock),
    .reset(regs_309_reset),
    .io_in(regs_309_io_in),
    .io_reset(regs_309_io_reset),
    .io_out(regs_309_io_out),
    .io_enable(regs_309_io_enable)
  );
  FringeFF regs_310 ( // @[RegFile.scala 66:20:@38596.4]
    .clock(regs_310_clock),
    .reset(regs_310_reset),
    .io_in(regs_310_io_in),
    .io_reset(regs_310_io_reset),
    .io_out(regs_310_io_out),
    .io_enable(regs_310_io_enable)
  );
  FringeFF regs_311 ( // @[RegFile.scala 66:20:@38610.4]
    .clock(regs_311_clock),
    .reset(regs_311_reset),
    .io_in(regs_311_io_in),
    .io_reset(regs_311_io_reset),
    .io_out(regs_311_io_out),
    .io_enable(regs_311_io_enable)
  );
  FringeFF regs_312 ( // @[RegFile.scala 66:20:@38624.4]
    .clock(regs_312_clock),
    .reset(regs_312_reset),
    .io_in(regs_312_io_in),
    .io_reset(regs_312_io_reset),
    .io_out(regs_312_io_out),
    .io_enable(regs_312_io_enable)
  );
  FringeFF regs_313 ( // @[RegFile.scala 66:20:@38638.4]
    .clock(regs_313_clock),
    .reset(regs_313_reset),
    .io_in(regs_313_io_in),
    .io_reset(regs_313_io_reset),
    .io_out(regs_313_io_out),
    .io_enable(regs_313_io_enable)
  );
  FringeFF regs_314 ( // @[RegFile.scala 66:20:@38652.4]
    .clock(regs_314_clock),
    .reset(regs_314_reset),
    .io_in(regs_314_io_in),
    .io_reset(regs_314_io_reset),
    .io_out(regs_314_io_out),
    .io_enable(regs_314_io_enable)
  );
  FringeFF regs_315 ( // @[RegFile.scala 66:20:@38666.4]
    .clock(regs_315_clock),
    .reset(regs_315_reset),
    .io_in(regs_315_io_in),
    .io_reset(regs_315_io_reset),
    .io_out(regs_315_io_out),
    .io_enable(regs_315_io_enable)
  );
  FringeFF regs_316 ( // @[RegFile.scala 66:20:@38680.4]
    .clock(regs_316_clock),
    .reset(regs_316_reset),
    .io_in(regs_316_io_in),
    .io_reset(regs_316_io_reset),
    .io_out(regs_316_io_out),
    .io_enable(regs_316_io_enable)
  );
  FringeFF regs_317 ( // @[RegFile.scala 66:20:@38694.4]
    .clock(regs_317_clock),
    .reset(regs_317_reset),
    .io_in(regs_317_io_in),
    .io_reset(regs_317_io_reset),
    .io_out(regs_317_io_out),
    .io_enable(regs_317_io_enable)
  );
  FringeFF regs_318 ( // @[RegFile.scala 66:20:@38708.4]
    .clock(regs_318_clock),
    .reset(regs_318_reset),
    .io_in(regs_318_io_in),
    .io_reset(regs_318_io_reset),
    .io_out(regs_318_io_out),
    .io_enable(regs_318_io_enable)
  );
  FringeFF regs_319 ( // @[RegFile.scala 66:20:@38722.4]
    .clock(regs_319_clock),
    .reset(regs_319_reset),
    .io_in(regs_319_io_in),
    .io_reset(regs_319_io_reset),
    .io_out(regs_319_io_out),
    .io_enable(regs_319_io_enable)
  );
  FringeFF regs_320 ( // @[RegFile.scala 66:20:@38736.4]
    .clock(regs_320_clock),
    .reset(regs_320_reset),
    .io_in(regs_320_io_in),
    .io_reset(regs_320_io_reset),
    .io_out(regs_320_io_out),
    .io_enable(regs_320_io_enable)
  );
  FringeFF regs_321 ( // @[RegFile.scala 66:20:@38750.4]
    .clock(regs_321_clock),
    .reset(regs_321_reset),
    .io_in(regs_321_io_in),
    .io_reset(regs_321_io_reset),
    .io_out(regs_321_io_out),
    .io_enable(regs_321_io_enable)
  );
  FringeFF regs_322 ( // @[RegFile.scala 66:20:@38764.4]
    .clock(regs_322_clock),
    .reset(regs_322_reset),
    .io_in(regs_322_io_in),
    .io_reset(regs_322_io_reset),
    .io_out(regs_322_io_out),
    .io_enable(regs_322_io_enable)
  );
  FringeFF regs_323 ( // @[RegFile.scala 66:20:@38778.4]
    .clock(regs_323_clock),
    .reset(regs_323_reset),
    .io_in(regs_323_io_in),
    .io_reset(regs_323_io_reset),
    .io_out(regs_323_io_out),
    .io_enable(regs_323_io_enable)
  );
  FringeFF regs_324 ( // @[RegFile.scala 66:20:@38792.4]
    .clock(regs_324_clock),
    .reset(regs_324_reset),
    .io_in(regs_324_io_in),
    .io_reset(regs_324_io_reset),
    .io_out(regs_324_io_out),
    .io_enable(regs_324_io_enable)
  );
  FringeFF regs_325 ( // @[RegFile.scala 66:20:@38806.4]
    .clock(regs_325_clock),
    .reset(regs_325_reset),
    .io_in(regs_325_io_in),
    .io_reset(regs_325_io_reset),
    .io_out(regs_325_io_out),
    .io_enable(regs_325_io_enable)
  );
  FringeFF regs_326 ( // @[RegFile.scala 66:20:@38820.4]
    .clock(regs_326_clock),
    .reset(regs_326_reset),
    .io_in(regs_326_io_in),
    .io_reset(regs_326_io_reset),
    .io_out(regs_326_io_out),
    .io_enable(regs_326_io_enable)
  );
  FringeFF regs_327 ( // @[RegFile.scala 66:20:@38834.4]
    .clock(regs_327_clock),
    .reset(regs_327_reset),
    .io_in(regs_327_io_in),
    .io_reset(regs_327_io_reset),
    .io_out(regs_327_io_out),
    .io_enable(regs_327_io_enable)
  );
  FringeFF regs_328 ( // @[RegFile.scala 66:20:@38848.4]
    .clock(regs_328_clock),
    .reset(regs_328_reset),
    .io_in(regs_328_io_in),
    .io_reset(regs_328_io_reset),
    .io_out(regs_328_io_out),
    .io_enable(regs_328_io_enable)
  );
  FringeFF regs_329 ( // @[RegFile.scala 66:20:@38862.4]
    .clock(regs_329_clock),
    .reset(regs_329_reset),
    .io_in(regs_329_io_in),
    .io_reset(regs_329_io_reset),
    .io_out(regs_329_io_out),
    .io_enable(regs_329_io_enable)
  );
  FringeFF regs_330 ( // @[RegFile.scala 66:20:@38876.4]
    .clock(regs_330_clock),
    .reset(regs_330_reset),
    .io_in(regs_330_io_in),
    .io_reset(regs_330_io_reset),
    .io_out(regs_330_io_out),
    .io_enable(regs_330_io_enable)
  );
  FringeFF regs_331 ( // @[RegFile.scala 66:20:@38890.4]
    .clock(regs_331_clock),
    .reset(regs_331_reset),
    .io_in(regs_331_io_in),
    .io_reset(regs_331_io_reset),
    .io_out(regs_331_io_out),
    .io_enable(regs_331_io_enable)
  );
  FringeFF regs_332 ( // @[RegFile.scala 66:20:@38904.4]
    .clock(regs_332_clock),
    .reset(regs_332_reset),
    .io_in(regs_332_io_in),
    .io_reset(regs_332_io_reset),
    .io_out(regs_332_io_out),
    .io_enable(regs_332_io_enable)
  );
  FringeFF regs_333 ( // @[RegFile.scala 66:20:@38918.4]
    .clock(regs_333_clock),
    .reset(regs_333_reset),
    .io_in(regs_333_io_in),
    .io_reset(regs_333_io_reset),
    .io_out(regs_333_io_out),
    .io_enable(regs_333_io_enable)
  );
  FringeFF regs_334 ( // @[RegFile.scala 66:20:@38932.4]
    .clock(regs_334_clock),
    .reset(regs_334_reset),
    .io_in(regs_334_io_in),
    .io_reset(regs_334_io_reset),
    .io_out(regs_334_io_out),
    .io_enable(regs_334_io_enable)
  );
  FringeFF regs_335 ( // @[RegFile.scala 66:20:@38946.4]
    .clock(regs_335_clock),
    .reset(regs_335_reset),
    .io_in(regs_335_io_in),
    .io_reset(regs_335_io_reset),
    .io_out(regs_335_io_out),
    .io_enable(regs_335_io_enable)
  );
  FringeFF regs_336 ( // @[RegFile.scala 66:20:@38960.4]
    .clock(regs_336_clock),
    .reset(regs_336_reset),
    .io_in(regs_336_io_in),
    .io_reset(regs_336_io_reset),
    .io_out(regs_336_io_out),
    .io_enable(regs_336_io_enable)
  );
  FringeFF regs_337 ( // @[RegFile.scala 66:20:@38974.4]
    .clock(regs_337_clock),
    .reset(regs_337_reset),
    .io_in(regs_337_io_in),
    .io_reset(regs_337_io_reset),
    .io_out(regs_337_io_out),
    .io_enable(regs_337_io_enable)
  );
  FringeFF regs_338 ( // @[RegFile.scala 66:20:@38988.4]
    .clock(regs_338_clock),
    .reset(regs_338_reset),
    .io_in(regs_338_io_in),
    .io_reset(regs_338_io_reset),
    .io_out(regs_338_io_out),
    .io_enable(regs_338_io_enable)
  );
  FringeFF regs_339 ( // @[RegFile.scala 66:20:@39002.4]
    .clock(regs_339_clock),
    .reset(regs_339_reset),
    .io_in(regs_339_io_in),
    .io_reset(regs_339_io_reset),
    .io_out(regs_339_io_out),
    .io_enable(regs_339_io_enable)
  );
  FringeFF regs_340 ( // @[RegFile.scala 66:20:@39016.4]
    .clock(regs_340_clock),
    .reset(regs_340_reset),
    .io_in(regs_340_io_in),
    .io_reset(regs_340_io_reset),
    .io_out(regs_340_io_out),
    .io_enable(regs_340_io_enable)
  );
  FringeFF regs_341 ( // @[RegFile.scala 66:20:@39030.4]
    .clock(regs_341_clock),
    .reset(regs_341_reset),
    .io_in(regs_341_io_in),
    .io_reset(regs_341_io_reset),
    .io_out(regs_341_io_out),
    .io_enable(regs_341_io_enable)
  );
  FringeFF regs_342 ( // @[RegFile.scala 66:20:@39044.4]
    .clock(regs_342_clock),
    .reset(regs_342_reset),
    .io_in(regs_342_io_in),
    .io_reset(regs_342_io_reset),
    .io_out(regs_342_io_out),
    .io_enable(regs_342_io_enable)
  );
  FringeFF regs_343 ( // @[RegFile.scala 66:20:@39058.4]
    .clock(regs_343_clock),
    .reset(regs_343_reset),
    .io_in(regs_343_io_in),
    .io_reset(regs_343_io_reset),
    .io_out(regs_343_io_out),
    .io_enable(regs_343_io_enable)
  );
  FringeFF regs_344 ( // @[RegFile.scala 66:20:@39072.4]
    .clock(regs_344_clock),
    .reset(regs_344_reset),
    .io_in(regs_344_io_in),
    .io_reset(regs_344_io_reset),
    .io_out(regs_344_io_out),
    .io_enable(regs_344_io_enable)
  );
  FringeFF regs_345 ( // @[RegFile.scala 66:20:@39086.4]
    .clock(regs_345_clock),
    .reset(regs_345_reset),
    .io_in(regs_345_io_in),
    .io_reset(regs_345_io_reset),
    .io_out(regs_345_io_out),
    .io_enable(regs_345_io_enable)
  );
  FringeFF regs_346 ( // @[RegFile.scala 66:20:@39100.4]
    .clock(regs_346_clock),
    .reset(regs_346_reset),
    .io_in(regs_346_io_in),
    .io_reset(regs_346_io_reset),
    .io_out(regs_346_io_out),
    .io_enable(regs_346_io_enable)
  );
  FringeFF regs_347 ( // @[RegFile.scala 66:20:@39114.4]
    .clock(regs_347_clock),
    .reset(regs_347_reset),
    .io_in(regs_347_io_in),
    .io_reset(regs_347_io_reset),
    .io_out(regs_347_io_out),
    .io_enable(regs_347_io_enable)
  );
  FringeFF regs_348 ( // @[RegFile.scala 66:20:@39128.4]
    .clock(regs_348_clock),
    .reset(regs_348_reset),
    .io_in(regs_348_io_in),
    .io_reset(regs_348_io_reset),
    .io_out(regs_348_io_out),
    .io_enable(regs_348_io_enable)
  );
  FringeFF regs_349 ( // @[RegFile.scala 66:20:@39142.4]
    .clock(regs_349_clock),
    .reset(regs_349_reset),
    .io_in(regs_349_io_in),
    .io_reset(regs_349_io_reset),
    .io_out(regs_349_io_out),
    .io_enable(regs_349_io_enable)
  );
  FringeFF regs_350 ( // @[RegFile.scala 66:20:@39156.4]
    .clock(regs_350_clock),
    .reset(regs_350_reset),
    .io_in(regs_350_io_in),
    .io_reset(regs_350_io_reset),
    .io_out(regs_350_io_out),
    .io_enable(regs_350_io_enable)
  );
  FringeFF regs_351 ( // @[RegFile.scala 66:20:@39170.4]
    .clock(regs_351_clock),
    .reset(regs_351_reset),
    .io_in(regs_351_io_in),
    .io_reset(regs_351_io_reset),
    .io_out(regs_351_io_out),
    .io_enable(regs_351_io_enable)
  );
  FringeFF regs_352 ( // @[RegFile.scala 66:20:@39184.4]
    .clock(regs_352_clock),
    .reset(regs_352_reset),
    .io_in(regs_352_io_in),
    .io_reset(regs_352_io_reset),
    .io_out(regs_352_io_out),
    .io_enable(regs_352_io_enable)
  );
  FringeFF regs_353 ( // @[RegFile.scala 66:20:@39198.4]
    .clock(regs_353_clock),
    .reset(regs_353_reset),
    .io_in(regs_353_io_in),
    .io_reset(regs_353_io_reset),
    .io_out(regs_353_io_out),
    .io_enable(regs_353_io_enable)
  );
  FringeFF regs_354 ( // @[RegFile.scala 66:20:@39212.4]
    .clock(regs_354_clock),
    .reset(regs_354_reset),
    .io_in(regs_354_io_in),
    .io_reset(regs_354_io_reset),
    .io_out(regs_354_io_out),
    .io_enable(regs_354_io_enable)
  );
  FringeFF regs_355 ( // @[RegFile.scala 66:20:@39226.4]
    .clock(regs_355_clock),
    .reset(regs_355_reset),
    .io_in(regs_355_io_in),
    .io_reset(regs_355_io_reset),
    .io_out(regs_355_io_out),
    .io_enable(regs_355_io_enable)
  );
  FringeFF regs_356 ( // @[RegFile.scala 66:20:@39240.4]
    .clock(regs_356_clock),
    .reset(regs_356_reset),
    .io_in(regs_356_io_in),
    .io_reset(regs_356_io_reset),
    .io_out(regs_356_io_out),
    .io_enable(regs_356_io_enable)
  );
  FringeFF regs_357 ( // @[RegFile.scala 66:20:@39254.4]
    .clock(regs_357_clock),
    .reset(regs_357_reset),
    .io_in(regs_357_io_in),
    .io_reset(regs_357_io_reset),
    .io_out(regs_357_io_out),
    .io_enable(regs_357_io_enable)
  );
  FringeFF regs_358 ( // @[RegFile.scala 66:20:@39268.4]
    .clock(regs_358_clock),
    .reset(regs_358_reset),
    .io_in(regs_358_io_in),
    .io_reset(regs_358_io_reset),
    .io_out(regs_358_io_out),
    .io_enable(regs_358_io_enable)
  );
  FringeFF regs_359 ( // @[RegFile.scala 66:20:@39282.4]
    .clock(regs_359_clock),
    .reset(regs_359_reset),
    .io_in(regs_359_io_in),
    .io_reset(regs_359_io_reset),
    .io_out(regs_359_io_out),
    .io_enable(regs_359_io_enable)
  );
  FringeFF regs_360 ( // @[RegFile.scala 66:20:@39296.4]
    .clock(regs_360_clock),
    .reset(regs_360_reset),
    .io_in(regs_360_io_in),
    .io_reset(regs_360_io_reset),
    .io_out(regs_360_io_out),
    .io_enable(regs_360_io_enable)
  );
  FringeFF regs_361 ( // @[RegFile.scala 66:20:@39310.4]
    .clock(regs_361_clock),
    .reset(regs_361_reset),
    .io_in(regs_361_io_in),
    .io_reset(regs_361_io_reset),
    .io_out(regs_361_io_out),
    .io_enable(regs_361_io_enable)
  );
  FringeFF regs_362 ( // @[RegFile.scala 66:20:@39324.4]
    .clock(regs_362_clock),
    .reset(regs_362_reset),
    .io_in(regs_362_io_in),
    .io_reset(regs_362_io_reset),
    .io_out(regs_362_io_out),
    .io_enable(regs_362_io_enable)
  );
  FringeFF regs_363 ( // @[RegFile.scala 66:20:@39338.4]
    .clock(regs_363_clock),
    .reset(regs_363_reset),
    .io_in(regs_363_io_in),
    .io_reset(regs_363_io_reset),
    .io_out(regs_363_io_out),
    .io_enable(regs_363_io_enable)
  );
  FringeFF regs_364 ( // @[RegFile.scala 66:20:@39352.4]
    .clock(regs_364_clock),
    .reset(regs_364_reset),
    .io_in(regs_364_io_in),
    .io_reset(regs_364_io_reset),
    .io_out(regs_364_io_out),
    .io_enable(regs_364_io_enable)
  );
  FringeFF regs_365 ( // @[RegFile.scala 66:20:@39366.4]
    .clock(regs_365_clock),
    .reset(regs_365_reset),
    .io_in(regs_365_io_in),
    .io_reset(regs_365_io_reset),
    .io_out(regs_365_io_out),
    .io_enable(regs_365_io_enable)
  );
  FringeFF regs_366 ( // @[RegFile.scala 66:20:@39380.4]
    .clock(regs_366_clock),
    .reset(regs_366_reset),
    .io_in(regs_366_io_in),
    .io_reset(regs_366_io_reset),
    .io_out(regs_366_io_out),
    .io_enable(regs_366_io_enable)
  );
  FringeFF regs_367 ( // @[RegFile.scala 66:20:@39394.4]
    .clock(regs_367_clock),
    .reset(regs_367_reset),
    .io_in(regs_367_io_in),
    .io_reset(regs_367_io_reset),
    .io_out(regs_367_io_out),
    .io_enable(regs_367_io_enable)
  );
  FringeFF regs_368 ( // @[RegFile.scala 66:20:@39408.4]
    .clock(regs_368_clock),
    .reset(regs_368_reset),
    .io_in(regs_368_io_in),
    .io_reset(regs_368_io_reset),
    .io_out(regs_368_io_out),
    .io_enable(regs_368_io_enable)
  );
  FringeFF regs_369 ( // @[RegFile.scala 66:20:@39422.4]
    .clock(regs_369_clock),
    .reset(regs_369_reset),
    .io_in(regs_369_io_in),
    .io_reset(regs_369_io_reset),
    .io_out(regs_369_io_out),
    .io_enable(regs_369_io_enable)
  );
  FringeFF regs_370 ( // @[RegFile.scala 66:20:@39436.4]
    .clock(regs_370_clock),
    .reset(regs_370_reset),
    .io_in(regs_370_io_in),
    .io_reset(regs_370_io_reset),
    .io_out(regs_370_io_out),
    .io_enable(regs_370_io_enable)
  );
  FringeFF regs_371 ( // @[RegFile.scala 66:20:@39450.4]
    .clock(regs_371_clock),
    .reset(regs_371_reset),
    .io_in(regs_371_io_in),
    .io_reset(regs_371_io_reset),
    .io_out(regs_371_io_out),
    .io_enable(regs_371_io_enable)
  );
  FringeFF regs_372 ( // @[RegFile.scala 66:20:@39464.4]
    .clock(regs_372_clock),
    .reset(regs_372_reset),
    .io_in(regs_372_io_in),
    .io_reset(regs_372_io_reset),
    .io_out(regs_372_io_out),
    .io_enable(regs_372_io_enable)
  );
  FringeFF regs_373 ( // @[RegFile.scala 66:20:@39478.4]
    .clock(regs_373_clock),
    .reset(regs_373_reset),
    .io_in(regs_373_io_in),
    .io_reset(regs_373_io_reset),
    .io_out(regs_373_io_out),
    .io_enable(regs_373_io_enable)
  );
  FringeFF regs_374 ( // @[RegFile.scala 66:20:@39492.4]
    .clock(regs_374_clock),
    .reset(regs_374_reset),
    .io_in(regs_374_io_in),
    .io_reset(regs_374_io_reset),
    .io_out(regs_374_io_out),
    .io_enable(regs_374_io_enable)
  );
  FringeFF regs_375 ( // @[RegFile.scala 66:20:@39506.4]
    .clock(regs_375_clock),
    .reset(regs_375_reset),
    .io_in(regs_375_io_in),
    .io_reset(regs_375_io_reset),
    .io_out(regs_375_io_out),
    .io_enable(regs_375_io_enable)
  );
  FringeFF regs_376 ( // @[RegFile.scala 66:20:@39520.4]
    .clock(regs_376_clock),
    .reset(regs_376_reset),
    .io_in(regs_376_io_in),
    .io_reset(regs_376_io_reset),
    .io_out(regs_376_io_out),
    .io_enable(regs_376_io_enable)
  );
  FringeFF regs_377 ( // @[RegFile.scala 66:20:@39534.4]
    .clock(regs_377_clock),
    .reset(regs_377_reset),
    .io_in(regs_377_io_in),
    .io_reset(regs_377_io_reset),
    .io_out(regs_377_io_out),
    .io_enable(regs_377_io_enable)
  );
  FringeFF regs_378 ( // @[RegFile.scala 66:20:@39548.4]
    .clock(regs_378_clock),
    .reset(regs_378_reset),
    .io_in(regs_378_io_in),
    .io_reset(regs_378_io_reset),
    .io_out(regs_378_io_out),
    .io_enable(regs_378_io_enable)
  );
  FringeFF regs_379 ( // @[RegFile.scala 66:20:@39562.4]
    .clock(regs_379_clock),
    .reset(regs_379_reset),
    .io_in(regs_379_io_in),
    .io_reset(regs_379_io_reset),
    .io_out(regs_379_io_out),
    .io_enable(regs_379_io_enable)
  );
  FringeFF regs_380 ( // @[RegFile.scala 66:20:@39576.4]
    .clock(regs_380_clock),
    .reset(regs_380_reset),
    .io_in(regs_380_io_in),
    .io_reset(regs_380_io_reset),
    .io_out(regs_380_io_out),
    .io_enable(regs_380_io_enable)
  );
  FringeFF regs_381 ( // @[RegFile.scala 66:20:@39590.4]
    .clock(regs_381_clock),
    .reset(regs_381_reset),
    .io_in(regs_381_io_in),
    .io_reset(regs_381_io_reset),
    .io_out(regs_381_io_out),
    .io_enable(regs_381_io_enable)
  );
  FringeFF regs_382 ( // @[RegFile.scala 66:20:@39604.4]
    .clock(regs_382_clock),
    .reset(regs_382_reset),
    .io_in(regs_382_io_in),
    .io_reset(regs_382_io_reset),
    .io_out(regs_382_io_out),
    .io_enable(regs_382_io_enable)
  );
  FringeFF regs_383 ( // @[RegFile.scala 66:20:@39618.4]
    .clock(regs_383_clock),
    .reset(regs_383_reset),
    .io_in(regs_383_io_in),
    .io_reset(regs_383_io_reset),
    .io_out(regs_383_io_out),
    .io_enable(regs_383_io_enable)
  );
  FringeFF regs_384 ( // @[RegFile.scala 66:20:@39632.4]
    .clock(regs_384_clock),
    .reset(regs_384_reset),
    .io_in(regs_384_io_in),
    .io_reset(regs_384_io_reset),
    .io_out(regs_384_io_out),
    .io_enable(regs_384_io_enable)
  );
  FringeFF regs_385 ( // @[RegFile.scala 66:20:@39646.4]
    .clock(regs_385_clock),
    .reset(regs_385_reset),
    .io_in(regs_385_io_in),
    .io_reset(regs_385_io_reset),
    .io_out(regs_385_io_out),
    .io_enable(regs_385_io_enable)
  );
  FringeFF regs_386 ( // @[RegFile.scala 66:20:@39660.4]
    .clock(regs_386_clock),
    .reset(regs_386_reset),
    .io_in(regs_386_io_in),
    .io_reset(regs_386_io_reset),
    .io_out(regs_386_io_out),
    .io_enable(regs_386_io_enable)
  );
  FringeFF regs_387 ( // @[RegFile.scala 66:20:@39674.4]
    .clock(regs_387_clock),
    .reset(regs_387_reset),
    .io_in(regs_387_io_in),
    .io_reset(regs_387_io_reset),
    .io_out(regs_387_io_out),
    .io_enable(regs_387_io_enable)
  );
  FringeFF regs_388 ( // @[RegFile.scala 66:20:@39688.4]
    .clock(regs_388_clock),
    .reset(regs_388_reset),
    .io_in(regs_388_io_in),
    .io_reset(regs_388_io_reset),
    .io_out(regs_388_io_out),
    .io_enable(regs_388_io_enable)
  );
  FringeFF regs_389 ( // @[RegFile.scala 66:20:@39702.4]
    .clock(regs_389_clock),
    .reset(regs_389_reset),
    .io_in(regs_389_io_in),
    .io_reset(regs_389_io_reset),
    .io_out(regs_389_io_out),
    .io_enable(regs_389_io_enable)
  );
  FringeFF regs_390 ( // @[RegFile.scala 66:20:@39716.4]
    .clock(regs_390_clock),
    .reset(regs_390_reset),
    .io_in(regs_390_io_in),
    .io_reset(regs_390_io_reset),
    .io_out(regs_390_io_out),
    .io_enable(regs_390_io_enable)
  );
  FringeFF regs_391 ( // @[RegFile.scala 66:20:@39730.4]
    .clock(regs_391_clock),
    .reset(regs_391_reset),
    .io_in(regs_391_io_in),
    .io_reset(regs_391_io_reset),
    .io_out(regs_391_io_out),
    .io_enable(regs_391_io_enable)
  );
  FringeFF regs_392 ( // @[RegFile.scala 66:20:@39744.4]
    .clock(regs_392_clock),
    .reset(regs_392_reset),
    .io_in(regs_392_io_in),
    .io_reset(regs_392_io_reset),
    .io_out(regs_392_io_out),
    .io_enable(regs_392_io_enable)
  );
  FringeFF regs_393 ( // @[RegFile.scala 66:20:@39758.4]
    .clock(regs_393_clock),
    .reset(regs_393_reset),
    .io_in(regs_393_io_in),
    .io_reset(regs_393_io_reset),
    .io_out(regs_393_io_out),
    .io_enable(regs_393_io_enable)
  );
  FringeFF regs_394 ( // @[RegFile.scala 66:20:@39772.4]
    .clock(regs_394_clock),
    .reset(regs_394_reset),
    .io_in(regs_394_io_in),
    .io_reset(regs_394_io_reset),
    .io_out(regs_394_io_out),
    .io_enable(regs_394_io_enable)
  );
  FringeFF regs_395 ( // @[RegFile.scala 66:20:@39786.4]
    .clock(regs_395_clock),
    .reset(regs_395_reset),
    .io_in(regs_395_io_in),
    .io_reset(regs_395_io_reset),
    .io_out(regs_395_io_out),
    .io_enable(regs_395_io_enable)
  );
  FringeFF regs_396 ( // @[RegFile.scala 66:20:@39800.4]
    .clock(regs_396_clock),
    .reset(regs_396_reset),
    .io_in(regs_396_io_in),
    .io_reset(regs_396_io_reset),
    .io_out(regs_396_io_out),
    .io_enable(regs_396_io_enable)
  );
  FringeFF regs_397 ( // @[RegFile.scala 66:20:@39814.4]
    .clock(regs_397_clock),
    .reset(regs_397_reset),
    .io_in(regs_397_io_in),
    .io_reset(regs_397_io_reset),
    .io_out(regs_397_io_out),
    .io_enable(regs_397_io_enable)
  );
  FringeFF regs_398 ( // @[RegFile.scala 66:20:@39828.4]
    .clock(regs_398_clock),
    .reset(regs_398_reset),
    .io_in(regs_398_io_in),
    .io_reset(regs_398_io_reset),
    .io_out(regs_398_io_out),
    .io_enable(regs_398_io_enable)
  );
  FringeFF regs_399 ( // @[RegFile.scala 66:20:@39842.4]
    .clock(regs_399_clock),
    .reset(regs_399_reset),
    .io_in(regs_399_io_in),
    .io_reset(regs_399_io_reset),
    .io_out(regs_399_io_out),
    .io_enable(regs_399_io_enable)
  );
  FringeFF regs_400 ( // @[RegFile.scala 66:20:@39856.4]
    .clock(regs_400_clock),
    .reset(regs_400_reset),
    .io_in(regs_400_io_in),
    .io_reset(regs_400_io_reset),
    .io_out(regs_400_io_out),
    .io_enable(regs_400_io_enable)
  );
  FringeFF regs_401 ( // @[RegFile.scala 66:20:@39870.4]
    .clock(regs_401_clock),
    .reset(regs_401_reset),
    .io_in(regs_401_io_in),
    .io_reset(regs_401_io_reset),
    .io_out(regs_401_io_out),
    .io_enable(regs_401_io_enable)
  );
  FringeFF regs_402 ( // @[RegFile.scala 66:20:@39884.4]
    .clock(regs_402_clock),
    .reset(regs_402_reset),
    .io_in(regs_402_io_in),
    .io_reset(regs_402_io_reset),
    .io_out(regs_402_io_out),
    .io_enable(regs_402_io_enable)
  );
  FringeFF regs_403 ( // @[RegFile.scala 66:20:@39898.4]
    .clock(regs_403_clock),
    .reset(regs_403_reset),
    .io_in(regs_403_io_in),
    .io_reset(regs_403_io_reset),
    .io_out(regs_403_io_out),
    .io_enable(regs_403_io_enable)
  );
  FringeFF regs_404 ( // @[RegFile.scala 66:20:@39912.4]
    .clock(regs_404_clock),
    .reset(regs_404_reset),
    .io_in(regs_404_io_in),
    .io_reset(regs_404_io_reset),
    .io_out(regs_404_io_out),
    .io_enable(regs_404_io_enable)
  );
  FringeFF regs_405 ( // @[RegFile.scala 66:20:@39926.4]
    .clock(regs_405_clock),
    .reset(regs_405_reset),
    .io_in(regs_405_io_in),
    .io_reset(regs_405_io_reset),
    .io_out(regs_405_io_out),
    .io_enable(regs_405_io_enable)
  );
  FringeFF regs_406 ( // @[RegFile.scala 66:20:@39940.4]
    .clock(regs_406_clock),
    .reset(regs_406_reset),
    .io_in(regs_406_io_in),
    .io_reset(regs_406_io_reset),
    .io_out(regs_406_io_out),
    .io_enable(regs_406_io_enable)
  );
  FringeFF regs_407 ( // @[RegFile.scala 66:20:@39954.4]
    .clock(regs_407_clock),
    .reset(regs_407_reset),
    .io_in(regs_407_io_in),
    .io_reset(regs_407_io_reset),
    .io_out(regs_407_io_out),
    .io_enable(regs_407_io_enable)
  );
  FringeFF regs_408 ( // @[RegFile.scala 66:20:@39968.4]
    .clock(regs_408_clock),
    .reset(regs_408_reset),
    .io_in(regs_408_io_in),
    .io_reset(regs_408_io_reset),
    .io_out(regs_408_io_out),
    .io_enable(regs_408_io_enable)
  );
  FringeFF regs_409 ( // @[RegFile.scala 66:20:@39982.4]
    .clock(regs_409_clock),
    .reset(regs_409_reset),
    .io_in(regs_409_io_in),
    .io_reset(regs_409_io_reset),
    .io_out(regs_409_io_out),
    .io_enable(regs_409_io_enable)
  );
  FringeFF regs_410 ( // @[RegFile.scala 66:20:@39996.4]
    .clock(regs_410_clock),
    .reset(regs_410_reset),
    .io_in(regs_410_io_in),
    .io_reset(regs_410_io_reset),
    .io_out(regs_410_io_out),
    .io_enable(regs_410_io_enable)
  );
  FringeFF regs_411 ( // @[RegFile.scala 66:20:@40010.4]
    .clock(regs_411_clock),
    .reset(regs_411_reset),
    .io_in(regs_411_io_in),
    .io_reset(regs_411_io_reset),
    .io_out(regs_411_io_out),
    .io_enable(regs_411_io_enable)
  );
  FringeFF regs_412 ( // @[RegFile.scala 66:20:@40024.4]
    .clock(regs_412_clock),
    .reset(regs_412_reset),
    .io_in(regs_412_io_in),
    .io_reset(regs_412_io_reset),
    .io_out(regs_412_io_out),
    .io_enable(regs_412_io_enable)
  );
  FringeFF regs_413 ( // @[RegFile.scala 66:20:@40038.4]
    .clock(regs_413_clock),
    .reset(regs_413_reset),
    .io_in(regs_413_io_in),
    .io_reset(regs_413_io_reset),
    .io_out(regs_413_io_out),
    .io_enable(regs_413_io_enable)
  );
  FringeFF regs_414 ( // @[RegFile.scala 66:20:@40052.4]
    .clock(regs_414_clock),
    .reset(regs_414_reset),
    .io_in(regs_414_io_in),
    .io_reset(regs_414_io_reset),
    .io_out(regs_414_io_out),
    .io_enable(regs_414_io_enable)
  );
  FringeFF regs_415 ( // @[RegFile.scala 66:20:@40066.4]
    .clock(regs_415_clock),
    .reset(regs_415_reset),
    .io_in(regs_415_io_in),
    .io_reset(regs_415_io_reset),
    .io_out(regs_415_io_out),
    .io_enable(regs_415_io_enable)
  );
  FringeFF regs_416 ( // @[RegFile.scala 66:20:@40080.4]
    .clock(regs_416_clock),
    .reset(regs_416_reset),
    .io_in(regs_416_io_in),
    .io_reset(regs_416_io_reset),
    .io_out(regs_416_io_out),
    .io_enable(regs_416_io_enable)
  );
  FringeFF regs_417 ( // @[RegFile.scala 66:20:@40094.4]
    .clock(regs_417_clock),
    .reset(regs_417_reset),
    .io_in(regs_417_io_in),
    .io_reset(regs_417_io_reset),
    .io_out(regs_417_io_out),
    .io_enable(regs_417_io_enable)
  );
  FringeFF regs_418 ( // @[RegFile.scala 66:20:@40108.4]
    .clock(regs_418_clock),
    .reset(regs_418_reset),
    .io_in(regs_418_io_in),
    .io_reset(regs_418_io_reset),
    .io_out(regs_418_io_out),
    .io_enable(regs_418_io_enable)
  );
  FringeFF regs_419 ( // @[RegFile.scala 66:20:@40122.4]
    .clock(regs_419_clock),
    .reset(regs_419_reset),
    .io_in(regs_419_io_in),
    .io_reset(regs_419_io_reset),
    .io_out(regs_419_io_out),
    .io_enable(regs_419_io_enable)
  );
  FringeFF regs_420 ( // @[RegFile.scala 66:20:@40136.4]
    .clock(regs_420_clock),
    .reset(regs_420_reset),
    .io_in(regs_420_io_in),
    .io_reset(regs_420_io_reset),
    .io_out(regs_420_io_out),
    .io_enable(regs_420_io_enable)
  );
  FringeFF regs_421 ( // @[RegFile.scala 66:20:@40150.4]
    .clock(regs_421_clock),
    .reset(regs_421_reset),
    .io_in(regs_421_io_in),
    .io_reset(regs_421_io_reset),
    .io_out(regs_421_io_out),
    .io_enable(regs_421_io_enable)
  );
  FringeFF regs_422 ( // @[RegFile.scala 66:20:@40164.4]
    .clock(regs_422_clock),
    .reset(regs_422_reset),
    .io_in(regs_422_io_in),
    .io_reset(regs_422_io_reset),
    .io_out(regs_422_io_out),
    .io_enable(regs_422_io_enable)
  );
  FringeFF regs_423 ( // @[RegFile.scala 66:20:@40178.4]
    .clock(regs_423_clock),
    .reset(regs_423_reset),
    .io_in(regs_423_io_in),
    .io_reset(regs_423_io_reset),
    .io_out(regs_423_io_out),
    .io_enable(regs_423_io_enable)
  );
  FringeFF regs_424 ( // @[RegFile.scala 66:20:@40192.4]
    .clock(regs_424_clock),
    .reset(regs_424_reset),
    .io_in(regs_424_io_in),
    .io_reset(regs_424_io_reset),
    .io_out(regs_424_io_out),
    .io_enable(regs_424_io_enable)
  );
  FringeFF regs_425 ( // @[RegFile.scala 66:20:@40206.4]
    .clock(regs_425_clock),
    .reset(regs_425_reset),
    .io_in(regs_425_io_in),
    .io_reset(regs_425_io_reset),
    .io_out(regs_425_io_out),
    .io_enable(regs_425_io_enable)
  );
  FringeFF regs_426 ( // @[RegFile.scala 66:20:@40220.4]
    .clock(regs_426_clock),
    .reset(regs_426_reset),
    .io_in(regs_426_io_in),
    .io_reset(regs_426_io_reset),
    .io_out(regs_426_io_out),
    .io_enable(regs_426_io_enable)
  );
  FringeFF regs_427 ( // @[RegFile.scala 66:20:@40234.4]
    .clock(regs_427_clock),
    .reset(regs_427_reset),
    .io_in(regs_427_io_in),
    .io_reset(regs_427_io_reset),
    .io_out(regs_427_io_out),
    .io_enable(regs_427_io_enable)
  );
  FringeFF regs_428 ( // @[RegFile.scala 66:20:@40248.4]
    .clock(regs_428_clock),
    .reset(regs_428_reset),
    .io_in(regs_428_io_in),
    .io_reset(regs_428_io_reset),
    .io_out(regs_428_io_out),
    .io_enable(regs_428_io_enable)
  );
  FringeFF regs_429 ( // @[RegFile.scala 66:20:@40262.4]
    .clock(regs_429_clock),
    .reset(regs_429_reset),
    .io_in(regs_429_io_in),
    .io_reset(regs_429_io_reset),
    .io_out(regs_429_io_out),
    .io_enable(regs_429_io_enable)
  );
  FringeFF regs_430 ( // @[RegFile.scala 66:20:@40276.4]
    .clock(regs_430_clock),
    .reset(regs_430_reset),
    .io_in(regs_430_io_in),
    .io_reset(regs_430_io_reset),
    .io_out(regs_430_io_out),
    .io_enable(regs_430_io_enable)
  );
  FringeFF regs_431 ( // @[RegFile.scala 66:20:@40290.4]
    .clock(regs_431_clock),
    .reset(regs_431_reset),
    .io_in(regs_431_io_in),
    .io_reset(regs_431_io_reset),
    .io_out(regs_431_io_out),
    .io_enable(regs_431_io_enable)
  );
  FringeFF regs_432 ( // @[RegFile.scala 66:20:@40304.4]
    .clock(regs_432_clock),
    .reset(regs_432_reset),
    .io_in(regs_432_io_in),
    .io_reset(regs_432_io_reset),
    .io_out(regs_432_io_out),
    .io_enable(regs_432_io_enable)
  );
  FringeFF regs_433 ( // @[RegFile.scala 66:20:@40318.4]
    .clock(regs_433_clock),
    .reset(regs_433_reset),
    .io_in(regs_433_io_in),
    .io_reset(regs_433_io_reset),
    .io_out(regs_433_io_out),
    .io_enable(regs_433_io_enable)
  );
  FringeFF regs_434 ( // @[RegFile.scala 66:20:@40332.4]
    .clock(regs_434_clock),
    .reset(regs_434_reset),
    .io_in(regs_434_io_in),
    .io_reset(regs_434_io_reset),
    .io_out(regs_434_io_out),
    .io_enable(regs_434_io_enable)
  );
  FringeFF regs_435 ( // @[RegFile.scala 66:20:@40346.4]
    .clock(regs_435_clock),
    .reset(regs_435_reset),
    .io_in(regs_435_io_in),
    .io_reset(regs_435_io_reset),
    .io_out(regs_435_io_out),
    .io_enable(regs_435_io_enable)
  );
  FringeFF regs_436 ( // @[RegFile.scala 66:20:@40360.4]
    .clock(regs_436_clock),
    .reset(regs_436_reset),
    .io_in(regs_436_io_in),
    .io_reset(regs_436_io_reset),
    .io_out(regs_436_io_out),
    .io_enable(regs_436_io_enable)
  );
  FringeFF regs_437 ( // @[RegFile.scala 66:20:@40374.4]
    .clock(regs_437_clock),
    .reset(regs_437_reset),
    .io_in(regs_437_io_in),
    .io_reset(regs_437_io_reset),
    .io_out(regs_437_io_out),
    .io_enable(regs_437_io_enable)
  );
  FringeFF regs_438 ( // @[RegFile.scala 66:20:@40388.4]
    .clock(regs_438_clock),
    .reset(regs_438_reset),
    .io_in(regs_438_io_in),
    .io_reset(regs_438_io_reset),
    .io_out(regs_438_io_out),
    .io_enable(regs_438_io_enable)
  );
  FringeFF regs_439 ( // @[RegFile.scala 66:20:@40402.4]
    .clock(regs_439_clock),
    .reset(regs_439_reset),
    .io_in(regs_439_io_in),
    .io_reset(regs_439_io_reset),
    .io_out(regs_439_io_out),
    .io_enable(regs_439_io_enable)
  );
  FringeFF regs_440 ( // @[RegFile.scala 66:20:@40416.4]
    .clock(regs_440_clock),
    .reset(regs_440_reset),
    .io_in(regs_440_io_in),
    .io_reset(regs_440_io_reset),
    .io_out(regs_440_io_out),
    .io_enable(regs_440_io_enable)
  );
  FringeFF regs_441 ( // @[RegFile.scala 66:20:@40430.4]
    .clock(regs_441_clock),
    .reset(regs_441_reset),
    .io_in(regs_441_io_in),
    .io_reset(regs_441_io_reset),
    .io_out(regs_441_io_out),
    .io_enable(regs_441_io_enable)
  );
  FringeFF regs_442 ( // @[RegFile.scala 66:20:@40444.4]
    .clock(regs_442_clock),
    .reset(regs_442_reset),
    .io_in(regs_442_io_in),
    .io_reset(regs_442_io_reset),
    .io_out(regs_442_io_out),
    .io_enable(regs_442_io_enable)
  );
  FringeFF regs_443 ( // @[RegFile.scala 66:20:@40458.4]
    .clock(regs_443_clock),
    .reset(regs_443_reset),
    .io_in(regs_443_io_in),
    .io_reset(regs_443_io_reset),
    .io_out(regs_443_io_out),
    .io_enable(regs_443_io_enable)
  );
  FringeFF regs_444 ( // @[RegFile.scala 66:20:@40472.4]
    .clock(regs_444_clock),
    .reset(regs_444_reset),
    .io_in(regs_444_io_in),
    .io_reset(regs_444_io_reset),
    .io_out(regs_444_io_out),
    .io_enable(regs_444_io_enable)
  );
  FringeFF regs_445 ( // @[RegFile.scala 66:20:@40486.4]
    .clock(regs_445_clock),
    .reset(regs_445_reset),
    .io_in(regs_445_io_in),
    .io_reset(regs_445_io_reset),
    .io_out(regs_445_io_out),
    .io_enable(regs_445_io_enable)
  );
  FringeFF regs_446 ( // @[RegFile.scala 66:20:@40500.4]
    .clock(regs_446_clock),
    .reset(regs_446_reset),
    .io_in(regs_446_io_in),
    .io_reset(regs_446_io_reset),
    .io_out(regs_446_io_out),
    .io_enable(regs_446_io_enable)
  );
  FringeFF regs_447 ( // @[RegFile.scala 66:20:@40514.4]
    .clock(regs_447_clock),
    .reset(regs_447_reset),
    .io_in(regs_447_io_in),
    .io_reset(regs_447_io_reset),
    .io_out(regs_447_io_out),
    .io_enable(regs_447_io_enable)
  );
  FringeFF regs_448 ( // @[RegFile.scala 66:20:@40528.4]
    .clock(regs_448_clock),
    .reset(regs_448_reset),
    .io_in(regs_448_io_in),
    .io_reset(regs_448_io_reset),
    .io_out(regs_448_io_out),
    .io_enable(regs_448_io_enable)
  );
  FringeFF regs_449 ( // @[RegFile.scala 66:20:@40542.4]
    .clock(regs_449_clock),
    .reset(regs_449_reset),
    .io_in(regs_449_io_in),
    .io_reset(regs_449_io_reset),
    .io_out(regs_449_io_out),
    .io_enable(regs_449_io_enable)
  );
  FringeFF regs_450 ( // @[RegFile.scala 66:20:@40556.4]
    .clock(regs_450_clock),
    .reset(regs_450_reset),
    .io_in(regs_450_io_in),
    .io_reset(regs_450_io_reset),
    .io_out(regs_450_io_out),
    .io_enable(regs_450_io_enable)
  );
  FringeFF regs_451 ( // @[RegFile.scala 66:20:@40570.4]
    .clock(regs_451_clock),
    .reset(regs_451_reset),
    .io_in(regs_451_io_in),
    .io_reset(regs_451_io_reset),
    .io_out(regs_451_io_out),
    .io_enable(regs_451_io_enable)
  );
  FringeFF regs_452 ( // @[RegFile.scala 66:20:@40584.4]
    .clock(regs_452_clock),
    .reset(regs_452_reset),
    .io_in(regs_452_io_in),
    .io_reset(regs_452_io_reset),
    .io_out(regs_452_io_out),
    .io_enable(regs_452_io_enable)
  );
  FringeFF regs_453 ( // @[RegFile.scala 66:20:@40598.4]
    .clock(regs_453_clock),
    .reset(regs_453_reset),
    .io_in(regs_453_io_in),
    .io_reset(regs_453_io_reset),
    .io_out(regs_453_io_out),
    .io_enable(regs_453_io_enable)
  );
  FringeFF regs_454 ( // @[RegFile.scala 66:20:@40612.4]
    .clock(regs_454_clock),
    .reset(regs_454_reset),
    .io_in(regs_454_io_in),
    .io_reset(regs_454_io_reset),
    .io_out(regs_454_io_out),
    .io_enable(regs_454_io_enable)
  );
  FringeFF regs_455 ( // @[RegFile.scala 66:20:@40626.4]
    .clock(regs_455_clock),
    .reset(regs_455_reset),
    .io_in(regs_455_io_in),
    .io_reset(regs_455_io_reset),
    .io_out(regs_455_io_out),
    .io_enable(regs_455_io_enable)
  );
  FringeFF regs_456 ( // @[RegFile.scala 66:20:@40640.4]
    .clock(regs_456_clock),
    .reset(regs_456_reset),
    .io_in(regs_456_io_in),
    .io_reset(regs_456_io_reset),
    .io_out(regs_456_io_out),
    .io_enable(regs_456_io_enable)
  );
  FringeFF regs_457 ( // @[RegFile.scala 66:20:@40654.4]
    .clock(regs_457_clock),
    .reset(regs_457_reset),
    .io_in(regs_457_io_in),
    .io_reset(regs_457_io_reset),
    .io_out(regs_457_io_out),
    .io_enable(regs_457_io_enable)
  );
  FringeFF regs_458 ( // @[RegFile.scala 66:20:@40668.4]
    .clock(regs_458_clock),
    .reset(regs_458_reset),
    .io_in(regs_458_io_in),
    .io_reset(regs_458_io_reset),
    .io_out(regs_458_io_out),
    .io_enable(regs_458_io_enable)
  );
  FringeFF regs_459 ( // @[RegFile.scala 66:20:@40682.4]
    .clock(regs_459_clock),
    .reset(regs_459_reset),
    .io_in(regs_459_io_in),
    .io_reset(regs_459_io_reset),
    .io_out(regs_459_io_out),
    .io_enable(regs_459_io_enable)
  );
  FringeFF regs_460 ( // @[RegFile.scala 66:20:@40696.4]
    .clock(regs_460_clock),
    .reset(regs_460_reset),
    .io_in(regs_460_io_in),
    .io_reset(regs_460_io_reset),
    .io_out(regs_460_io_out),
    .io_enable(regs_460_io_enable)
  );
  FringeFF regs_461 ( // @[RegFile.scala 66:20:@40710.4]
    .clock(regs_461_clock),
    .reset(regs_461_reset),
    .io_in(regs_461_io_in),
    .io_reset(regs_461_io_reset),
    .io_out(regs_461_io_out),
    .io_enable(regs_461_io_enable)
  );
  FringeFF regs_462 ( // @[RegFile.scala 66:20:@40724.4]
    .clock(regs_462_clock),
    .reset(regs_462_reset),
    .io_in(regs_462_io_in),
    .io_reset(regs_462_io_reset),
    .io_out(regs_462_io_out),
    .io_enable(regs_462_io_enable)
  );
  FringeFF regs_463 ( // @[RegFile.scala 66:20:@40738.4]
    .clock(regs_463_clock),
    .reset(regs_463_reset),
    .io_in(regs_463_io_in),
    .io_reset(regs_463_io_reset),
    .io_out(regs_463_io_out),
    .io_enable(regs_463_io_enable)
  );
  FringeFF regs_464 ( // @[RegFile.scala 66:20:@40752.4]
    .clock(regs_464_clock),
    .reset(regs_464_reset),
    .io_in(regs_464_io_in),
    .io_reset(regs_464_io_reset),
    .io_out(regs_464_io_out),
    .io_enable(regs_464_io_enable)
  );
  FringeFF regs_465 ( // @[RegFile.scala 66:20:@40766.4]
    .clock(regs_465_clock),
    .reset(regs_465_reset),
    .io_in(regs_465_io_in),
    .io_reset(regs_465_io_reset),
    .io_out(regs_465_io_out),
    .io_enable(regs_465_io_enable)
  );
  FringeFF regs_466 ( // @[RegFile.scala 66:20:@40780.4]
    .clock(regs_466_clock),
    .reset(regs_466_reset),
    .io_in(regs_466_io_in),
    .io_reset(regs_466_io_reset),
    .io_out(regs_466_io_out),
    .io_enable(regs_466_io_enable)
  );
  FringeFF regs_467 ( // @[RegFile.scala 66:20:@40794.4]
    .clock(regs_467_clock),
    .reset(regs_467_reset),
    .io_in(regs_467_io_in),
    .io_reset(regs_467_io_reset),
    .io_out(regs_467_io_out),
    .io_enable(regs_467_io_enable)
  );
  FringeFF regs_468 ( // @[RegFile.scala 66:20:@40808.4]
    .clock(regs_468_clock),
    .reset(regs_468_reset),
    .io_in(regs_468_io_in),
    .io_reset(regs_468_io_reset),
    .io_out(regs_468_io_out),
    .io_enable(regs_468_io_enable)
  );
  FringeFF regs_469 ( // @[RegFile.scala 66:20:@40822.4]
    .clock(regs_469_clock),
    .reset(regs_469_reset),
    .io_in(regs_469_io_in),
    .io_reset(regs_469_io_reset),
    .io_out(regs_469_io_out),
    .io_enable(regs_469_io_enable)
  );
  FringeFF regs_470 ( // @[RegFile.scala 66:20:@40836.4]
    .clock(regs_470_clock),
    .reset(regs_470_reset),
    .io_in(regs_470_io_in),
    .io_reset(regs_470_io_reset),
    .io_out(regs_470_io_out),
    .io_enable(regs_470_io_enable)
  );
  FringeFF regs_471 ( // @[RegFile.scala 66:20:@40850.4]
    .clock(regs_471_clock),
    .reset(regs_471_reset),
    .io_in(regs_471_io_in),
    .io_reset(regs_471_io_reset),
    .io_out(regs_471_io_out),
    .io_enable(regs_471_io_enable)
  );
  FringeFF regs_472 ( // @[RegFile.scala 66:20:@40864.4]
    .clock(regs_472_clock),
    .reset(regs_472_reset),
    .io_in(regs_472_io_in),
    .io_reset(regs_472_io_reset),
    .io_out(regs_472_io_out),
    .io_enable(regs_472_io_enable)
  );
  FringeFF regs_473 ( // @[RegFile.scala 66:20:@40878.4]
    .clock(regs_473_clock),
    .reset(regs_473_reset),
    .io_in(regs_473_io_in),
    .io_reset(regs_473_io_reset),
    .io_out(regs_473_io_out),
    .io_enable(regs_473_io_enable)
  );
  FringeFF regs_474 ( // @[RegFile.scala 66:20:@40892.4]
    .clock(regs_474_clock),
    .reset(regs_474_reset),
    .io_in(regs_474_io_in),
    .io_reset(regs_474_io_reset),
    .io_out(regs_474_io_out),
    .io_enable(regs_474_io_enable)
  );
  FringeFF regs_475 ( // @[RegFile.scala 66:20:@40906.4]
    .clock(regs_475_clock),
    .reset(regs_475_reset),
    .io_in(regs_475_io_in),
    .io_reset(regs_475_io_reset),
    .io_out(regs_475_io_out),
    .io_enable(regs_475_io_enable)
  );
  FringeFF regs_476 ( // @[RegFile.scala 66:20:@40920.4]
    .clock(regs_476_clock),
    .reset(regs_476_reset),
    .io_in(regs_476_io_in),
    .io_reset(regs_476_io_reset),
    .io_out(regs_476_io_out),
    .io_enable(regs_476_io_enable)
  );
  FringeFF regs_477 ( // @[RegFile.scala 66:20:@40934.4]
    .clock(regs_477_clock),
    .reset(regs_477_reset),
    .io_in(regs_477_io_in),
    .io_reset(regs_477_io_reset),
    .io_out(regs_477_io_out),
    .io_enable(regs_477_io_enable)
  );
  FringeFF regs_478 ( // @[RegFile.scala 66:20:@40948.4]
    .clock(regs_478_clock),
    .reset(regs_478_reset),
    .io_in(regs_478_io_in),
    .io_reset(regs_478_io_reset),
    .io_out(regs_478_io_out),
    .io_enable(regs_478_io_enable)
  );
  FringeFF regs_479 ( // @[RegFile.scala 66:20:@40962.4]
    .clock(regs_479_clock),
    .reset(regs_479_reset),
    .io_in(regs_479_io_in),
    .io_reset(regs_479_io_reset),
    .io_out(regs_479_io_out),
    .io_enable(regs_479_io_enable)
  );
  FringeFF regs_480 ( // @[RegFile.scala 66:20:@40976.4]
    .clock(regs_480_clock),
    .reset(regs_480_reset),
    .io_in(regs_480_io_in),
    .io_reset(regs_480_io_reset),
    .io_out(regs_480_io_out),
    .io_enable(regs_480_io_enable)
  );
  FringeFF regs_481 ( // @[RegFile.scala 66:20:@40990.4]
    .clock(regs_481_clock),
    .reset(regs_481_reset),
    .io_in(regs_481_io_in),
    .io_reset(regs_481_io_reset),
    .io_out(regs_481_io_out),
    .io_enable(regs_481_io_enable)
  );
  FringeFF regs_482 ( // @[RegFile.scala 66:20:@41004.4]
    .clock(regs_482_clock),
    .reset(regs_482_reset),
    .io_in(regs_482_io_in),
    .io_reset(regs_482_io_reset),
    .io_out(regs_482_io_out),
    .io_enable(regs_482_io_enable)
  );
  FringeFF regs_483 ( // @[RegFile.scala 66:20:@41018.4]
    .clock(regs_483_clock),
    .reset(regs_483_reset),
    .io_in(regs_483_io_in),
    .io_reset(regs_483_io_reset),
    .io_out(regs_483_io_out),
    .io_enable(regs_483_io_enable)
  );
  FringeFF regs_484 ( // @[RegFile.scala 66:20:@41032.4]
    .clock(regs_484_clock),
    .reset(regs_484_reset),
    .io_in(regs_484_io_in),
    .io_reset(regs_484_io_reset),
    .io_out(regs_484_io_out),
    .io_enable(regs_484_io_enable)
  );
  FringeFF regs_485 ( // @[RegFile.scala 66:20:@41046.4]
    .clock(regs_485_clock),
    .reset(regs_485_reset),
    .io_in(regs_485_io_in),
    .io_reset(regs_485_io_reset),
    .io_out(regs_485_io_out),
    .io_enable(regs_485_io_enable)
  );
  FringeFF regs_486 ( // @[RegFile.scala 66:20:@41060.4]
    .clock(regs_486_clock),
    .reset(regs_486_reset),
    .io_in(regs_486_io_in),
    .io_reset(regs_486_io_reset),
    .io_out(regs_486_io_out),
    .io_enable(regs_486_io_enable)
  );
  FringeFF regs_487 ( // @[RegFile.scala 66:20:@41074.4]
    .clock(regs_487_clock),
    .reset(regs_487_reset),
    .io_in(regs_487_io_in),
    .io_reset(regs_487_io_reset),
    .io_out(regs_487_io_out),
    .io_enable(regs_487_io_enable)
  );
  FringeFF regs_488 ( // @[RegFile.scala 66:20:@41088.4]
    .clock(regs_488_clock),
    .reset(regs_488_reset),
    .io_in(regs_488_io_in),
    .io_reset(regs_488_io_reset),
    .io_out(regs_488_io_out),
    .io_enable(regs_488_io_enable)
  );
  FringeFF regs_489 ( // @[RegFile.scala 66:20:@41102.4]
    .clock(regs_489_clock),
    .reset(regs_489_reset),
    .io_in(regs_489_io_in),
    .io_reset(regs_489_io_reset),
    .io_out(regs_489_io_out),
    .io_enable(regs_489_io_enable)
  );
  FringeFF regs_490 ( // @[RegFile.scala 66:20:@41116.4]
    .clock(regs_490_clock),
    .reset(regs_490_reset),
    .io_in(regs_490_io_in),
    .io_reset(regs_490_io_reset),
    .io_out(regs_490_io_out),
    .io_enable(regs_490_io_enable)
  );
  FringeFF regs_491 ( // @[RegFile.scala 66:20:@41130.4]
    .clock(regs_491_clock),
    .reset(regs_491_reset),
    .io_in(regs_491_io_in),
    .io_reset(regs_491_io_reset),
    .io_out(regs_491_io_out),
    .io_enable(regs_491_io_enable)
  );
  FringeFF regs_492 ( // @[RegFile.scala 66:20:@41144.4]
    .clock(regs_492_clock),
    .reset(regs_492_reset),
    .io_in(regs_492_io_in),
    .io_reset(regs_492_io_reset),
    .io_out(regs_492_io_out),
    .io_enable(regs_492_io_enable)
  );
  FringeFF regs_493 ( // @[RegFile.scala 66:20:@41158.4]
    .clock(regs_493_clock),
    .reset(regs_493_reset),
    .io_in(regs_493_io_in),
    .io_reset(regs_493_io_reset),
    .io_out(regs_493_io_out),
    .io_enable(regs_493_io_enable)
  );
  FringeFF regs_494 ( // @[RegFile.scala 66:20:@41172.4]
    .clock(regs_494_clock),
    .reset(regs_494_reset),
    .io_in(regs_494_io_in),
    .io_reset(regs_494_io_reset),
    .io_out(regs_494_io_out),
    .io_enable(regs_494_io_enable)
  );
  FringeFF regs_495 ( // @[RegFile.scala 66:20:@41186.4]
    .clock(regs_495_clock),
    .reset(regs_495_reset),
    .io_in(regs_495_io_in),
    .io_reset(regs_495_io_reset),
    .io_out(regs_495_io_out),
    .io_enable(regs_495_io_enable)
  );
  FringeFF regs_496 ( // @[RegFile.scala 66:20:@41200.4]
    .clock(regs_496_clock),
    .reset(regs_496_reset),
    .io_in(regs_496_io_in),
    .io_reset(regs_496_io_reset),
    .io_out(regs_496_io_out),
    .io_enable(regs_496_io_enable)
  );
  FringeFF regs_497 ( // @[RegFile.scala 66:20:@41214.4]
    .clock(regs_497_clock),
    .reset(regs_497_reset),
    .io_in(regs_497_io_in),
    .io_reset(regs_497_io_reset),
    .io_out(regs_497_io_out),
    .io_enable(regs_497_io_enable)
  );
  FringeFF regs_498 ( // @[RegFile.scala 66:20:@41228.4]
    .clock(regs_498_clock),
    .reset(regs_498_reset),
    .io_in(regs_498_io_in),
    .io_reset(regs_498_io_reset),
    .io_out(regs_498_io_out),
    .io_enable(regs_498_io_enable)
  );
  FringeFF regs_499 ( // @[RegFile.scala 66:20:@41242.4]
    .clock(regs_499_clock),
    .reset(regs_499_reset),
    .io_in(regs_499_io_in),
    .io_reset(regs_499_io_reset),
    .io_out(regs_499_io_out),
    .io_enable(regs_499_io_enable)
  );
  FringeFF regs_500 ( // @[RegFile.scala 66:20:@41256.4]
    .clock(regs_500_clock),
    .reset(regs_500_reset),
    .io_in(regs_500_io_in),
    .io_reset(regs_500_io_reset),
    .io_out(regs_500_io_out),
    .io_enable(regs_500_io_enable)
  );
  FringeFF regs_501 ( // @[RegFile.scala 66:20:@41270.4]
    .clock(regs_501_clock),
    .reset(regs_501_reset),
    .io_in(regs_501_io_in),
    .io_reset(regs_501_io_reset),
    .io_out(regs_501_io_out),
    .io_enable(regs_501_io_enable)
  );
  FringeFF regs_502 ( // @[RegFile.scala 66:20:@41284.4]
    .clock(regs_502_clock),
    .reset(regs_502_reset),
    .io_in(regs_502_io_in),
    .io_reset(regs_502_io_reset),
    .io_out(regs_502_io_out),
    .io_enable(regs_502_io_enable)
  );
  MuxN rport ( // @[RegFile.scala 95:21:@41298.4]
    .io_ins_0(rport_io_ins_0),
    .io_ins_1(rport_io_ins_1),
    .io_ins_2(rport_io_ins_2),
    .io_ins_3(rport_io_ins_3),
    .io_ins_4(rport_io_ins_4),
    .io_ins_5(rport_io_ins_5),
    .io_ins_6(rport_io_ins_6),
    .io_ins_7(rport_io_ins_7),
    .io_ins_8(rport_io_ins_8),
    .io_ins_9(rport_io_ins_9),
    .io_ins_10(rport_io_ins_10),
    .io_ins_11(rport_io_ins_11),
    .io_ins_12(rport_io_ins_12),
    .io_ins_13(rport_io_ins_13),
    .io_ins_14(rport_io_ins_14),
    .io_ins_15(rport_io_ins_15),
    .io_ins_16(rport_io_ins_16),
    .io_ins_17(rport_io_ins_17),
    .io_ins_18(rport_io_ins_18),
    .io_ins_19(rport_io_ins_19),
    .io_ins_20(rport_io_ins_20),
    .io_ins_21(rport_io_ins_21),
    .io_ins_22(rport_io_ins_22),
    .io_ins_23(rport_io_ins_23),
    .io_ins_24(rport_io_ins_24),
    .io_ins_25(rport_io_ins_25),
    .io_ins_26(rport_io_ins_26),
    .io_ins_27(rport_io_ins_27),
    .io_ins_28(rport_io_ins_28),
    .io_ins_29(rport_io_ins_29),
    .io_ins_30(rport_io_ins_30),
    .io_ins_31(rport_io_ins_31),
    .io_ins_32(rport_io_ins_32),
    .io_ins_33(rport_io_ins_33),
    .io_ins_34(rport_io_ins_34),
    .io_ins_35(rport_io_ins_35),
    .io_ins_36(rport_io_ins_36),
    .io_ins_37(rport_io_ins_37),
    .io_ins_38(rport_io_ins_38),
    .io_ins_39(rport_io_ins_39),
    .io_ins_40(rport_io_ins_40),
    .io_ins_41(rport_io_ins_41),
    .io_ins_42(rport_io_ins_42),
    .io_ins_43(rport_io_ins_43),
    .io_ins_44(rport_io_ins_44),
    .io_ins_45(rport_io_ins_45),
    .io_ins_46(rport_io_ins_46),
    .io_ins_47(rport_io_ins_47),
    .io_ins_48(rport_io_ins_48),
    .io_ins_49(rport_io_ins_49),
    .io_ins_50(rport_io_ins_50),
    .io_ins_51(rport_io_ins_51),
    .io_ins_52(rport_io_ins_52),
    .io_ins_53(rport_io_ins_53),
    .io_ins_54(rport_io_ins_54),
    .io_ins_55(rport_io_ins_55),
    .io_ins_56(rport_io_ins_56),
    .io_ins_57(rport_io_ins_57),
    .io_ins_58(rport_io_ins_58),
    .io_ins_59(rport_io_ins_59),
    .io_ins_60(rport_io_ins_60),
    .io_ins_61(rport_io_ins_61),
    .io_ins_62(rport_io_ins_62),
    .io_ins_63(rport_io_ins_63),
    .io_ins_64(rport_io_ins_64),
    .io_ins_65(rport_io_ins_65),
    .io_ins_66(rport_io_ins_66),
    .io_ins_67(rport_io_ins_67),
    .io_ins_68(rport_io_ins_68),
    .io_ins_69(rport_io_ins_69),
    .io_ins_70(rport_io_ins_70),
    .io_ins_71(rport_io_ins_71),
    .io_ins_72(rport_io_ins_72),
    .io_ins_73(rport_io_ins_73),
    .io_ins_74(rport_io_ins_74),
    .io_ins_75(rport_io_ins_75),
    .io_ins_76(rport_io_ins_76),
    .io_ins_77(rport_io_ins_77),
    .io_ins_78(rport_io_ins_78),
    .io_ins_79(rport_io_ins_79),
    .io_ins_80(rport_io_ins_80),
    .io_ins_81(rport_io_ins_81),
    .io_ins_82(rport_io_ins_82),
    .io_ins_83(rport_io_ins_83),
    .io_ins_84(rport_io_ins_84),
    .io_ins_85(rport_io_ins_85),
    .io_ins_86(rport_io_ins_86),
    .io_ins_87(rport_io_ins_87),
    .io_ins_88(rport_io_ins_88),
    .io_ins_89(rport_io_ins_89),
    .io_ins_90(rport_io_ins_90),
    .io_ins_91(rport_io_ins_91),
    .io_ins_92(rport_io_ins_92),
    .io_ins_93(rport_io_ins_93),
    .io_ins_94(rport_io_ins_94),
    .io_ins_95(rport_io_ins_95),
    .io_ins_96(rport_io_ins_96),
    .io_ins_97(rport_io_ins_97),
    .io_ins_98(rport_io_ins_98),
    .io_ins_99(rport_io_ins_99),
    .io_ins_100(rport_io_ins_100),
    .io_ins_101(rport_io_ins_101),
    .io_ins_102(rport_io_ins_102),
    .io_ins_103(rport_io_ins_103),
    .io_ins_104(rport_io_ins_104),
    .io_ins_105(rport_io_ins_105),
    .io_ins_106(rport_io_ins_106),
    .io_ins_107(rport_io_ins_107),
    .io_ins_108(rport_io_ins_108),
    .io_ins_109(rport_io_ins_109),
    .io_ins_110(rport_io_ins_110),
    .io_ins_111(rport_io_ins_111),
    .io_ins_112(rport_io_ins_112),
    .io_ins_113(rport_io_ins_113),
    .io_ins_114(rport_io_ins_114),
    .io_ins_115(rport_io_ins_115),
    .io_ins_116(rport_io_ins_116),
    .io_ins_117(rport_io_ins_117),
    .io_ins_118(rport_io_ins_118),
    .io_ins_119(rport_io_ins_119),
    .io_ins_120(rport_io_ins_120),
    .io_ins_121(rport_io_ins_121),
    .io_ins_122(rport_io_ins_122),
    .io_ins_123(rport_io_ins_123),
    .io_ins_124(rport_io_ins_124),
    .io_ins_125(rport_io_ins_125),
    .io_ins_126(rport_io_ins_126),
    .io_ins_127(rport_io_ins_127),
    .io_ins_128(rport_io_ins_128),
    .io_ins_129(rport_io_ins_129),
    .io_ins_130(rport_io_ins_130),
    .io_ins_131(rport_io_ins_131),
    .io_ins_132(rport_io_ins_132),
    .io_ins_133(rport_io_ins_133),
    .io_ins_134(rport_io_ins_134),
    .io_ins_135(rport_io_ins_135),
    .io_ins_136(rport_io_ins_136),
    .io_ins_137(rport_io_ins_137),
    .io_ins_138(rport_io_ins_138),
    .io_ins_139(rport_io_ins_139),
    .io_ins_140(rport_io_ins_140),
    .io_ins_141(rport_io_ins_141),
    .io_ins_142(rport_io_ins_142),
    .io_ins_143(rport_io_ins_143),
    .io_ins_144(rport_io_ins_144),
    .io_ins_145(rport_io_ins_145),
    .io_ins_146(rport_io_ins_146),
    .io_ins_147(rport_io_ins_147),
    .io_ins_148(rport_io_ins_148),
    .io_ins_149(rport_io_ins_149),
    .io_ins_150(rport_io_ins_150),
    .io_ins_151(rport_io_ins_151),
    .io_ins_152(rport_io_ins_152),
    .io_ins_153(rport_io_ins_153),
    .io_ins_154(rport_io_ins_154),
    .io_ins_155(rport_io_ins_155),
    .io_ins_156(rport_io_ins_156),
    .io_ins_157(rport_io_ins_157),
    .io_ins_158(rport_io_ins_158),
    .io_ins_159(rport_io_ins_159),
    .io_ins_160(rport_io_ins_160),
    .io_ins_161(rport_io_ins_161),
    .io_ins_162(rport_io_ins_162),
    .io_ins_163(rport_io_ins_163),
    .io_ins_164(rport_io_ins_164),
    .io_ins_165(rport_io_ins_165),
    .io_ins_166(rport_io_ins_166),
    .io_ins_167(rport_io_ins_167),
    .io_ins_168(rport_io_ins_168),
    .io_ins_169(rport_io_ins_169),
    .io_ins_170(rport_io_ins_170),
    .io_ins_171(rport_io_ins_171),
    .io_ins_172(rport_io_ins_172),
    .io_ins_173(rport_io_ins_173),
    .io_ins_174(rport_io_ins_174),
    .io_ins_175(rport_io_ins_175),
    .io_ins_176(rport_io_ins_176),
    .io_ins_177(rport_io_ins_177),
    .io_ins_178(rport_io_ins_178),
    .io_ins_179(rport_io_ins_179),
    .io_ins_180(rport_io_ins_180),
    .io_ins_181(rport_io_ins_181),
    .io_ins_182(rport_io_ins_182),
    .io_ins_183(rport_io_ins_183),
    .io_ins_184(rport_io_ins_184),
    .io_ins_185(rport_io_ins_185),
    .io_ins_186(rport_io_ins_186),
    .io_ins_187(rport_io_ins_187),
    .io_ins_188(rport_io_ins_188),
    .io_ins_189(rport_io_ins_189),
    .io_ins_190(rport_io_ins_190),
    .io_ins_191(rport_io_ins_191),
    .io_ins_192(rport_io_ins_192),
    .io_ins_193(rport_io_ins_193),
    .io_ins_194(rport_io_ins_194),
    .io_ins_195(rport_io_ins_195),
    .io_ins_196(rport_io_ins_196),
    .io_ins_197(rport_io_ins_197),
    .io_ins_198(rport_io_ins_198),
    .io_ins_199(rport_io_ins_199),
    .io_ins_200(rport_io_ins_200),
    .io_ins_201(rport_io_ins_201),
    .io_ins_202(rport_io_ins_202),
    .io_ins_203(rport_io_ins_203),
    .io_ins_204(rport_io_ins_204),
    .io_ins_205(rport_io_ins_205),
    .io_ins_206(rport_io_ins_206),
    .io_ins_207(rport_io_ins_207),
    .io_ins_208(rport_io_ins_208),
    .io_ins_209(rport_io_ins_209),
    .io_ins_210(rport_io_ins_210),
    .io_ins_211(rport_io_ins_211),
    .io_ins_212(rport_io_ins_212),
    .io_ins_213(rport_io_ins_213),
    .io_ins_214(rport_io_ins_214),
    .io_ins_215(rport_io_ins_215),
    .io_ins_216(rport_io_ins_216),
    .io_ins_217(rport_io_ins_217),
    .io_ins_218(rport_io_ins_218),
    .io_ins_219(rport_io_ins_219),
    .io_ins_220(rport_io_ins_220),
    .io_ins_221(rport_io_ins_221),
    .io_ins_222(rport_io_ins_222),
    .io_ins_223(rport_io_ins_223),
    .io_ins_224(rport_io_ins_224),
    .io_ins_225(rport_io_ins_225),
    .io_ins_226(rport_io_ins_226),
    .io_ins_227(rport_io_ins_227),
    .io_ins_228(rport_io_ins_228),
    .io_ins_229(rport_io_ins_229),
    .io_ins_230(rport_io_ins_230),
    .io_ins_231(rport_io_ins_231),
    .io_ins_232(rport_io_ins_232),
    .io_ins_233(rport_io_ins_233),
    .io_ins_234(rport_io_ins_234),
    .io_ins_235(rport_io_ins_235),
    .io_ins_236(rport_io_ins_236),
    .io_ins_237(rport_io_ins_237),
    .io_ins_238(rport_io_ins_238),
    .io_ins_239(rport_io_ins_239),
    .io_ins_240(rport_io_ins_240),
    .io_ins_241(rport_io_ins_241),
    .io_ins_242(rport_io_ins_242),
    .io_ins_243(rport_io_ins_243),
    .io_ins_244(rport_io_ins_244),
    .io_ins_245(rport_io_ins_245),
    .io_ins_246(rport_io_ins_246),
    .io_ins_247(rport_io_ins_247),
    .io_ins_248(rport_io_ins_248),
    .io_ins_249(rport_io_ins_249),
    .io_ins_250(rport_io_ins_250),
    .io_ins_251(rport_io_ins_251),
    .io_ins_252(rport_io_ins_252),
    .io_ins_253(rport_io_ins_253),
    .io_ins_254(rport_io_ins_254),
    .io_ins_255(rport_io_ins_255),
    .io_ins_256(rport_io_ins_256),
    .io_ins_257(rport_io_ins_257),
    .io_ins_258(rport_io_ins_258),
    .io_ins_259(rport_io_ins_259),
    .io_ins_260(rport_io_ins_260),
    .io_ins_261(rport_io_ins_261),
    .io_ins_262(rport_io_ins_262),
    .io_ins_263(rport_io_ins_263),
    .io_ins_264(rport_io_ins_264),
    .io_ins_265(rport_io_ins_265),
    .io_ins_266(rport_io_ins_266),
    .io_ins_267(rport_io_ins_267),
    .io_ins_268(rport_io_ins_268),
    .io_ins_269(rport_io_ins_269),
    .io_ins_270(rport_io_ins_270),
    .io_ins_271(rport_io_ins_271),
    .io_ins_272(rport_io_ins_272),
    .io_ins_273(rport_io_ins_273),
    .io_ins_274(rport_io_ins_274),
    .io_ins_275(rport_io_ins_275),
    .io_ins_276(rport_io_ins_276),
    .io_ins_277(rport_io_ins_277),
    .io_ins_278(rport_io_ins_278),
    .io_ins_279(rport_io_ins_279),
    .io_ins_280(rport_io_ins_280),
    .io_ins_281(rport_io_ins_281),
    .io_ins_282(rport_io_ins_282),
    .io_ins_283(rport_io_ins_283),
    .io_ins_284(rport_io_ins_284),
    .io_ins_285(rport_io_ins_285),
    .io_ins_286(rport_io_ins_286),
    .io_ins_287(rport_io_ins_287),
    .io_ins_288(rport_io_ins_288),
    .io_ins_289(rport_io_ins_289),
    .io_ins_290(rport_io_ins_290),
    .io_ins_291(rport_io_ins_291),
    .io_ins_292(rport_io_ins_292),
    .io_ins_293(rport_io_ins_293),
    .io_ins_294(rport_io_ins_294),
    .io_ins_295(rport_io_ins_295),
    .io_ins_296(rport_io_ins_296),
    .io_ins_297(rport_io_ins_297),
    .io_ins_298(rport_io_ins_298),
    .io_ins_299(rport_io_ins_299),
    .io_ins_300(rport_io_ins_300),
    .io_ins_301(rport_io_ins_301),
    .io_ins_302(rport_io_ins_302),
    .io_ins_303(rport_io_ins_303),
    .io_ins_304(rport_io_ins_304),
    .io_ins_305(rport_io_ins_305),
    .io_ins_306(rport_io_ins_306),
    .io_ins_307(rport_io_ins_307),
    .io_ins_308(rport_io_ins_308),
    .io_ins_309(rport_io_ins_309),
    .io_ins_310(rport_io_ins_310),
    .io_ins_311(rport_io_ins_311),
    .io_ins_312(rport_io_ins_312),
    .io_ins_313(rport_io_ins_313),
    .io_ins_314(rport_io_ins_314),
    .io_ins_315(rport_io_ins_315),
    .io_ins_316(rport_io_ins_316),
    .io_ins_317(rport_io_ins_317),
    .io_ins_318(rport_io_ins_318),
    .io_ins_319(rport_io_ins_319),
    .io_ins_320(rport_io_ins_320),
    .io_ins_321(rport_io_ins_321),
    .io_ins_322(rport_io_ins_322),
    .io_ins_323(rport_io_ins_323),
    .io_ins_324(rport_io_ins_324),
    .io_ins_325(rport_io_ins_325),
    .io_ins_326(rport_io_ins_326),
    .io_ins_327(rport_io_ins_327),
    .io_ins_328(rport_io_ins_328),
    .io_ins_329(rport_io_ins_329),
    .io_ins_330(rport_io_ins_330),
    .io_ins_331(rport_io_ins_331),
    .io_ins_332(rport_io_ins_332),
    .io_ins_333(rport_io_ins_333),
    .io_ins_334(rport_io_ins_334),
    .io_ins_335(rport_io_ins_335),
    .io_ins_336(rport_io_ins_336),
    .io_ins_337(rport_io_ins_337),
    .io_ins_338(rport_io_ins_338),
    .io_ins_339(rport_io_ins_339),
    .io_ins_340(rport_io_ins_340),
    .io_ins_341(rport_io_ins_341),
    .io_ins_342(rport_io_ins_342),
    .io_ins_343(rport_io_ins_343),
    .io_ins_344(rport_io_ins_344),
    .io_ins_345(rport_io_ins_345),
    .io_ins_346(rport_io_ins_346),
    .io_ins_347(rport_io_ins_347),
    .io_ins_348(rport_io_ins_348),
    .io_ins_349(rport_io_ins_349),
    .io_ins_350(rport_io_ins_350),
    .io_ins_351(rport_io_ins_351),
    .io_ins_352(rport_io_ins_352),
    .io_ins_353(rport_io_ins_353),
    .io_ins_354(rport_io_ins_354),
    .io_ins_355(rport_io_ins_355),
    .io_ins_356(rport_io_ins_356),
    .io_ins_357(rport_io_ins_357),
    .io_ins_358(rport_io_ins_358),
    .io_ins_359(rport_io_ins_359),
    .io_ins_360(rport_io_ins_360),
    .io_ins_361(rport_io_ins_361),
    .io_ins_362(rport_io_ins_362),
    .io_ins_363(rport_io_ins_363),
    .io_ins_364(rport_io_ins_364),
    .io_ins_365(rport_io_ins_365),
    .io_ins_366(rport_io_ins_366),
    .io_ins_367(rport_io_ins_367),
    .io_ins_368(rport_io_ins_368),
    .io_ins_369(rport_io_ins_369),
    .io_ins_370(rport_io_ins_370),
    .io_ins_371(rport_io_ins_371),
    .io_ins_372(rport_io_ins_372),
    .io_ins_373(rport_io_ins_373),
    .io_ins_374(rport_io_ins_374),
    .io_ins_375(rport_io_ins_375),
    .io_ins_376(rport_io_ins_376),
    .io_ins_377(rport_io_ins_377),
    .io_ins_378(rport_io_ins_378),
    .io_ins_379(rport_io_ins_379),
    .io_ins_380(rport_io_ins_380),
    .io_ins_381(rport_io_ins_381),
    .io_ins_382(rport_io_ins_382),
    .io_ins_383(rport_io_ins_383),
    .io_ins_384(rport_io_ins_384),
    .io_ins_385(rport_io_ins_385),
    .io_ins_386(rport_io_ins_386),
    .io_ins_387(rport_io_ins_387),
    .io_ins_388(rport_io_ins_388),
    .io_ins_389(rport_io_ins_389),
    .io_ins_390(rport_io_ins_390),
    .io_ins_391(rport_io_ins_391),
    .io_ins_392(rport_io_ins_392),
    .io_ins_393(rport_io_ins_393),
    .io_ins_394(rport_io_ins_394),
    .io_ins_395(rport_io_ins_395),
    .io_ins_396(rport_io_ins_396),
    .io_ins_397(rport_io_ins_397),
    .io_ins_398(rport_io_ins_398),
    .io_ins_399(rport_io_ins_399),
    .io_ins_400(rport_io_ins_400),
    .io_ins_401(rport_io_ins_401),
    .io_ins_402(rport_io_ins_402),
    .io_ins_403(rport_io_ins_403),
    .io_ins_404(rport_io_ins_404),
    .io_ins_405(rport_io_ins_405),
    .io_ins_406(rport_io_ins_406),
    .io_ins_407(rport_io_ins_407),
    .io_ins_408(rport_io_ins_408),
    .io_ins_409(rport_io_ins_409),
    .io_ins_410(rport_io_ins_410),
    .io_ins_411(rport_io_ins_411),
    .io_ins_412(rport_io_ins_412),
    .io_ins_413(rport_io_ins_413),
    .io_ins_414(rport_io_ins_414),
    .io_ins_415(rport_io_ins_415),
    .io_ins_416(rport_io_ins_416),
    .io_ins_417(rport_io_ins_417),
    .io_ins_418(rport_io_ins_418),
    .io_ins_419(rport_io_ins_419),
    .io_ins_420(rport_io_ins_420),
    .io_ins_421(rport_io_ins_421),
    .io_ins_422(rport_io_ins_422),
    .io_ins_423(rport_io_ins_423),
    .io_ins_424(rport_io_ins_424),
    .io_ins_425(rport_io_ins_425),
    .io_ins_426(rport_io_ins_426),
    .io_ins_427(rport_io_ins_427),
    .io_ins_428(rport_io_ins_428),
    .io_ins_429(rport_io_ins_429),
    .io_ins_430(rport_io_ins_430),
    .io_ins_431(rport_io_ins_431),
    .io_ins_432(rport_io_ins_432),
    .io_ins_433(rport_io_ins_433),
    .io_ins_434(rport_io_ins_434),
    .io_ins_435(rport_io_ins_435),
    .io_ins_436(rport_io_ins_436),
    .io_ins_437(rport_io_ins_437),
    .io_ins_438(rport_io_ins_438),
    .io_ins_439(rport_io_ins_439),
    .io_ins_440(rport_io_ins_440),
    .io_ins_441(rport_io_ins_441),
    .io_ins_442(rport_io_ins_442),
    .io_ins_443(rport_io_ins_443),
    .io_ins_444(rport_io_ins_444),
    .io_ins_445(rport_io_ins_445),
    .io_ins_446(rport_io_ins_446),
    .io_ins_447(rport_io_ins_447),
    .io_ins_448(rport_io_ins_448),
    .io_ins_449(rport_io_ins_449),
    .io_ins_450(rport_io_ins_450),
    .io_ins_451(rport_io_ins_451),
    .io_ins_452(rport_io_ins_452),
    .io_ins_453(rport_io_ins_453),
    .io_ins_454(rport_io_ins_454),
    .io_ins_455(rport_io_ins_455),
    .io_ins_456(rport_io_ins_456),
    .io_ins_457(rport_io_ins_457),
    .io_ins_458(rport_io_ins_458),
    .io_ins_459(rport_io_ins_459),
    .io_ins_460(rport_io_ins_460),
    .io_ins_461(rport_io_ins_461),
    .io_ins_462(rport_io_ins_462),
    .io_ins_463(rport_io_ins_463),
    .io_ins_464(rport_io_ins_464),
    .io_ins_465(rport_io_ins_465),
    .io_ins_466(rport_io_ins_466),
    .io_ins_467(rport_io_ins_467),
    .io_ins_468(rport_io_ins_468),
    .io_ins_469(rport_io_ins_469),
    .io_ins_470(rport_io_ins_470),
    .io_ins_471(rport_io_ins_471),
    .io_ins_472(rport_io_ins_472),
    .io_ins_473(rport_io_ins_473),
    .io_ins_474(rport_io_ins_474),
    .io_ins_475(rport_io_ins_475),
    .io_ins_476(rport_io_ins_476),
    .io_ins_477(rport_io_ins_477),
    .io_ins_478(rport_io_ins_478),
    .io_ins_479(rport_io_ins_479),
    .io_ins_480(rport_io_ins_480),
    .io_ins_481(rport_io_ins_481),
    .io_ins_482(rport_io_ins_482),
    .io_ins_483(rport_io_ins_483),
    .io_ins_484(rport_io_ins_484),
    .io_ins_485(rport_io_ins_485),
    .io_ins_486(rport_io_ins_486),
    .io_ins_487(rport_io_ins_487),
    .io_ins_488(rport_io_ins_488),
    .io_ins_489(rport_io_ins_489),
    .io_ins_490(rport_io_ins_490),
    .io_ins_491(rport_io_ins_491),
    .io_ins_492(rport_io_ins_492),
    .io_ins_493(rport_io_ins_493),
    .io_ins_494(rport_io_ins_494),
    .io_ins_495(rport_io_ins_495),
    .io_ins_496(rport_io_ins_496),
    .io_ins_497(rport_io_ins_497),
    .io_ins_498(rport_io_ins_498),
    .io_ins_499(rport_io_ins_499),
    .io_ins_500(rport_io_ins_500),
    .io_ins_501(rport_io_ins_501),
    .io_ins_502(rport_io_ins_502),
    .io_sel(rport_io_sel),
    .io_out(rport_io_out)
  );
  assign _T_3076 = io_waddr == 32'h0; // @[RegFile.scala 80:42:@34258.4]
  assign _T_3082 = io_waddr == 32'h1; // @[RegFile.scala 68:46:@34270.4]
  assign _T_3083 = io_wen & _T_3082; // @[RegFile.scala 68:34:@34271.4]
  assign _T_3096 = io_waddr == 32'h2; // @[RegFile.scala 80:42:@34289.4]
  assign _T_3102 = io_waddr == 32'h3; // @[RegFile.scala 74:80:@34301.4]
  assign _T_3103 = io_wen & _T_3102; // @[RegFile.scala 74:68:@34302.4]
  assign io_rdata = rport_io_out; // @[RegFile.scala 107:14:@42309.4]
  assign io_argIns_0 = regs_0_io_out; // @[RegFile.scala 111:13:@42314.4]
  assign io_argIns_1 = regs_1_io_out; // @[RegFile.scala 111:13:@42315.4]
  assign io_argIns_2 = regs_2_io_out; // @[RegFile.scala 111:13:@42316.4]
  assign regs_0_clock = clock; // @[:@34256.4]
  assign regs_0_reset = reset; // @[:@34257.4 RegFile.scala 82:16:@34263.4]
  assign regs_0_io_in = io_wdata; // @[RegFile.scala 81:16:@34261.4]
  assign regs_0_io_reset = reset; // @[RegFile.scala 83:19:@34265.4]
  assign regs_0_io_enable = io_wen & _T_3076; // @[RegFile.scala 80:20:@34260.4]
  assign regs_1_clock = clock; // @[:@34268.4]
  assign regs_1_reset = reset; // @[:@34269.4 RegFile.scala 70:16:@34281.4]
  assign regs_1_io_in = _T_3083 ? io_wdata : io_argOuts_0_bits; // @[RegFile.scala 69:16:@34279.4]
  assign regs_1_io_reset = reset; // @[RegFile.scala 72:19:@34284.4]
  assign regs_1_io_enable = _T_3083 ? _T_3083 : io_argOuts_0_valid; // @[RegFile.scala 68:20:@34275.4]
  assign regs_2_clock = clock; // @[:@34287.4]
  assign regs_2_reset = reset; // @[:@34288.4 RegFile.scala 82:16:@34294.4]
  assign regs_2_io_in = io_wdata; // @[RegFile.scala 81:16:@34292.4]
  assign regs_2_io_reset = reset; // @[RegFile.scala 83:19:@34296.4]
  assign regs_2_io_enable = io_wen & _T_3096; // @[RegFile.scala 80:20:@34291.4]
  assign regs_3_clock = clock; // @[:@34299.4]
  assign regs_3_reset = io_reset; // @[:@34300.4 RegFile.scala 76:16:@34307.4]
  assign regs_3_io_in = io_argOuts_1_valid ? io_argOuts_1_bits : io_wdata; // @[RegFile.scala 75:16:@34306.4]
  assign regs_3_io_reset = reset; // @[RegFile.scala 78:19:@34310.4]
  assign regs_3_io_enable = io_argOuts_1_valid | _T_3103; // @[RegFile.scala 74:20:@34304.4]
  assign regs_4_clock = clock; // @[:@34313.4]
  assign regs_4_reset = io_reset; // @[:@34314.4 RegFile.scala 76:16:@34321.4]
  assign regs_4_io_in = 64'h0; // @[RegFile.scala 75:16:@34320.4]
  assign regs_4_io_reset = reset; // @[RegFile.scala 78:19:@34324.4]
  assign regs_4_io_enable = 1'h1; // @[RegFile.scala 74:20:@34318.4]
  assign regs_5_clock = clock; // @[:@34327.4]
  assign regs_5_reset = io_reset; // @[:@34328.4 RegFile.scala 76:16:@34335.4]
  assign regs_5_io_in = 64'h0; // @[RegFile.scala 75:16:@34334.4]
  assign regs_5_io_reset = reset; // @[RegFile.scala 78:19:@34338.4]
  assign regs_5_io_enable = 1'h1; // @[RegFile.scala 74:20:@34332.4]
  assign regs_6_clock = clock; // @[:@34341.4]
  assign regs_6_reset = io_reset; // @[:@34342.4 RegFile.scala 76:16:@34349.4]
  assign regs_6_io_in = 64'h0; // @[RegFile.scala 75:16:@34348.4]
  assign regs_6_io_reset = reset; // @[RegFile.scala 78:19:@34352.4]
  assign regs_6_io_enable = 1'h1; // @[RegFile.scala 74:20:@34346.4]
  assign regs_7_clock = clock; // @[:@34355.4]
  assign regs_7_reset = io_reset; // @[:@34356.4 RegFile.scala 76:16:@34363.4]
  assign regs_7_io_in = 64'h0; // @[RegFile.scala 75:16:@34362.4]
  assign regs_7_io_reset = reset; // @[RegFile.scala 78:19:@34366.4]
  assign regs_7_io_enable = 1'h1; // @[RegFile.scala 74:20:@34360.4]
  assign regs_8_clock = clock; // @[:@34369.4]
  assign regs_8_reset = io_reset; // @[:@34370.4 RegFile.scala 76:16:@34377.4]
  assign regs_8_io_in = 64'h0; // @[RegFile.scala 75:16:@34376.4]
  assign regs_8_io_reset = reset; // @[RegFile.scala 78:19:@34380.4]
  assign regs_8_io_enable = 1'h1; // @[RegFile.scala 74:20:@34374.4]
  assign regs_9_clock = clock; // @[:@34383.4]
  assign regs_9_reset = io_reset; // @[:@34384.4 RegFile.scala 76:16:@34391.4]
  assign regs_9_io_in = 64'h0; // @[RegFile.scala 75:16:@34390.4]
  assign regs_9_io_reset = reset; // @[RegFile.scala 78:19:@34394.4]
  assign regs_9_io_enable = 1'h1; // @[RegFile.scala 74:20:@34388.4]
  assign regs_10_clock = clock; // @[:@34397.4]
  assign regs_10_reset = io_reset; // @[:@34398.4 RegFile.scala 76:16:@34405.4]
  assign regs_10_io_in = 64'h0; // @[RegFile.scala 75:16:@34404.4]
  assign regs_10_io_reset = reset; // @[RegFile.scala 78:19:@34408.4]
  assign regs_10_io_enable = 1'h1; // @[RegFile.scala 74:20:@34402.4]
  assign regs_11_clock = clock; // @[:@34411.4]
  assign regs_11_reset = io_reset; // @[:@34412.4 RegFile.scala 76:16:@34419.4]
  assign regs_11_io_in = 64'h0; // @[RegFile.scala 75:16:@34418.4]
  assign regs_11_io_reset = reset; // @[RegFile.scala 78:19:@34422.4]
  assign regs_11_io_enable = 1'h1; // @[RegFile.scala 74:20:@34416.4]
  assign regs_12_clock = clock; // @[:@34425.4]
  assign regs_12_reset = io_reset; // @[:@34426.4 RegFile.scala 76:16:@34433.4]
  assign regs_12_io_in = 64'h0; // @[RegFile.scala 75:16:@34432.4]
  assign regs_12_io_reset = reset; // @[RegFile.scala 78:19:@34436.4]
  assign regs_12_io_enable = 1'h1; // @[RegFile.scala 74:20:@34430.4]
  assign regs_13_clock = clock; // @[:@34439.4]
  assign regs_13_reset = io_reset; // @[:@34440.4 RegFile.scala 76:16:@34447.4]
  assign regs_13_io_in = 64'h0; // @[RegFile.scala 75:16:@34446.4]
  assign regs_13_io_reset = reset; // @[RegFile.scala 78:19:@34450.4]
  assign regs_13_io_enable = 1'h1; // @[RegFile.scala 74:20:@34444.4]
  assign regs_14_clock = clock; // @[:@34453.4]
  assign regs_14_reset = io_reset; // @[:@34454.4 RegFile.scala 76:16:@34461.4]
  assign regs_14_io_in = 64'h0; // @[RegFile.scala 75:16:@34460.4]
  assign regs_14_io_reset = reset; // @[RegFile.scala 78:19:@34464.4]
  assign regs_14_io_enable = 1'h1; // @[RegFile.scala 74:20:@34458.4]
  assign regs_15_clock = clock; // @[:@34467.4]
  assign regs_15_reset = io_reset; // @[:@34468.4 RegFile.scala 76:16:@34475.4]
  assign regs_15_io_in = 64'h0; // @[RegFile.scala 75:16:@34474.4]
  assign regs_15_io_reset = reset; // @[RegFile.scala 78:19:@34478.4]
  assign regs_15_io_enable = 1'h1; // @[RegFile.scala 74:20:@34472.4]
  assign regs_16_clock = clock; // @[:@34481.4]
  assign regs_16_reset = io_reset; // @[:@34482.4 RegFile.scala 76:16:@34489.4]
  assign regs_16_io_in = 64'h0; // @[RegFile.scala 75:16:@34488.4]
  assign regs_16_io_reset = reset; // @[RegFile.scala 78:19:@34492.4]
  assign regs_16_io_enable = 1'h1; // @[RegFile.scala 74:20:@34486.4]
  assign regs_17_clock = clock; // @[:@34495.4]
  assign regs_17_reset = io_reset; // @[:@34496.4 RegFile.scala 76:16:@34503.4]
  assign regs_17_io_in = 64'h0; // @[RegFile.scala 75:16:@34502.4]
  assign regs_17_io_reset = reset; // @[RegFile.scala 78:19:@34506.4]
  assign regs_17_io_enable = 1'h1; // @[RegFile.scala 74:20:@34500.4]
  assign regs_18_clock = clock; // @[:@34509.4]
  assign regs_18_reset = io_reset; // @[:@34510.4 RegFile.scala 76:16:@34517.4]
  assign regs_18_io_in = 64'h0; // @[RegFile.scala 75:16:@34516.4]
  assign regs_18_io_reset = reset; // @[RegFile.scala 78:19:@34520.4]
  assign regs_18_io_enable = 1'h1; // @[RegFile.scala 74:20:@34514.4]
  assign regs_19_clock = clock; // @[:@34523.4]
  assign regs_19_reset = io_reset; // @[:@34524.4 RegFile.scala 76:16:@34531.4]
  assign regs_19_io_in = 64'h0; // @[RegFile.scala 75:16:@34530.4]
  assign regs_19_io_reset = reset; // @[RegFile.scala 78:19:@34534.4]
  assign regs_19_io_enable = 1'h1; // @[RegFile.scala 74:20:@34528.4]
  assign regs_20_clock = clock; // @[:@34537.4]
  assign regs_20_reset = io_reset; // @[:@34538.4 RegFile.scala 76:16:@34545.4]
  assign regs_20_io_in = 64'h0; // @[RegFile.scala 75:16:@34544.4]
  assign regs_20_io_reset = reset; // @[RegFile.scala 78:19:@34548.4]
  assign regs_20_io_enable = 1'h1; // @[RegFile.scala 74:20:@34542.4]
  assign regs_21_clock = clock; // @[:@34551.4]
  assign regs_21_reset = io_reset; // @[:@34552.4 RegFile.scala 76:16:@34559.4]
  assign regs_21_io_in = 64'h0; // @[RegFile.scala 75:16:@34558.4]
  assign regs_21_io_reset = reset; // @[RegFile.scala 78:19:@34562.4]
  assign regs_21_io_enable = 1'h1; // @[RegFile.scala 74:20:@34556.4]
  assign regs_22_clock = clock; // @[:@34565.4]
  assign regs_22_reset = io_reset; // @[:@34566.4 RegFile.scala 76:16:@34573.4]
  assign regs_22_io_in = 64'h0; // @[RegFile.scala 75:16:@34572.4]
  assign regs_22_io_reset = reset; // @[RegFile.scala 78:19:@34576.4]
  assign regs_22_io_enable = 1'h1; // @[RegFile.scala 74:20:@34570.4]
  assign regs_23_clock = clock; // @[:@34579.4]
  assign regs_23_reset = io_reset; // @[:@34580.4 RegFile.scala 76:16:@34587.4]
  assign regs_23_io_in = 64'h0; // @[RegFile.scala 75:16:@34586.4]
  assign regs_23_io_reset = reset; // @[RegFile.scala 78:19:@34590.4]
  assign regs_23_io_enable = 1'h1; // @[RegFile.scala 74:20:@34584.4]
  assign regs_24_clock = clock; // @[:@34593.4]
  assign regs_24_reset = io_reset; // @[:@34594.4 RegFile.scala 76:16:@34601.4]
  assign regs_24_io_in = 64'h0; // @[RegFile.scala 75:16:@34600.4]
  assign regs_24_io_reset = reset; // @[RegFile.scala 78:19:@34604.4]
  assign regs_24_io_enable = 1'h1; // @[RegFile.scala 74:20:@34598.4]
  assign regs_25_clock = clock; // @[:@34607.4]
  assign regs_25_reset = io_reset; // @[:@34608.4 RegFile.scala 76:16:@34615.4]
  assign regs_25_io_in = 64'h0; // @[RegFile.scala 75:16:@34614.4]
  assign regs_25_io_reset = reset; // @[RegFile.scala 78:19:@34618.4]
  assign regs_25_io_enable = 1'h1; // @[RegFile.scala 74:20:@34612.4]
  assign regs_26_clock = clock; // @[:@34621.4]
  assign regs_26_reset = io_reset; // @[:@34622.4 RegFile.scala 76:16:@34629.4]
  assign regs_26_io_in = 64'h0; // @[RegFile.scala 75:16:@34628.4]
  assign regs_26_io_reset = reset; // @[RegFile.scala 78:19:@34632.4]
  assign regs_26_io_enable = 1'h1; // @[RegFile.scala 74:20:@34626.4]
  assign regs_27_clock = clock; // @[:@34635.4]
  assign regs_27_reset = io_reset; // @[:@34636.4 RegFile.scala 76:16:@34643.4]
  assign regs_27_io_in = 64'h0; // @[RegFile.scala 75:16:@34642.4]
  assign regs_27_io_reset = reset; // @[RegFile.scala 78:19:@34646.4]
  assign regs_27_io_enable = 1'h1; // @[RegFile.scala 74:20:@34640.4]
  assign regs_28_clock = clock; // @[:@34649.4]
  assign regs_28_reset = io_reset; // @[:@34650.4 RegFile.scala 76:16:@34657.4]
  assign regs_28_io_in = 64'h0; // @[RegFile.scala 75:16:@34656.4]
  assign regs_28_io_reset = reset; // @[RegFile.scala 78:19:@34660.4]
  assign regs_28_io_enable = 1'h1; // @[RegFile.scala 74:20:@34654.4]
  assign regs_29_clock = clock; // @[:@34663.4]
  assign regs_29_reset = io_reset; // @[:@34664.4 RegFile.scala 76:16:@34671.4]
  assign regs_29_io_in = 64'h0; // @[RegFile.scala 75:16:@34670.4]
  assign regs_29_io_reset = reset; // @[RegFile.scala 78:19:@34674.4]
  assign regs_29_io_enable = 1'h1; // @[RegFile.scala 74:20:@34668.4]
  assign regs_30_clock = clock; // @[:@34677.4]
  assign regs_30_reset = io_reset; // @[:@34678.4 RegFile.scala 76:16:@34685.4]
  assign regs_30_io_in = 64'h0; // @[RegFile.scala 75:16:@34684.4]
  assign regs_30_io_reset = reset; // @[RegFile.scala 78:19:@34688.4]
  assign regs_30_io_enable = 1'h1; // @[RegFile.scala 74:20:@34682.4]
  assign regs_31_clock = clock; // @[:@34691.4]
  assign regs_31_reset = io_reset; // @[:@34692.4 RegFile.scala 76:16:@34699.4]
  assign regs_31_io_in = 64'h0; // @[RegFile.scala 75:16:@34698.4]
  assign regs_31_io_reset = reset; // @[RegFile.scala 78:19:@34702.4]
  assign regs_31_io_enable = 1'h1; // @[RegFile.scala 74:20:@34696.4]
  assign regs_32_clock = clock; // @[:@34705.4]
  assign regs_32_reset = io_reset; // @[:@34706.4 RegFile.scala 76:16:@34713.4]
  assign regs_32_io_in = 64'h0; // @[RegFile.scala 75:16:@34712.4]
  assign regs_32_io_reset = reset; // @[RegFile.scala 78:19:@34716.4]
  assign regs_32_io_enable = 1'h1; // @[RegFile.scala 74:20:@34710.4]
  assign regs_33_clock = clock; // @[:@34719.4]
  assign regs_33_reset = io_reset; // @[:@34720.4 RegFile.scala 76:16:@34727.4]
  assign regs_33_io_in = 64'h0; // @[RegFile.scala 75:16:@34726.4]
  assign regs_33_io_reset = reset; // @[RegFile.scala 78:19:@34730.4]
  assign regs_33_io_enable = 1'h1; // @[RegFile.scala 74:20:@34724.4]
  assign regs_34_clock = clock; // @[:@34733.4]
  assign regs_34_reset = io_reset; // @[:@34734.4 RegFile.scala 76:16:@34741.4]
  assign regs_34_io_in = 64'h0; // @[RegFile.scala 75:16:@34740.4]
  assign regs_34_io_reset = reset; // @[RegFile.scala 78:19:@34744.4]
  assign regs_34_io_enable = 1'h1; // @[RegFile.scala 74:20:@34738.4]
  assign regs_35_clock = clock; // @[:@34747.4]
  assign regs_35_reset = io_reset; // @[:@34748.4 RegFile.scala 76:16:@34755.4]
  assign regs_35_io_in = 64'h0; // @[RegFile.scala 75:16:@34754.4]
  assign regs_35_io_reset = reset; // @[RegFile.scala 78:19:@34758.4]
  assign regs_35_io_enable = 1'h1; // @[RegFile.scala 74:20:@34752.4]
  assign regs_36_clock = clock; // @[:@34761.4]
  assign regs_36_reset = io_reset; // @[:@34762.4 RegFile.scala 76:16:@34769.4]
  assign regs_36_io_in = 64'h0; // @[RegFile.scala 75:16:@34768.4]
  assign regs_36_io_reset = reset; // @[RegFile.scala 78:19:@34772.4]
  assign regs_36_io_enable = 1'h1; // @[RegFile.scala 74:20:@34766.4]
  assign regs_37_clock = clock; // @[:@34775.4]
  assign regs_37_reset = io_reset; // @[:@34776.4 RegFile.scala 76:16:@34783.4]
  assign regs_37_io_in = 64'h0; // @[RegFile.scala 75:16:@34782.4]
  assign regs_37_io_reset = reset; // @[RegFile.scala 78:19:@34786.4]
  assign regs_37_io_enable = 1'h1; // @[RegFile.scala 74:20:@34780.4]
  assign regs_38_clock = clock; // @[:@34789.4]
  assign regs_38_reset = io_reset; // @[:@34790.4 RegFile.scala 76:16:@34797.4]
  assign regs_38_io_in = 64'h0; // @[RegFile.scala 75:16:@34796.4]
  assign regs_38_io_reset = reset; // @[RegFile.scala 78:19:@34800.4]
  assign regs_38_io_enable = 1'h1; // @[RegFile.scala 74:20:@34794.4]
  assign regs_39_clock = clock; // @[:@34803.4]
  assign regs_39_reset = io_reset; // @[:@34804.4 RegFile.scala 76:16:@34811.4]
  assign regs_39_io_in = 64'h0; // @[RegFile.scala 75:16:@34810.4]
  assign regs_39_io_reset = reset; // @[RegFile.scala 78:19:@34814.4]
  assign regs_39_io_enable = 1'h1; // @[RegFile.scala 74:20:@34808.4]
  assign regs_40_clock = clock; // @[:@34817.4]
  assign regs_40_reset = io_reset; // @[:@34818.4 RegFile.scala 76:16:@34825.4]
  assign regs_40_io_in = 64'h0; // @[RegFile.scala 75:16:@34824.4]
  assign regs_40_io_reset = reset; // @[RegFile.scala 78:19:@34828.4]
  assign regs_40_io_enable = 1'h1; // @[RegFile.scala 74:20:@34822.4]
  assign regs_41_clock = clock; // @[:@34831.4]
  assign regs_41_reset = io_reset; // @[:@34832.4 RegFile.scala 76:16:@34839.4]
  assign regs_41_io_in = 64'h0; // @[RegFile.scala 75:16:@34838.4]
  assign regs_41_io_reset = reset; // @[RegFile.scala 78:19:@34842.4]
  assign regs_41_io_enable = 1'h1; // @[RegFile.scala 74:20:@34836.4]
  assign regs_42_clock = clock; // @[:@34845.4]
  assign regs_42_reset = io_reset; // @[:@34846.4 RegFile.scala 76:16:@34853.4]
  assign regs_42_io_in = 64'h0; // @[RegFile.scala 75:16:@34852.4]
  assign regs_42_io_reset = reset; // @[RegFile.scala 78:19:@34856.4]
  assign regs_42_io_enable = 1'h1; // @[RegFile.scala 74:20:@34850.4]
  assign regs_43_clock = clock; // @[:@34859.4]
  assign regs_43_reset = io_reset; // @[:@34860.4 RegFile.scala 76:16:@34867.4]
  assign regs_43_io_in = 64'h0; // @[RegFile.scala 75:16:@34866.4]
  assign regs_43_io_reset = reset; // @[RegFile.scala 78:19:@34870.4]
  assign regs_43_io_enable = 1'h1; // @[RegFile.scala 74:20:@34864.4]
  assign regs_44_clock = clock; // @[:@34873.4]
  assign regs_44_reset = io_reset; // @[:@34874.4 RegFile.scala 76:16:@34881.4]
  assign regs_44_io_in = 64'h0; // @[RegFile.scala 75:16:@34880.4]
  assign regs_44_io_reset = reset; // @[RegFile.scala 78:19:@34884.4]
  assign regs_44_io_enable = 1'h1; // @[RegFile.scala 74:20:@34878.4]
  assign regs_45_clock = clock; // @[:@34887.4]
  assign regs_45_reset = io_reset; // @[:@34888.4 RegFile.scala 76:16:@34895.4]
  assign regs_45_io_in = 64'h0; // @[RegFile.scala 75:16:@34894.4]
  assign regs_45_io_reset = reset; // @[RegFile.scala 78:19:@34898.4]
  assign regs_45_io_enable = 1'h1; // @[RegFile.scala 74:20:@34892.4]
  assign regs_46_clock = clock; // @[:@34901.4]
  assign regs_46_reset = io_reset; // @[:@34902.4 RegFile.scala 76:16:@34909.4]
  assign regs_46_io_in = 64'h0; // @[RegFile.scala 75:16:@34908.4]
  assign regs_46_io_reset = reset; // @[RegFile.scala 78:19:@34912.4]
  assign regs_46_io_enable = 1'h1; // @[RegFile.scala 74:20:@34906.4]
  assign regs_47_clock = clock; // @[:@34915.4]
  assign regs_47_reset = io_reset; // @[:@34916.4 RegFile.scala 76:16:@34923.4]
  assign regs_47_io_in = 64'h0; // @[RegFile.scala 75:16:@34922.4]
  assign regs_47_io_reset = reset; // @[RegFile.scala 78:19:@34926.4]
  assign regs_47_io_enable = 1'h1; // @[RegFile.scala 74:20:@34920.4]
  assign regs_48_clock = clock; // @[:@34929.4]
  assign regs_48_reset = io_reset; // @[:@34930.4 RegFile.scala 76:16:@34937.4]
  assign regs_48_io_in = 64'h0; // @[RegFile.scala 75:16:@34936.4]
  assign regs_48_io_reset = reset; // @[RegFile.scala 78:19:@34940.4]
  assign regs_48_io_enable = 1'h1; // @[RegFile.scala 74:20:@34934.4]
  assign regs_49_clock = clock; // @[:@34943.4]
  assign regs_49_reset = io_reset; // @[:@34944.4 RegFile.scala 76:16:@34951.4]
  assign regs_49_io_in = 64'h0; // @[RegFile.scala 75:16:@34950.4]
  assign regs_49_io_reset = reset; // @[RegFile.scala 78:19:@34954.4]
  assign regs_49_io_enable = 1'h1; // @[RegFile.scala 74:20:@34948.4]
  assign regs_50_clock = clock; // @[:@34957.4]
  assign regs_50_reset = io_reset; // @[:@34958.4 RegFile.scala 76:16:@34965.4]
  assign regs_50_io_in = 64'h0; // @[RegFile.scala 75:16:@34964.4]
  assign regs_50_io_reset = reset; // @[RegFile.scala 78:19:@34968.4]
  assign regs_50_io_enable = 1'h1; // @[RegFile.scala 74:20:@34962.4]
  assign regs_51_clock = clock; // @[:@34971.4]
  assign regs_51_reset = io_reset; // @[:@34972.4 RegFile.scala 76:16:@34979.4]
  assign regs_51_io_in = 64'h0; // @[RegFile.scala 75:16:@34978.4]
  assign regs_51_io_reset = reset; // @[RegFile.scala 78:19:@34982.4]
  assign regs_51_io_enable = 1'h1; // @[RegFile.scala 74:20:@34976.4]
  assign regs_52_clock = clock; // @[:@34985.4]
  assign regs_52_reset = io_reset; // @[:@34986.4 RegFile.scala 76:16:@34993.4]
  assign regs_52_io_in = 64'h0; // @[RegFile.scala 75:16:@34992.4]
  assign regs_52_io_reset = reset; // @[RegFile.scala 78:19:@34996.4]
  assign regs_52_io_enable = 1'h1; // @[RegFile.scala 74:20:@34990.4]
  assign regs_53_clock = clock; // @[:@34999.4]
  assign regs_53_reset = io_reset; // @[:@35000.4 RegFile.scala 76:16:@35007.4]
  assign regs_53_io_in = 64'h0; // @[RegFile.scala 75:16:@35006.4]
  assign regs_53_io_reset = reset; // @[RegFile.scala 78:19:@35010.4]
  assign regs_53_io_enable = 1'h1; // @[RegFile.scala 74:20:@35004.4]
  assign regs_54_clock = clock; // @[:@35013.4]
  assign regs_54_reset = io_reset; // @[:@35014.4 RegFile.scala 76:16:@35021.4]
  assign regs_54_io_in = 64'h0; // @[RegFile.scala 75:16:@35020.4]
  assign regs_54_io_reset = reset; // @[RegFile.scala 78:19:@35024.4]
  assign regs_54_io_enable = 1'h1; // @[RegFile.scala 74:20:@35018.4]
  assign regs_55_clock = clock; // @[:@35027.4]
  assign regs_55_reset = io_reset; // @[:@35028.4 RegFile.scala 76:16:@35035.4]
  assign regs_55_io_in = 64'h0; // @[RegFile.scala 75:16:@35034.4]
  assign regs_55_io_reset = reset; // @[RegFile.scala 78:19:@35038.4]
  assign regs_55_io_enable = 1'h1; // @[RegFile.scala 74:20:@35032.4]
  assign regs_56_clock = clock; // @[:@35041.4]
  assign regs_56_reset = io_reset; // @[:@35042.4 RegFile.scala 76:16:@35049.4]
  assign regs_56_io_in = 64'h0; // @[RegFile.scala 75:16:@35048.4]
  assign regs_56_io_reset = reset; // @[RegFile.scala 78:19:@35052.4]
  assign regs_56_io_enable = 1'h1; // @[RegFile.scala 74:20:@35046.4]
  assign regs_57_clock = clock; // @[:@35055.4]
  assign regs_57_reset = io_reset; // @[:@35056.4 RegFile.scala 76:16:@35063.4]
  assign regs_57_io_in = 64'h0; // @[RegFile.scala 75:16:@35062.4]
  assign regs_57_io_reset = reset; // @[RegFile.scala 78:19:@35066.4]
  assign regs_57_io_enable = 1'h1; // @[RegFile.scala 74:20:@35060.4]
  assign regs_58_clock = clock; // @[:@35069.4]
  assign regs_58_reset = io_reset; // @[:@35070.4 RegFile.scala 76:16:@35077.4]
  assign regs_58_io_in = 64'h0; // @[RegFile.scala 75:16:@35076.4]
  assign regs_58_io_reset = reset; // @[RegFile.scala 78:19:@35080.4]
  assign regs_58_io_enable = 1'h1; // @[RegFile.scala 74:20:@35074.4]
  assign regs_59_clock = clock; // @[:@35083.4]
  assign regs_59_reset = io_reset; // @[:@35084.4 RegFile.scala 76:16:@35091.4]
  assign regs_59_io_in = 64'h0; // @[RegFile.scala 75:16:@35090.4]
  assign regs_59_io_reset = reset; // @[RegFile.scala 78:19:@35094.4]
  assign regs_59_io_enable = 1'h1; // @[RegFile.scala 74:20:@35088.4]
  assign regs_60_clock = clock; // @[:@35097.4]
  assign regs_60_reset = io_reset; // @[:@35098.4 RegFile.scala 76:16:@35105.4]
  assign regs_60_io_in = 64'h0; // @[RegFile.scala 75:16:@35104.4]
  assign regs_60_io_reset = reset; // @[RegFile.scala 78:19:@35108.4]
  assign regs_60_io_enable = 1'h1; // @[RegFile.scala 74:20:@35102.4]
  assign regs_61_clock = clock; // @[:@35111.4]
  assign regs_61_reset = io_reset; // @[:@35112.4 RegFile.scala 76:16:@35119.4]
  assign regs_61_io_in = 64'h0; // @[RegFile.scala 75:16:@35118.4]
  assign regs_61_io_reset = reset; // @[RegFile.scala 78:19:@35122.4]
  assign regs_61_io_enable = 1'h1; // @[RegFile.scala 74:20:@35116.4]
  assign regs_62_clock = clock; // @[:@35125.4]
  assign regs_62_reset = io_reset; // @[:@35126.4 RegFile.scala 76:16:@35133.4]
  assign regs_62_io_in = 64'h0; // @[RegFile.scala 75:16:@35132.4]
  assign regs_62_io_reset = reset; // @[RegFile.scala 78:19:@35136.4]
  assign regs_62_io_enable = 1'h1; // @[RegFile.scala 74:20:@35130.4]
  assign regs_63_clock = clock; // @[:@35139.4]
  assign regs_63_reset = io_reset; // @[:@35140.4 RegFile.scala 76:16:@35147.4]
  assign regs_63_io_in = 64'h0; // @[RegFile.scala 75:16:@35146.4]
  assign regs_63_io_reset = reset; // @[RegFile.scala 78:19:@35150.4]
  assign regs_63_io_enable = 1'h1; // @[RegFile.scala 74:20:@35144.4]
  assign regs_64_clock = clock; // @[:@35153.4]
  assign regs_64_reset = io_reset; // @[:@35154.4 RegFile.scala 76:16:@35161.4]
  assign regs_64_io_in = 64'h0; // @[RegFile.scala 75:16:@35160.4]
  assign regs_64_io_reset = reset; // @[RegFile.scala 78:19:@35164.4]
  assign regs_64_io_enable = 1'h1; // @[RegFile.scala 74:20:@35158.4]
  assign regs_65_clock = clock; // @[:@35167.4]
  assign regs_65_reset = io_reset; // @[:@35168.4 RegFile.scala 76:16:@35175.4]
  assign regs_65_io_in = 64'h0; // @[RegFile.scala 75:16:@35174.4]
  assign regs_65_io_reset = reset; // @[RegFile.scala 78:19:@35178.4]
  assign regs_65_io_enable = 1'h1; // @[RegFile.scala 74:20:@35172.4]
  assign regs_66_clock = clock; // @[:@35181.4]
  assign regs_66_reset = io_reset; // @[:@35182.4 RegFile.scala 76:16:@35189.4]
  assign regs_66_io_in = 64'h0; // @[RegFile.scala 75:16:@35188.4]
  assign regs_66_io_reset = reset; // @[RegFile.scala 78:19:@35192.4]
  assign regs_66_io_enable = 1'h1; // @[RegFile.scala 74:20:@35186.4]
  assign regs_67_clock = clock; // @[:@35195.4]
  assign regs_67_reset = io_reset; // @[:@35196.4 RegFile.scala 76:16:@35203.4]
  assign regs_67_io_in = 64'h0; // @[RegFile.scala 75:16:@35202.4]
  assign regs_67_io_reset = reset; // @[RegFile.scala 78:19:@35206.4]
  assign regs_67_io_enable = 1'h1; // @[RegFile.scala 74:20:@35200.4]
  assign regs_68_clock = clock; // @[:@35209.4]
  assign regs_68_reset = io_reset; // @[:@35210.4 RegFile.scala 76:16:@35217.4]
  assign regs_68_io_in = 64'h0; // @[RegFile.scala 75:16:@35216.4]
  assign regs_68_io_reset = reset; // @[RegFile.scala 78:19:@35220.4]
  assign regs_68_io_enable = 1'h1; // @[RegFile.scala 74:20:@35214.4]
  assign regs_69_clock = clock; // @[:@35223.4]
  assign regs_69_reset = io_reset; // @[:@35224.4 RegFile.scala 76:16:@35231.4]
  assign regs_69_io_in = 64'h0; // @[RegFile.scala 75:16:@35230.4]
  assign regs_69_io_reset = reset; // @[RegFile.scala 78:19:@35234.4]
  assign regs_69_io_enable = 1'h1; // @[RegFile.scala 74:20:@35228.4]
  assign regs_70_clock = clock; // @[:@35237.4]
  assign regs_70_reset = io_reset; // @[:@35238.4 RegFile.scala 76:16:@35245.4]
  assign regs_70_io_in = 64'h0; // @[RegFile.scala 75:16:@35244.4]
  assign regs_70_io_reset = reset; // @[RegFile.scala 78:19:@35248.4]
  assign regs_70_io_enable = 1'h1; // @[RegFile.scala 74:20:@35242.4]
  assign regs_71_clock = clock; // @[:@35251.4]
  assign regs_71_reset = io_reset; // @[:@35252.4 RegFile.scala 76:16:@35259.4]
  assign regs_71_io_in = 64'h0; // @[RegFile.scala 75:16:@35258.4]
  assign regs_71_io_reset = reset; // @[RegFile.scala 78:19:@35262.4]
  assign regs_71_io_enable = 1'h1; // @[RegFile.scala 74:20:@35256.4]
  assign regs_72_clock = clock; // @[:@35265.4]
  assign regs_72_reset = io_reset; // @[:@35266.4 RegFile.scala 76:16:@35273.4]
  assign regs_72_io_in = 64'h0; // @[RegFile.scala 75:16:@35272.4]
  assign regs_72_io_reset = reset; // @[RegFile.scala 78:19:@35276.4]
  assign regs_72_io_enable = 1'h1; // @[RegFile.scala 74:20:@35270.4]
  assign regs_73_clock = clock; // @[:@35279.4]
  assign regs_73_reset = io_reset; // @[:@35280.4 RegFile.scala 76:16:@35287.4]
  assign regs_73_io_in = 64'h0; // @[RegFile.scala 75:16:@35286.4]
  assign regs_73_io_reset = reset; // @[RegFile.scala 78:19:@35290.4]
  assign regs_73_io_enable = 1'h1; // @[RegFile.scala 74:20:@35284.4]
  assign regs_74_clock = clock; // @[:@35293.4]
  assign regs_74_reset = io_reset; // @[:@35294.4 RegFile.scala 76:16:@35301.4]
  assign regs_74_io_in = 64'h0; // @[RegFile.scala 75:16:@35300.4]
  assign regs_74_io_reset = reset; // @[RegFile.scala 78:19:@35304.4]
  assign regs_74_io_enable = 1'h1; // @[RegFile.scala 74:20:@35298.4]
  assign regs_75_clock = clock; // @[:@35307.4]
  assign regs_75_reset = io_reset; // @[:@35308.4 RegFile.scala 76:16:@35315.4]
  assign regs_75_io_in = 64'h0; // @[RegFile.scala 75:16:@35314.4]
  assign regs_75_io_reset = reset; // @[RegFile.scala 78:19:@35318.4]
  assign regs_75_io_enable = 1'h1; // @[RegFile.scala 74:20:@35312.4]
  assign regs_76_clock = clock; // @[:@35321.4]
  assign regs_76_reset = io_reset; // @[:@35322.4 RegFile.scala 76:16:@35329.4]
  assign regs_76_io_in = 64'h0; // @[RegFile.scala 75:16:@35328.4]
  assign regs_76_io_reset = reset; // @[RegFile.scala 78:19:@35332.4]
  assign regs_76_io_enable = 1'h1; // @[RegFile.scala 74:20:@35326.4]
  assign regs_77_clock = clock; // @[:@35335.4]
  assign regs_77_reset = io_reset; // @[:@35336.4 RegFile.scala 76:16:@35343.4]
  assign regs_77_io_in = 64'h0; // @[RegFile.scala 75:16:@35342.4]
  assign regs_77_io_reset = reset; // @[RegFile.scala 78:19:@35346.4]
  assign regs_77_io_enable = 1'h1; // @[RegFile.scala 74:20:@35340.4]
  assign regs_78_clock = clock; // @[:@35349.4]
  assign regs_78_reset = io_reset; // @[:@35350.4 RegFile.scala 76:16:@35357.4]
  assign regs_78_io_in = 64'h0; // @[RegFile.scala 75:16:@35356.4]
  assign regs_78_io_reset = reset; // @[RegFile.scala 78:19:@35360.4]
  assign regs_78_io_enable = 1'h1; // @[RegFile.scala 74:20:@35354.4]
  assign regs_79_clock = clock; // @[:@35363.4]
  assign regs_79_reset = io_reset; // @[:@35364.4 RegFile.scala 76:16:@35371.4]
  assign regs_79_io_in = 64'h0; // @[RegFile.scala 75:16:@35370.4]
  assign regs_79_io_reset = reset; // @[RegFile.scala 78:19:@35374.4]
  assign regs_79_io_enable = 1'h1; // @[RegFile.scala 74:20:@35368.4]
  assign regs_80_clock = clock; // @[:@35377.4]
  assign regs_80_reset = io_reset; // @[:@35378.4 RegFile.scala 76:16:@35385.4]
  assign regs_80_io_in = 64'h0; // @[RegFile.scala 75:16:@35384.4]
  assign regs_80_io_reset = reset; // @[RegFile.scala 78:19:@35388.4]
  assign regs_80_io_enable = 1'h1; // @[RegFile.scala 74:20:@35382.4]
  assign regs_81_clock = clock; // @[:@35391.4]
  assign regs_81_reset = io_reset; // @[:@35392.4 RegFile.scala 76:16:@35399.4]
  assign regs_81_io_in = 64'h0; // @[RegFile.scala 75:16:@35398.4]
  assign regs_81_io_reset = reset; // @[RegFile.scala 78:19:@35402.4]
  assign regs_81_io_enable = 1'h1; // @[RegFile.scala 74:20:@35396.4]
  assign regs_82_clock = clock; // @[:@35405.4]
  assign regs_82_reset = io_reset; // @[:@35406.4 RegFile.scala 76:16:@35413.4]
  assign regs_82_io_in = 64'h0; // @[RegFile.scala 75:16:@35412.4]
  assign regs_82_io_reset = reset; // @[RegFile.scala 78:19:@35416.4]
  assign regs_82_io_enable = 1'h1; // @[RegFile.scala 74:20:@35410.4]
  assign regs_83_clock = clock; // @[:@35419.4]
  assign regs_83_reset = io_reset; // @[:@35420.4 RegFile.scala 76:16:@35427.4]
  assign regs_83_io_in = 64'h0; // @[RegFile.scala 75:16:@35426.4]
  assign regs_83_io_reset = reset; // @[RegFile.scala 78:19:@35430.4]
  assign regs_83_io_enable = 1'h1; // @[RegFile.scala 74:20:@35424.4]
  assign regs_84_clock = clock; // @[:@35433.4]
  assign regs_84_reset = io_reset; // @[:@35434.4 RegFile.scala 76:16:@35441.4]
  assign regs_84_io_in = 64'h0; // @[RegFile.scala 75:16:@35440.4]
  assign regs_84_io_reset = reset; // @[RegFile.scala 78:19:@35444.4]
  assign regs_84_io_enable = 1'h1; // @[RegFile.scala 74:20:@35438.4]
  assign regs_85_clock = clock; // @[:@35447.4]
  assign regs_85_reset = io_reset; // @[:@35448.4 RegFile.scala 76:16:@35455.4]
  assign regs_85_io_in = 64'h0; // @[RegFile.scala 75:16:@35454.4]
  assign regs_85_io_reset = reset; // @[RegFile.scala 78:19:@35458.4]
  assign regs_85_io_enable = 1'h1; // @[RegFile.scala 74:20:@35452.4]
  assign regs_86_clock = clock; // @[:@35461.4]
  assign regs_86_reset = io_reset; // @[:@35462.4 RegFile.scala 76:16:@35469.4]
  assign regs_86_io_in = 64'h0; // @[RegFile.scala 75:16:@35468.4]
  assign regs_86_io_reset = reset; // @[RegFile.scala 78:19:@35472.4]
  assign regs_86_io_enable = 1'h1; // @[RegFile.scala 74:20:@35466.4]
  assign regs_87_clock = clock; // @[:@35475.4]
  assign regs_87_reset = io_reset; // @[:@35476.4 RegFile.scala 76:16:@35483.4]
  assign regs_87_io_in = 64'h0; // @[RegFile.scala 75:16:@35482.4]
  assign regs_87_io_reset = reset; // @[RegFile.scala 78:19:@35486.4]
  assign regs_87_io_enable = 1'h1; // @[RegFile.scala 74:20:@35480.4]
  assign regs_88_clock = clock; // @[:@35489.4]
  assign regs_88_reset = io_reset; // @[:@35490.4 RegFile.scala 76:16:@35497.4]
  assign regs_88_io_in = 64'h0; // @[RegFile.scala 75:16:@35496.4]
  assign regs_88_io_reset = reset; // @[RegFile.scala 78:19:@35500.4]
  assign regs_88_io_enable = 1'h1; // @[RegFile.scala 74:20:@35494.4]
  assign regs_89_clock = clock; // @[:@35503.4]
  assign regs_89_reset = io_reset; // @[:@35504.4 RegFile.scala 76:16:@35511.4]
  assign regs_89_io_in = 64'h0; // @[RegFile.scala 75:16:@35510.4]
  assign regs_89_io_reset = reset; // @[RegFile.scala 78:19:@35514.4]
  assign regs_89_io_enable = 1'h1; // @[RegFile.scala 74:20:@35508.4]
  assign regs_90_clock = clock; // @[:@35517.4]
  assign regs_90_reset = io_reset; // @[:@35518.4 RegFile.scala 76:16:@35525.4]
  assign regs_90_io_in = 64'h0; // @[RegFile.scala 75:16:@35524.4]
  assign regs_90_io_reset = reset; // @[RegFile.scala 78:19:@35528.4]
  assign regs_90_io_enable = 1'h1; // @[RegFile.scala 74:20:@35522.4]
  assign regs_91_clock = clock; // @[:@35531.4]
  assign regs_91_reset = io_reset; // @[:@35532.4 RegFile.scala 76:16:@35539.4]
  assign regs_91_io_in = 64'h0; // @[RegFile.scala 75:16:@35538.4]
  assign regs_91_io_reset = reset; // @[RegFile.scala 78:19:@35542.4]
  assign regs_91_io_enable = 1'h1; // @[RegFile.scala 74:20:@35536.4]
  assign regs_92_clock = clock; // @[:@35545.4]
  assign regs_92_reset = io_reset; // @[:@35546.4 RegFile.scala 76:16:@35553.4]
  assign regs_92_io_in = 64'h0; // @[RegFile.scala 75:16:@35552.4]
  assign regs_92_io_reset = reset; // @[RegFile.scala 78:19:@35556.4]
  assign regs_92_io_enable = 1'h1; // @[RegFile.scala 74:20:@35550.4]
  assign regs_93_clock = clock; // @[:@35559.4]
  assign regs_93_reset = io_reset; // @[:@35560.4 RegFile.scala 76:16:@35567.4]
  assign regs_93_io_in = 64'h0; // @[RegFile.scala 75:16:@35566.4]
  assign regs_93_io_reset = reset; // @[RegFile.scala 78:19:@35570.4]
  assign regs_93_io_enable = 1'h1; // @[RegFile.scala 74:20:@35564.4]
  assign regs_94_clock = clock; // @[:@35573.4]
  assign regs_94_reset = io_reset; // @[:@35574.4 RegFile.scala 76:16:@35581.4]
  assign regs_94_io_in = 64'h0; // @[RegFile.scala 75:16:@35580.4]
  assign regs_94_io_reset = reset; // @[RegFile.scala 78:19:@35584.4]
  assign regs_94_io_enable = 1'h1; // @[RegFile.scala 74:20:@35578.4]
  assign regs_95_clock = clock; // @[:@35587.4]
  assign regs_95_reset = io_reset; // @[:@35588.4 RegFile.scala 76:16:@35595.4]
  assign regs_95_io_in = 64'h0; // @[RegFile.scala 75:16:@35594.4]
  assign regs_95_io_reset = reset; // @[RegFile.scala 78:19:@35598.4]
  assign regs_95_io_enable = 1'h1; // @[RegFile.scala 74:20:@35592.4]
  assign regs_96_clock = clock; // @[:@35601.4]
  assign regs_96_reset = io_reset; // @[:@35602.4 RegFile.scala 76:16:@35609.4]
  assign regs_96_io_in = 64'h0; // @[RegFile.scala 75:16:@35608.4]
  assign regs_96_io_reset = reset; // @[RegFile.scala 78:19:@35612.4]
  assign regs_96_io_enable = 1'h1; // @[RegFile.scala 74:20:@35606.4]
  assign regs_97_clock = clock; // @[:@35615.4]
  assign regs_97_reset = io_reset; // @[:@35616.4 RegFile.scala 76:16:@35623.4]
  assign regs_97_io_in = 64'h0; // @[RegFile.scala 75:16:@35622.4]
  assign regs_97_io_reset = reset; // @[RegFile.scala 78:19:@35626.4]
  assign regs_97_io_enable = 1'h1; // @[RegFile.scala 74:20:@35620.4]
  assign regs_98_clock = clock; // @[:@35629.4]
  assign regs_98_reset = io_reset; // @[:@35630.4 RegFile.scala 76:16:@35637.4]
  assign regs_98_io_in = 64'h0; // @[RegFile.scala 75:16:@35636.4]
  assign regs_98_io_reset = reset; // @[RegFile.scala 78:19:@35640.4]
  assign regs_98_io_enable = 1'h1; // @[RegFile.scala 74:20:@35634.4]
  assign regs_99_clock = clock; // @[:@35643.4]
  assign regs_99_reset = io_reset; // @[:@35644.4 RegFile.scala 76:16:@35651.4]
  assign regs_99_io_in = 64'h0; // @[RegFile.scala 75:16:@35650.4]
  assign regs_99_io_reset = reset; // @[RegFile.scala 78:19:@35654.4]
  assign regs_99_io_enable = 1'h1; // @[RegFile.scala 74:20:@35648.4]
  assign regs_100_clock = clock; // @[:@35657.4]
  assign regs_100_reset = io_reset; // @[:@35658.4 RegFile.scala 76:16:@35665.4]
  assign regs_100_io_in = 64'h0; // @[RegFile.scala 75:16:@35664.4]
  assign regs_100_io_reset = reset; // @[RegFile.scala 78:19:@35668.4]
  assign regs_100_io_enable = 1'h1; // @[RegFile.scala 74:20:@35662.4]
  assign regs_101_clock = clock; // @[:@35671.4]
  assign regs_101_reset = io_reset; // @[:@35672.4 RegFile.scala 76:16:@35679.4]
  assign regs_101_io_in = 64'h0; // @[RegFile.scala 75:16:@35678.4]
  assign regs_101_io_reset = reset; // @[RegFile.scala 78:19:@35682.4]
  assign regs_101_io_enable = 1'h1; // @[RegFile.scala 74:20:@35676.4]
  assign regs_102_clock = clock; // @[:@35685.4]
  assign regs_102_reset = io_reset; // @[:@35686.4 RegFile.scala 76:16:@35693.4]
  assign regs_102_io_in = 64'h0; // @[RegFile.scala 75:16:@35692.4]
  assign regs_102_io_reset = reset; // @[RegFile.scala 78:19:@35696.4]
  assign regs_102_io_enable = 1'h1; // @[RegFile.scala 74:20:@35690.4]
  assign regs_103_clock = clock; // @[:@35699.4]
  assign regs_103_reset = io_reset; // @[:@35700.4 RegFile.scala 76:16:@35707.4]
  assign regs_103_io_in = 64'h0; // @[RegFile.scala 75:16:@35706.4]
  assign regs_103_io_reset = reset; // @[RegFile.scala 78:19:@35710.4]
  assign regs_103_io_enable = 1'h1; // @[RegFile.scala 74:20:@35704.4]
  assign regs_104_clock = clock; // @[:@35713.4]
  assign regs_104_reset = io_reset; // @[:@35714.4 RegFile.scala 76:16:@35721.4]
  assign regs_104_io_in = 64'h0; // @[RegFile.scala 75:16:@35720.4]
  assign regs_104_io_reset = reset; // @[RegFile.scala 78:19:@35724.4]
  assign regs_104_io_enable = 1'h1; // @[RegFile.scala 74:20:@35718.4]
  assign regs_105_clock = clock; // @[:@35727.4]
  assign regs_105_reset = io_reset; // @[:@35728.4 RegFile.scala 76:16:@35735.4]
  assign regs_105_io_in = 64'h0; // @[RegFile.scala 75:16:@35734.4]
  assign regs_105_io_reset = reset; // @[RegFile.scala 78:19:@35738.4]
  assign regs_105_io_enable = 1'h1; // @[RegFile.scala 74:20:@35732.4]
  assign regs_106_clock = clock; // @[:@35741.4]
  assign regs_106_reset = io_reset; // @[:@35742.4 RegFile.scala 76:16:@35749.4]
  assign regs_106_io_in = 64'h0; // @[RegFile.scala 75:16:@35748.4]
  assign regs_106_io_reset = reset; // @[RegFile.scala 78:19:@35752.4]
  assign regs_106_io_enable = 1'h1; // @[RegFile.scala 74:20:@35746.4]
  assign regs_107_clock = clock; // @[:@35755.4]
  assign regs_107_reset = io_reset; // @[:@35756.4 RegFile.scala 76:16:@35763.4]
  assign regs_107_io_in = 64'h0; // @[RegFile.scala 75:16:@35762.4]
  assign regs_107_io_reset = reset; // @[RegFile.scala 78:19:@35766.4]
  assign regs_107_io_enable = 1'h1; // @[RegFile.scala 74:20:@35760.4]
  assign regs_108_clock = clock; // @[:@35769.4]
  assign regs_108_reset = io_reset; // @[:@35770.4 RegFile.scala 76:16:@35777.4]
  assign regs_108_io_in = 64'h0; // @[RegFile.scala 75:16:@35776.4]
  assign regs_108_io_reset = reset; // @[RegFile.scala 78:19:@35780.4]
  assign regs_108_io_enable = 1'h1; // @[RegFile.scala 74:20:@35774.4]
  assign regs_109_clock = clock; // @[:@35783.4]
  assign regs_109_reset = io_reset; // @[:@35784.4 RegFile.scala 76:16:@35791.4]
  assign regs_109_io_in = 64'h0; // @[RegFile.scala 75:16:@35790.4]
  assign regs_109_io_reset = reset; // @[RegFile.scala 78:19:@35794.4]
  assign regs_109_io_enable = 1'h1; // @[RegFile.scala 74:20:@35788.4]
  assign regs_110_clock = clock; // @[:@35797.4]
  assign regs_110_reset = io_reset; // @[:@35798.4 RegFile.scala 76:16:@35805.4]
  assign regs_110_io_in = 64'h0; // @[RegFile.scala 75:16:@35804.4]
  assign regs_110_io_reset = reset; // @[RegFile.scala 78:19:@35808.4]
  assign regs_110_io_enable = 1'h1; // @[RegFile.scala 74:20:@35802.4]
  assign regs_111_clock = clock; // @[:@35811.4]
  assign regs_111_reset = io_reset; // @[:@35812.4 RegFile.scala 76:16:@35819.4]
  assign regs_111_io_in = 64'h0; // @[RegFile.scala 75:16:@35818.4]
  assign regs_111_io_reset = reset; // @[RegFile.scala 78:19:@35822.4]
  assign regs_111_io_enable = 1'h1; // @[RegFile.scala 74:20:@35816.4]
  assign regs_112_clock = clock; // @[:@35825.4]
  assign regs_112_reset = io_reset; // @[:@35826.4 RegFile.scala 76:16:@35833.4]
  assign regs_112_io_in = 64'h0; // @[RegFile.scala 75:16:@35832.4]
  assign regs_112_io_reset = reset; // @[RegFile.scala 78:19:@35836.4]
  assign regs_112_io_enable = 1'h1; // @[RegFile.scala 74:20:@35830.4]
  assign regs_113_clock = clock; // @[:@35839.4]
  assign regs_113_reset = io_reset; // @[:@35840.4 RegFile.scala 76:16:@35847.4]
  assign regs_113_io_in = 64'h0; // @[RegFile.scala 75:16:@35846.4]
  assign regs_113_io_reset = reset; // @[RegFile.scala 78:19:@35850.4]
  assign regs_113_io_enable = 1'h1; // @[RegFile.scala 74:20:@35844.4]
  assign regs_114_clock = clock; // @[:@35853.4]
  assign regs_114_reset = io_reset; // @[:@35854.4 RegFile.scala 76:16:@35861.4]
  assign regs_114_io_in = 64'h0; // @[RegFile.scala 75:16:@35860.4]
  assign regs_114_io_reset = reset; // @[RegFile.scala 78:19:@35864.4]
  assign regs_114_io_enable = 1'h1; // @[RegFile.scala 74:20:@35858.4]
  assign regs_115_clock = clock; // @[:@35867.4]
  assign regs_115_reset = io_reset; // @[:@35868.4 RegFile.scala 76:16:@35875.4]
  assign regs_115_io_in = 64'h0; // @[RegFile.scala 75:16:@35874.4]
  assign regs_115_io_reset = reset; // @[RegFile.scala 78:19:@35878.4]
  assign regs_115_io_enable = 1'h1; // @[RegFile.scala 74:20:@35872.4]
  assign regs_116_clock = clock; // @[:@35881.4]
  assign regs_116_reset = io_reset; // @[:@35882.4 RegFile.scala 76:16:@35889.4]
  assign regs_116_io_in = 64'h0; // @[RegFile.scala 75:16:@35888.4]
  assign regs_116_io_reset = reset; // @[RegFile.scala 78:19:@35892.4]
  assign regs_116_io_enable = 1'h1; // @[RegFile.scala 74:20:@35886.4]
  assign regs_117_clock = clock; // @[:@35895.4]
  assign regs_117_reset = io_reset; // @[:@35896.4 RegFile.scala 76:16:@35903.4]
  assign regs_117_io_in = 64'h0; // @[RegFile.scala 75:16:@35902.4]
  assign regs_117_io_reset = reset; // @[RegFile.scala 78:19:@35906.4]
  assign regs_117_io_enable = 1'h1; // @[RegFile.scala 74:20:@35900.4]
  assign regs_118_clock = clock; // @[:@35909.4]
  assign regs_118_reset = io_reset; // @[:@35910.4 RegFile.scala 76:16:@35917.4]
  assign regs_118_io_in = 64'h0; // @[RegFile.scala 75:16:@35916.4]
  assign regs_118_io_reset = reset; // @[RegFile.scala 78:19:@35920.4]
  assign regs_118_io_enable = 1'h1; // @[RegFile.scala 74:20:@35914.4]
  assign regs_119_clock = clock; // @[:@35923.4]
  assign regs_119_reset = io_reset; // @[:@35924.4 RegFile.scala 76:16:@35931.4]
  assign regs_119_io_in = 64'h0; // @[RegFile.scala 75:16:@35930.4]
  assign regs_119_io_reset = reset; // @[RegFile.scala 78:19:@35934.4]
  assign regs_119_io_enable = 1'h1; // @[RegFile.scala 74:20:@35928.4]
  assign regs_120_clock = clock; // @[:@35937.4]
  assign regs_120_reset = io_reset; // @[:@35938.4 RegFile.scala 76:16:@35945.4]
  assign regs_120_io_in = 64'h0; // @[RegFile.scala 75:16:@35944.4]
  assign regs_120_io_reset = reset; // @[RegFile.scala 78:19:@35948.4]
  assign regs_120_io_enable = 1'h1; // @[RegFile.scala 74:20:@35942.4]
  assign regs_121_clock = clock; // @[:@35951.4]
  assign regs_121_reset = io_reset; // @[:@35952.4 RegFile.scala 76:16:@35959.4]
  assign regs_121_io_in = 64'h0; // @[RegFile.scala 75:16:@35958.4]
  assign regs_121_io_reset = reset; // @[RegFile.scala 78:19:@35962.4]
  assign regs_121_io_enable = 1'h1; // @[RegFile.scala 74:20:@35956.4]
  assign regs_122_clock = clock; // @[:@35965.4]
  assign regs_122_reset = io_reset; // @[:@35966.4 RegFile.scala 76:16:@35973.4]
  assign regs_122_io_in = 64'h0; // @[RegFile.scala 75:16:@35972.4]
  assign regs_122_io_reset = reset; // @[RegFile.scala 78:19:@35976.4]
  assign regs_122_io_enable = 1'h1; // @[RegFile.scala 74:20:@35970.4]
  assign regs_123_clock = clock; // @[:@35979.4]
  assign regs_123_reset = io_reset; // @[:@35980.4 RegFile.scala 76:16:@35987.4]
  assign regs_123_io_in = 64'h0; // @[RegFile.scala 75:16:@35986.4]
  assign regs_123_io_reset = reset; // @[RegFile.scala 78:19:@35990.4]
  assign regs_123_io_enable = 1'h1; // @[RegFile.scala 74:20:@35984.4]
  assign regs_124_clock = clock; // @[:@35993.4]
  assign regs_124_reset = io_reset; // @[:@35994.4 RegFile.scala 76:16:@36001.4]
  assign regs_124_io_in = 64'h0; // @[RegFile.scala 75:16:@36000.4]
  assign regs_124_io_reset = reset; // @[RegFile.scala 78:19:@36004.4]
  assign regs_124_io_enable = 1'h1; // @[RegFile.scala 74:20:@35998.4]
  assign regs_125_clock = clock; // @[:@36007.4]
  assign regs_125_reset = io_reset; // @[:@36008.4 RegFile.scala 76:16:@36015.4]
  assign regs_125_io_in = 64'h0; // @[RegFile.scala 75:16:@36014.4]
  assign regs_125_io_reset = reset; // @[RegFile.scala 78:19:@36018.4]
  assign regs_125_io_enable = 1'h1; // @[RegFile.scala 74:20:@36012.4]
  assign regs_126_clock = clock; // @[:@36021.4]
  assign regs_126_reset = io_reset; // @[:@36022.4 RegFile.scala 76:16:@36029.4]
  assign regs_126_io_in = 64'h0; // @[RegFile.scala 75:16:@36028.4]
  assign regs_126_io_reset = reset; // @[RegFile.scala 78:19:@36032.4]
  assign regs_126_io_enable = 1'h1; // @[RegFile.scala 74:20:@36026.4]
  assign regs_127_clock = clock; // @[:@36035.4]
  assign regs_127_reset = io_reset; // @[:@36036.4 RegFile.scala 76:16:@36043.4]
  assign regs_127_io_in = 64'h0; // @[RegFile.scala 75:16:@36042.4]
  assign regs_127_io_reset = reset; // @[RegFile.scala 78:19:@36046.4]
  assign regs_127_io_enable = 1'h1; // @[RegFile.scala 74:20:@36040.4]
  assign regs_128_clock = clock; // @[:@36049.4]
  assign regs_128_reset = io_reset; // @[:@36050.4 RegFile.scala 76:16:@36057.4]
  assign regs_128_io_in = 64'h0; // @[RegFile.scala 75:16:@36056.4]
  assign regs_128_io_reset = reset; // @[RegFile.scala 78:19:@36060.4]
  assign regs_128_io_enable = 1'h1; // @[RegFile.scala 74:20:@36054.4]
  assign regs_129_clock = clock; // @[:@36063.4]
  assign regs_129_reset = io_reset; // @[:@36064.4 RegFile.scala 76:16:@36071.4]
  assign regs_129_io_in = 64'h0; // @[RegFile.scala 75:16:@36070.4]
  assign regs_129_io_reset = reset; // @[RegFile.scala 78:19:@36074.4]
  assign regs_129_io_enable = 1'h1; // @[RegFile.scala 74:20:@36068.4]
  assign regs_130_clock = clock; // @[:@36077.4]
  assign regs_130_reset = io_reset; // @[:@36078.4 RegFile.scala 76:16:@36085.4]
  assign regs_130_io_in = 64'h0; // @[RegFile.scala 75:16:@36084.4]
  assign regs_130_io_reset = reset; // @[RegFile.scala 78:19:@36088.4]
  assign regs_130_io_enable = 1'h1; // @[RegFile.scala 74:20:@36082.4]
  assign regs_131_clock = clock; // @[:@36091.4]
  assign regs_131_reset = io_reset; // @[:@36092.4 RegFile.scala 76:16:@36099.4]
  assign regs_131_io_in = 64'h0; // @[RegFile.scala 75:16:@36098.4]
  assign regs_131_io_reset = reset; // @[RegFile.scala 78:19:@36102.4]
  assign regs_131_io_enable = 1'h1; // @[RegFile.scala 74:20:@36096.4]
  assign regs_132_clock = clock; // @[:@36105.4]
  assign regs_132_reset = io_reset; // @[:@36106.4 RegFile.scala 76:16:@36113.4]
  assign regs_132_io_in = 64'h0; // @[RegFile.scala 75:16:@36112.4]
  assign regs_132_io_reset = reset; // @[RegFile.scala 78:19:@36116.4]
  assign regs_132_io_enable = 1'h1; // @[RegFile.scala 74:20:@36110.4]
  assign regs_133_clock = clock; // @[:@36119.4]
  assign regs_133_reset = io_reset; // @[:@36120.4 RegFile.scala 76:16:@36127.4]
  assign regs_133_io_in = 64'h0; // @[RegFile.scala 75:16:@36126.4]
  assign regs_133_io_reset = reset; // @[RegFile.scala 78:19:@36130.4]
  assign regs_133_io_enable = 1'h1; // @[RegFile.scala 74:20:@36124.4]
  assign regs_134_clock = clock; // @[:@36133.4]
  assign regs_134_reset = io_reset; // @[:@36134.4 RegFile.scala 76:16:@36141.4]
  assign regs_134_io_in = 64'h0; // @[RegFile.scala 75:16:@36140.4]
  assign regs_134_io_reset = reset; // @[RegFile.scala 78:19:@36144.4]
  assign regs_134_io_enable = 1'h1; // @[RegFile.scala 74:20:@36138.4]
  assign regs_135_clock = clock; // @[:@36147.4]
  assign regs_135_reset = io_reset; // @[:@36148.4 RegFile.scala 76:16:@36155.4]
  assign regs_135_io_in = 64'h0; // @[RegFile.scala 75:16:@36154.4]
  assign regs_135_io_reset = reset; // @[RegFile.scala 78:19:@36158.4]
  assign regs_135_io_enable = 1'h1; // @[RegFile.scala 74:20:@36152.4]
  assign regs_136_clock = clock; // @[:@36161.4]
  assign regs_136_reset = io_reset; // @[:@36162.4 RegFile.scala 76:16:@36169.4]
  assign regs_136_io_in = 64'h0; // @[RegFile.scala 75:16:@36168.4]
  assign regs_136_io_reset = reset; // @[RegFile.scala 78:19:@36172.4]
  assign regs_136_io_enable = 1'h1; // @[RegFile.scala 74:20:@36166.4]
  assign regs_137_clock = clock; // @[:@36175.4]
  assign regs_137_reset = io_reset; // @[:@36176.4 RegFile.scala 76:16:@36183.4]
  assign regs_137_io_in = 64'h0; // @[RegFile.scala 75:16:@36182.4]
  assign regs_137_io_reset = reset; // @[RegFile.scala 78:19:@36186.4]
  assign regs_137_io_enable = 1'h1; // @[RegFile.scala 74:20:@36180.4]
  assign regs_138_clock = clock; // @[:@36189.4]
  assign regs_138_reset = io_reset; // @[:@36190.4 RegFile.scala 76:16:@36197.4]
  assign regs_138_io_in = 64'h0; // @[RegFile.scala 75:16:@36196.4]
  assign regs_138_io_reset = reset; // @[RegFile.scala 78:19:@36200.4]
  assign regs_138_io_enable = 1'h1; // @[RegFile.scala 74:20:@36194.4]
  assign regs_139_clock = clock; // @[:@36203.4]
  assign regs_139_reset = io_reset; // @[:@36204.4 RegFile.scala 76:16:@36211.4]
  assign regs_139_io_in = 64'h0; // @[RegFile.scala 75:16:@36210.4]
  assign regs_139_io_reset = reset; // @[RegFile.scala 78:19:@36214.4]
  assign regs_139_io_enable = 1'h1; // @[RegFile.scala 74:20:@36208.4]
  assign regs_140_clock = clock; // @[:@36217.4]
  assign regs_140_reset = io_reset; // @[:@36218.4 RegFile.scala 76:16:@36225.4]
  assign regs_140_io_in = 64'h0; // @[RegFile.scala 75:16:@36224.4]
  assign regs_140_io_reset = reset; // @[RegFile.scala 78:19:@36228.4]
  assign regs_140_io_enable = 1'h1; // @[RegFile.scala 74:20:@36222.4]
  assign regs_141_clock = clock; // @[:@36231.4]
  assign regs_141_reset = io_reset; // @[:@36232.4 RegFile.scala 76:16:@36239.4]
  assign regs_141_io_in = 64'h0; // @[RegFile.scala 75:16:@36238.4]
  assign regs_141_io_reset = reset; // @[RegFile.scala 78:19:@36242.4]
  assign regs_141_io_enable = 1'h1; // @[RegFile.scala 74:20:@36236.4]
  assign regs_142_clock = clock; // @[:@36245.4]
  assign regs_142_reset = io_reset; // @[:@36246.4 RegFile.scala 76:16:@36253.4]
  assign regs_142_io_in = 64'h0; // @[RegFile.scala 75:16:@36252.4]
  assign regs_142_io_reset = reset; // @[RegFile.scala 78:19:@36256.4]
  assign regs_142_io_enable = 1'h1; // @[RegFile.scala 74:20:@36250.4]
  assign regs_143_clock = clock; // @[:@36259.4]
  assign regs_143_reset = io_reset; // @[:@36260.4 RegFile.scala 76:16:@36267.4]
  assign regs_143_io_in = 64'h0; // @[RegFile.scala 75:16:@36266.4]
  assign regs_143_io_reset = reset; // @[RegFile.scala 78:19:@36270.4]
  assign regs_143_io_enable = 1'h1; // @[RegFile.scala 74:20:@36264.4]
  assign regs_144_clock = clock; // @[:@36273.4]
  assign regs_144_reset = io_reset; // @[:@36274.4 RegFile.scala 76:16:@36281.4]
  assign regs_144_io_in = 64'h0; // @[RegFile.scala 75:16:@36280.4]
  assign regs_144_io_reset = reset; // @[RegFile.scala 78:19:@36284.4]
  assign regs_144_io_enable = 1'h1; // @[RegFile.scala 74:20:@36278.4]
  assign regs_145_clock = clock; // @[:@36287.4]
  assign regs_145_reset = io_reset; // @[:@36288.4 RegFile.scala 76:16:@36295.4]
  assign regs_145_io_in = 64'h0; // @[RegFile.scala 75:16:@36294.4]
  assign regs_145_io_reset = reset; // @[RegFile.scala 78:19:@36298.4]
  assign regs_145_io_enable = 1'h1; // @[RegFile.scala 74:20:@36292.4]
  assign regs_146_clock = clock; // @[:@36301.4]
  assign regs_146_reset = io_reset; // @[:@36302.4 RegFile.scala 76:16:@36309.4]
  assign regs_146_io_in = 64'h0; // @[RegFile.scala 75:16:@36308.4]
  assign regs_146_io_reset = reset; // @[RegFile.scala 78:19:@36312.4]
  assign regs_146_io_enable = 1'h1; // @[RegFile.scala 74:20:@36306.4]
  assign regs_147_clock = clock; // @[:@36315.4]
  assign regs_147_reset = io_reset; // @[:@36316.4 RegFile.scala 76:16:@36323.4]
  assign regs_147_io_in = 64'h0; // @[RegFile.scala 75:16:@36322.4]
  assign regs_147_io_reset = reset; // @[RegFile.scala 78:19:@36326.4]
  assign regs_147_io_enable = 1'h1; // @[RegFile.scala 74:20:@36320.4]
  assign regs_148_clock = clock; // @[:@36329.4]
  assign regs_148_reset = io_reset; // @[:@36330.4 RegFile.scala 76:16:@36337.4]
  assign regs_148_io_in = 64'h0; // @[RegFile.scala 75:16:@36336.4]
  assign regs_148_io_reset = reset; // @[RegFile.scala 78:19:@36340.4]
  assign regs_148_io_enable = 1'h1; // @[RegFile.scala 74:20:@36334.4]
  assign regs_149_clock = clock; // @[:@36343.4]
  assign regs_149_reset = io_reset; // @[:@36344.4 RegFile.scala 76:16:@36351.4]
  assign regs_149_io_in = 64'h0; // @[RegFile.scala 75:16:@36350.4]
  assign regs_149_io_reset = reset; // @[RegFile.scala 78:19:@36354.4]
  assign regs_149_io_enable = 1'h1; // @[RegFile.scala 74:20:@36348.4]
  assign regs_150_clock = clock; // @[:@36357.4]
  assign regs_150_reset = io_reset; // @[:@36358.4 RegFile.scala 76:16:@36365.4]
  assign regs_150_io_in = 64'h0; // @[RegFile.scala 75:16:@36364.4]
  assign regs_150_io_reset = reset; // @[RegFile.scala 78:19:@36368.4]
  assign regs_150_io_enable = 1'h1; // @[RegFile.scala 74:20:@36362.4]
  assign regs_151_clock = clock; // @[:@36371.4]
  assign regs_151_reset = io_reset; // @[:@36372.4 RegFile.scala 76:16:@36379.4]
  assign regs_151_io_in = 64'h0; // @[RegFile.scala 75:16:@36378.4]
  assign regs_151_io_reset = reset; // @[RegFile.scala 78:19:@36382.4]
  assign regs_151_io_enable = 1'h1; // @[RegFile.scala 74:20:@36376.4]
  assign regs_152_clock = clock; // @[:@36385.4]
  assign regs_152_reset = io_reset; // @[:@36386.4 RegFile.scala 76:16:@36393.4]
  assign regs_152_io_in = 64'h0; // @[RegFile.scala 75:16:@36392.4]
  assign regs_152_io_reset = reset; // @[RegFile.scala 78:19:@36396.4]
  assign regs_152_io_enable = 1'h1; // @[RegFile.scala 74:20:@36390.4]
  assign regs_153_clock = clock; // @[:@36399.4]
  assign regs_153_reset = io_reset; // @[:@36400.4 RegFile.scala 76:16:@36407.4]
  assign regs_153_io_in = 64'h0; // @[RegFile.scala 75:16:@36406.4]
  assign regs_153_io_reset = reset; // @[RegFile.scala 78:19:@36410.4]
  assign regs_153_io_enable = 1'h1; // @[RegFile.scala 74:20:@36404.4]
  assign regs_154_clock = clock; // @[:@36413.4]
  assign regs_154_reset = io_reset; // @[:@36414.4 RegFile.scala 76:16:@36421.4]
  assign regs_154_io_in = 64'h0; // @[RegFile.scala 75:16:@36420.4]
  assign regs_154_io_reset = reset; // @[RegFile.scala 78:19:@36424.4]
  assign regs_154_io_enable = 1'h1; // @[RegFile.scala 74:20:@36418.4]
  assign regs_155_clock = clock; // @[:@36427.4]
  assign regs_155_reset = io_reset; // @[:@36428.4 RegFile.scala 76:16:@36435.4]
  assign regs_155_io_in = 64'h0; // @[RegFile.scala 75:16:@36434.4]
  assign regs_155_io_reset = reset; // @[RegFile.scala 78:19:@36438.4]
  assign regs_155_io_enable = 1'h1; // @[RegFile.scala 74:20:@36432.4]
  assign regs_156_clock = clock; // @[:@36441.4]
  assign regs_156_reset = io_reset; // @[:@36442.4 RegFile.scala 76:16:@36449.4]
  assign regs_156_io_in = 64'h0; // @[RegFile.scala 75:16:@36448.4]
  assign regs_156_io_reset = reset; // @[RegFile.scala 78:19:@36452.4]
  assign regs_156_io_enable = 1'h1; // @[RegFile.scala 74:20:@36446.4]
  assign regs_157_clock = clock; // @[:@36455.4]
  assign regs_157_reset = io_reset; // @[:@36456.4 RegFile.scala 76:16:@36463.4]
  assign regs_157_io_in = 64'h0; // @[RegFile.scala 75:16:@36462.4]
  assign regs_157_io_reset = reset; // @[RegFile.scala 78:19:@36466.4]
  assign regs_157_io_enable = 1'h1; // @[RegFile.scala 74:20:@36460.4]
  assign regs_158_clock = clock; // @[:@36469.4]
  assign regs_158_reset = io_reset; // @[:@36470.4 RegFile.scala 76:16:@36477.4]
  assign regs_158_io_in = 64'h0; // @[RegFile.scala 75:16:@36476.4]
  assign regs_158_io_reset = reset; // @[RegFile.scala 78:19:@36480.4]
  assign regs_158_io_enable = 1'h1; // @[RegFile.scala 74:20:@36474.4]
  assign regs_159_clock = clock; // @[:@36483.4]
  assign regs_159_reset = io_reset; // @[:@36484.4 RegFile.scala 76:16:@36491.4]
  assign regs_159_io_in = 64'h0; // @[RegFile.scala 75:16:@36490.4]
  assign regs_159_io_reset = reset; // @[RegFile.scala 78:19:@36494.4]
  assign regs_159_io_enable = 1'h1; // @[RegFile.scala 74:20:@36488.4]
  assign regs_160_clock = clock; // @[:@36497.4]
  assign regs_160_reset = io_reset; // @[:@36498.4 RegFile.scala 76:16:@36505.4]
  assign regs_160_io_in = 64'h0; // @[RegFile.scala 75:16:@36504.4]
  assign regs_160_io_reset = reset; // @[RegFile.scala 78:19:@36508.4]
  assign regs_160_io_enable = 1'h1; // @[RegFile.scala 74:20:@36502.4]
  assign regs_161_clock = clock; // @[:@36511.4]
  assign regs_161_reset = io_reset; // @[:@36512.4 RegFile.scala 76:16:@36519.4]
  assign regs_161_io_in = 64'h0; // @[RegFile.scala 75:16:@36518.4]
  assign regs_161_io_reset = reset; // @[RegFile.scala 78:19:@36522.4]
  assign regs_161_io_enable = 1'h1; // @[RegFile.scala 74:20:@36516.4]
  assign regs_162_clock = clock; // @[:@36525.4]
  assign regs_162_reset = io_reset; // @[:@36526.4 RegFile.scala 76:16:@36533.4]
  assign regs_162_io_in = 64'h0; // @[RegFile.scala 75:16:@36532.4]
  assign regs_162_io_reset = reset; // @[RegFile.scala 78:19:@36536.4]
  assign regs_162_io_enable = 1'h1; // @[RegFile.scala 74:20:@36530.4]
  assign regs_163_clock = clock; // @[:@36539.4]
  assign regs_163_reset = io_reset; // @[:@36540.4 RegFile.scala 76:16:@36547.4]
  assign regs_163_io_in = 64'h0; // @[RegFile.scala 75:16:@36546.4]
  assign regs_163_io_reset = reset; // @[RegFile.scala 78:19:@36550.4]
  assign regs_163_io_enable = 1'h1; // @[RegFile.scala 74:20:@36544.4]
  assign regs_164_clock = clock; // @[:@36553.4]
  assign regs_164_reset = io_reset; // @[:@36554.4 RegFile.scala 76:16:@36561.4]
  assign regs_164_io_in = 64'h0; // @[RegFile.scala 75:16:@36560.4]
  assign regs_164_io_reset = reset; // @[RegFile.scala 78:19:@36564.4]
  assign regs_164_io_enable = 1'h1; // @[RegFile.scala 74:20:@36558.4]
  assign regs_165_clock = clock; // @[:@36567.4]
  assign regs_165_reset = io_reset; // @[:@36568.4 RegFile.scala 76:16:@36575.4]
  assign regs_165_io_in = 64'h0; // @[RegFile.scala 75:16:@36574.4]
  assign regs_165_io_reset = reset; // @[RegFile.scala 78:19:@36578.4]
  assign regs_165_io_enable = 1'h1; // @[RegFile.scala 74:20:@36572.4]
  assign regs_166_clock = clock; // @[:@36581.4]
  assign regs_166_reset = io_reset; // @[:@36582.4 RegFile.scala 76:16:@36589.4]
  assign regs_166_io_in = 64'h0; // @[RegFile.scala 75:16:@36588.4]
  assign regs_166_io_reset = reset; // @[RegFile.scala 78:19:@36592.4]
  assign regs_166_io_enable = 1'h1; // @[RegFile.scala 74:20:@36586.4]
  assign regs_167_clock = clock; // @[:@36595.4]
  assign regs_167_reset = io_reset; // @[:@36596.4 RegFile.scala 76:16:@36603.4]
  assign regs_167_io_in = 64'h0; // @[RegFile.scala 75:16:@36602.4]
  assign regs_167_io_reset = reset; // @[RegFile.scala 78:19:@36606.4]
  assign regs_167_io_enable = 1'h1; // @[RegFile.scala 74:20:@36600.4]
  assign regs_168_clock = clock; // @[:@36609.4]
  assign regs_168_reset = io_reset; // @[:@36610.4 RegFile.scala 76:16:@36617.4]
  assign regs_168_io_in = 64'h0; // @[RegFile.scala 75:16:@36616.4]
  assign regs_168_io_reset = reset; // @[RegFile.scala 78:19:@36620.4]
  assign regs_168_io_enable = 1'h1; // @[RegFile.scala 74:20:@36614.4]
  assign regs_169_clock = clock; // @[:@36623.4]
  assign regs_169_reset = io_reset; // @[:@36624.4 RegFile.scala 76:16:@36631.4]
  assign regs_169_io_in = 64'h0; // @[RegFile.scala 75:16:@36630.4]
  assign regs_169_io_reset = reset; // @[RegFile.scala 78:19:@36634.4]
  assign regs_169_io_enable = 1'h1; // @[RegFile.scala 74:20:@36628.4]
  assign regs_170_clock = clock; // @[:@36637.4]
  assign regs_170_reset = io_reset; // @[:@36638.4 RegFile.scala 76:16:@36645.4]
  assign regs_170_io_in = 64'h0; // @[RegFile.scala 75:16:@36644.4]
  assign regs_170_io_reset = reset; // @[RegFile.scala 78:19:@36648.4]
  assign regs_170_io_enable = 1'h1; // @[RegFile.scala 74:20:@36642.4]
  assign regs_171_clock = clock; // @[:@36651.4]
  assign regs_171_reset = io_reset; // @[:@36652.4 RegFile.scala 76:16:@36659.4]
  assign regs_171_io_in = 64'h0; // @[RegFile.scala 75:16:@36658.4]
  assign regs_171_io_reset = reset; // @[RegFile.scala 78:19:@36662.4]
  assign regs_171_io_enable = 1'h1; // @[RegFile.scala 74:20:@36656.4]
  assign regs_172_clock = clock; // @[:@36665.4]
  assign regs_172_reset = io_reset; // @[:@36666.4 RegFile.scala 76:16:@36673.4]
  assign regs_172_io_in = 64'h0; // @[RegFile.scala 75:16:@36672.4]
  assign regs_172_io_reset = reset; // @[RegFile.scala 78:19:@36676.4]
  assign regs_172_io_enable = 1'h1; // @[RegFile.scala 74:20:@36670.4]
  assign regs_173_clock = clock; // @[:@36679.4]
  assign regs_173_reset = io_reset; // @[:@36680.4 RegFile.scala 76:16:@36687.4]
  assign regs_173_io_in = 64'h0; // @[RegFile.scala 75:16:@36686.4]
  assign regs_173_io_reset = reset; // @[RegFile.scala 78:19:@36690.4]
  assign regs_173_io_enable = 1'h1; // @[RegFile.scala 74:20:@36684.4]
  assign regs_174_clock = clock; // @[:@36693.4]
  assign regs_174_reset = io_reset; // @[:@36694.4 RegFile.scala 76:16:@36701.4]
  assign regs_174_io_in = 64'h0; // @[RegFile.scala 75:16:@36700.4]
  assign regs_174_io_reset = reset; // @[RegFile.scala 78:19:@36704.4]
  assign regs_174_io_enable = 1'h1; // @[RegFile.scala 74:20:@36698.4]
  assign regs_175_clock = clock; // @[:@36707.4]
  assign regs_175_reset = io_reset; // @[:@36708.4 RegFile.scala 76:16:@36715.4]
  assign regs_175_io_in = 64'h0; // @[RegFile.scala 75:16:@36714.4]
  assign regs_175_io_reset = reset; // @[RegFile.scala 78:19:@36718.4]
  assign regs_175_io_enable = 1'h1; // @[RegFile.scala 74:20:@36712.4]
  assign regs_176_clock = clock; // @[:@36721.4]
  assign regs_176_reset = io_reset; // @[:@36722.4 RegFile.scala 76:16:@36729.4]
  assign regs_176_io_in = 64'h0; // @[RegFile.scala 75:16:@36728.4]
  assign regs_176_io_reset = reset; // @[RegFile.scala 78:19:@36732.4]
  assign regs_176_io_enable = 1'h1; // @[RegFile.scala 74:20:@36726.4]
  assign regs_177_clock = clock; // @[:@36735.4]
  assign regs_177_reset = io_reset; // @[:@36736.4 RegFile.scala 76:16:@36743.4]
  assign regs_177_io_in = 64'h0; // @[RegFile.scala 75:16:@36742.4]
  assign regs_177_io_reset = reset; // @[RegFile.scala 78:19:@36746.4]
  assign regs_177_io_enable = 1'h1; // @[RegFile.scala 74:20:@36740.4]
  assign regs_178_clock = clock; // @[:@36749.4]
  assign regs_178_reset = io_reset; // @[:@36750.4 RegFile.scala 76:16:@36757.4]
  assign regs_178_io_in = 64'h0; // @[RegFile.scala 75:16:@36756.4]
  assign regs_178_io_reset = reset; // @[RegFile.scala 78:19:@36760.4]
  assign regs_178_io_enable = 1'h1; // @[RegFile.scala 74:20:@36754.4]
  assign regs_179_clock = clock; // @[:@36763.4]
  assign regs_179_reset = io_reset; // @[:@36764.4 RegFile.scala 76:16:@36771.4]
  assign regs_179_io_in = 64'h0; // @[RegFile.scala 75:16:@36770.4]
  assign regs_179_io_reset = reset; // @[RegFile.scala 78:19:@36774.4]
  assign regs_179_io_enable = 1'h1; // @[RegFile.scala 74:20:@36768.4]
  assign regs_180_clock = clock; // @[:@36777.4]
  assign regs_180_reset = io_reset; // @[:@36778.4 RegFile.scala 76:16:@36785.4]
  assign regs_180_io_in = 64'h0; // @[RegFile.scala 75:16:@36784.4]
  assign regs_180_io_reset = reset; // @[RegFile.scala 78:19:@36788.4]
  assign regs_180_io_enable = 1'h1; // @[RegFile.scala 74:20:@36782.4]
  assign regs_181_clock = clock; // @[:@36791.4]
  assign regs_181_reset = io_reset; // @[:@36792.4 RegFile.scala 76:16:@36799.4]
  assign regs_181_io_in = 64'h0; // @[RegFile.scala 75:16:@36798.4]
  assign regs_181_io_reset = reset; // @[RegFile.scala 78:19:@36802.4]
  assign regs_181_io_enable = 1'h1; // @[RegFile.scala 74:20:@36796.4]
  assign regs_182_clock = clock; // @[:@36805.4]
  assign regs_182_reset = io_reset; // @[:@36806.4 RegFile.scala 76:16:@36813.4]
  assign regs_182_io_in = 64'h0; // @[RegFile.scala 75:16:@36812.4]
  assign regs_182_io_reset = reset; // @[RegFile.scala 78:19:@36816.4]
  assign regs_182_io_enable = 1'h1; // @[RegFile.scala 74:20:@36810.4]
  assign regs_183_clock = clock; // @[:@36819.4]
  assign regs_183_reset = io_reset; // @[:@36820.4 RegFile.scala 76:16:@36827.4]
  assign regs_183_io_in = 64'h0; // @[RegFile.scala 75:16:@36826.4]
  assign regs_183_io_reset = reset; // @[RegFile.scala 78:19:@36830.4]
  assign regs_183_io_enable = 1'h1; // @[RegFile.scala 74:20:@36824.4]
  assign regs_184_clock = clock; // @[:@36833.4]
  assign regs_184_reset = io_reset; // @[:@36834.4 RegFile.scala 76:16:@36841.4]
  assign regs_184_io_in = 64'h0; // @[RegFile.scala 75:16:@36840.4]
  assign regs_184_io_reset = reset; // @[RegFile.scala 78:19:@36844.4]
  assign regs_184_io_enable = 1'h1; // @[RegFile.scala 74:20:@36838.4]
  assign regs_185_clock = clock; // @[:@36847.4]
  assign regs_185_reset = io_reset; // @[:@36848.4 RegFile.scala 76:16:@36855.4]
  assign regs_185_io_in = 64'h0; // @[RegFile.scala 75:16:@36854.4]
  assign regs_185_io_reset = reset; // @[RegFile.scala 78:19:@36858.4]
  assign regs_185_io_enable = 1'h1; // @[RegFile.scala 74:20:@36852.4]
  assign regs_186_clock = clock; // @[:@36861.4]
  assign regs_186_reset = io_reset; // @[:@36862.4 RegFile.scala 76:16:@36869.4]
  assign regs_186_io_in = 64'h0; // @[RegFile.scala 75:16:@36868.4]
  assign regs_186_io_reset = reset; // @[RegFile.scala 78:19:@36872.4]
  assign regs_186_io_enable = 1'h1; // @[RegFile.scala 74:20:@36866.4]
  assign regs_187_clock = clock; // @[:@36875.4]
  assign regs_187_reset = io_reset; // @[:@36876.4 RegFile.scala 76:16:@36883.4]
  assign regs_187_io_in = 64'h0; // @[RegFile.scala 75:16:@36882.4]
  assign regs_187_io_reset = reset; // @[RegFile.scala 78:19:@36886.4]
  assign regs_187_io_enable = 1'h1; // @[RegFile.scala 74:20:@36880.4]
  assign regs_188_clock = clock; // @[:@36889.4]
  assign regs_188_reset = io_reset; // @[:@36890.4 RegFile.scala 76:16:@36897.4]
  assign regs_188_io_in = 64'h0; // @[RegFile.scala 75:16:@36896.4]
  assign regs_188_io_reset = reset; // @[RegFile.scala 78:19:@36900.4]
  assign regs_188_io_enable = 1'h1; // @[RegFile.scala 74:20:@36894.4]
  assign regs_189_clock = clock; // @[:@36903.4]
  assign regs_189_reset = io_reset; // @[:@36904.4 RegFile.scala 76:16:@36911.4]
  assign regs_189_io_in = 64'h0; // @[RegFile.scala 75:16:@36910.4]
  assign regs_189_io_reset = reset; // @[RegFile.scala 78:19:@36914.4]
  assign regs_189_io_enable = 1'h1; // @[RegFile.scala 74:20:@36908.4]
  assign regs_190_clock = clock; // @[:@36917.4]
  assign regs_190_reset = io_reset; // @[:@36918.4 RegFile.scala 76:16:@36925.4]
  assign regs_190_io_in = 64'h0; // @[RegFile.scala 75:16:@36924.4]
  assign regs_190_io_reset = reset; // @[RegFile.scala 78:19:@36928.4]
  assign regs_190_io_enable = 1'h1; // @[RegFile.scala 74:20:@36922.4]
  assign regs_191_clock = clock; // @[:@36931.4]
  assign regs_191_reset = io_reset; // @[:@36932.4 RegFile.scala 76:16:@36939.4]
  assign regs_191_io_in = 64'h0; // @[RegFile.scala 75:16:@36938.4]
  assign regs_191_io_reset = reset; // @[RegFile.scala 78:19:@36942.4]
  assign regs_191_io_enable = 1'h1; // @[RegFile.scala 74:20:@36936.4]
  assign regs_192_clock = clock; // @[:@36945.4]
  assign regs_192_reset = io_reset; // @[:@36946.4 RegFile.scala 76:16:@36953.4]
  assign regs_192_io_in = 64'h0; // @[RegFile.scala 75:16:@36952.4]
  assign regs_192_io_reset = reset; // @[RegFile.scala 78:19:@36956.4]
  assign regs_192_io_enable = 1'h1; // @[RegFile.scala 74:20:@36950.4]
  assign regs_193_clock = clock; // @[:@36959.4]
  assign regs_193_reset = io_reset; // @[:@36960.4 RegFile.scala 76:16:@36967.4]
  assign regs_193_io_in = 64'h0; // @[RegFile.scala 75:16:@36966.4]
  assign regs_193_io_reset = reset; // @[RegFile.scala 78:19:@36970.4]
  assign regs_193_io_enable = 1'h1; // @[RegFile.scala 74:20:@36964.4]
  assign regs_194_clock = clock; // @[:@36973.4]
  assign regs_194_reset = io_reset; // @[:@36974.4 RegFile.scala 76:16:@36981.4]
  assign regs_194_io_in = 64'h0; // @[RegFile.scala 75:16:@36980.4]
  assign regs_194_io_reset = reset; // @[RegFile.scala 78:19:@36984.4]
  assign regs_194_io_enable = 1'h1; // @[RegFile.scala 74:20:@36978.4]
  assign regs_195_clock = clock; // @[:@36987.4]
  assign regs_195_reset = io_reset; // @[:@36988.4 RegFile.scala 76:16:@36995.4]
  assign regs_195_io_in = 64'h0; // @[RegFile.scala 75:16:@36994.4]
  assign regs_195_io_reset = reset; // @[RegFile.scala 78:19:@36998.4]
  assign regs_195_io_enable = 1'h1; // @[RegFile.scala 74:20:@36992.4]
  assign regs_196_clock = clock; // @[:@37001.4]
  assign regs_196_reset = io_reset; // @[:@37002.4 RegFile.scala 76:16:@37009.4]
  assign regs_196_io_in = 64'h0; // @[RegFile.scala 75:16:@37008.4]
  assign regs_196_io_reset = reset; // @[RegFile.scala 78:19:@37012.4]
  assign regs_196_io_enable = 1'h1; // @[RegFile.scala 74:20:@37006.4]
  assign regs_197_clock = clock; // @[:@37015.4]
  assign regs_197_reset = io_reset; // @[:@37016.4 RegFile.scala 76:16:@37023.4]
  assign regs_197_io_in = 64'h0; // @[RegFile.scala 75:16:@37022.4]
  assign regs_197_io_reset = reset; // @[RegFile.scala 78:19:@37026.4]
  assign regs_197_io_enable = 1'h1; // @[RegFile.scala 74:20:@37020.4]
  assign regs_198_clock = clock; // @[:@37029.4]
  assign regs_198_reset = io_reset; // @[:@37030.4 RegFile.scala 76:16:@37037.4]
  assign regs_198_io_in = 64'h0; // @[RegFile.scala 75:16:@37036.4]
  assign regs_198_io_reset = reset; // @[RegFile.scala 78:19:@37040.4]
  assign regs_198_io_enable = 1'h1; // @[RegFile.scala 74:20:@37034.4]
  assign regs_199_clock = clock; // @[:@37043.4]
  assign regs_199_reset = io_reset; // @[:@37044.4 RegFile.scala 76:16:@37051.4]
  assign regs_199_io_in = 64'h0; // @[RegFile.scala 75:16:@37050.4]
  assign regs_199_io_reset = reset; // @[RegFile.scala 78:19:@37054.4]
  assign regs_199_io_enable = 1'h1; // @[RegFile.scala 74:20:@37048.4]
  assign regs_200_clock = clock; // @[:@37057.4]
  assign regs_200_reset = io_reset; // @[:@37058.4 RegFile.scala 76:16:@37065.4]
  assign regs_200_io_in = 64'h0; // @[RegFile.scala 75:16:@37064.4]
  assign regs_200_io_reset = reset; // @[RegFile.scala 78:19:@37068.4]
  assign regs_200_io_enable = 1'h1; // @[RegFile.scala 74:20:@37062.4]
  assign regs_201_clock = clock; // @[:@37071.4]
  assign regs_201_reset = io_reset; // @[:@37072.4 RegFile.scala 76:16:@37079.4]
  assign regs_201_io_in = 64'h0; // @[RegFile.scala 75:16:@37078.4]
  assign regs_201_io_reset = reset; // @[RegFile.scala 78:19:@37082.4]
  assign regs_201_io_enable = 1'h1; // @[RegFile.scala 74:20:@37076.4]
  assign regs_202_clock = clock; // @[:@37085.4]
  assign regs_202_reset = io_reset; // @[:@37086.4 RegFile.scala 76:16:@37093.4]
  assign regs_202_io_in = 64'h0; // @[RegFile.scala 75:16:@37092.4]
  assign regs_202_io_reset = reset; // @[RegFile.scala 78:19:@37096.4]
  assign regs_202_io_enable = 1'h1; // @[RegFile.scala 74:20:@37090.4]
  assign regs_203_clock = clock; // @[:@37099.4]
  assign regs_203_reset = io_reset; // @[:@37100.4 RegFile.scala 76:16:@37107.4]
  assign regs_203_io_in = 64'h0; // @[RegFile.scala 75:16:@37106.4]
  assign regs_203_io_reset = reset; // @[RegFile.scala 78:19:@37110.4]
  assign regs_203_io_enable = 1'h1; // @[RegFile.scala 74:20:@37104.4]
  assign regs_204_clock = clock; // @[:@37113.4]
  assign regs_204_reset = io_reset; // @[:@37114.4 RegFile.scala 76:16:@37121.4]
  assign regs_204_io_in = 64'h0; // @[RegFile.scala 75:16:@37120.4]
  assign regs_204_io_reset = reset; // @[RegFile.scala 78:19:@37124.4]
  assign regs_204_io_enable = 1'h1; // @[RegFile.scala 74:20:@37118.4]
  assign regs_205_clock = clock; // @[:@37127.4]
  assign regs_205_reset = io_reset; // @[:@37128.4 RegFile.scala 76:16:@37135.4]
  assign regs_205_io_in = 64'h0; // @[RegFile.scala 75:16:@37134.4]
  assign regs_205_io_reset = reset; // @[RegFile.scala 78:19:@37138.4]
  assign regs_205_io_enable = 1'h1; // @[RegFile.scala 74:20:@37132.4]
  assign regs_206_clock = clock; // @[:@37141.4]
  assign regs_206_reset = io_reset; // @[:@37142.4 RegFile.scala 76:16:@37149.4]
  assign regs_206_io_in = 64'h0; // @[RegFile.scala 75:16:@37148.4]
  assign regs_206_io_reset = reset; // @[RegFile.scala 78:19:@37152.4]
  assign regs_206_io_enable = 1'h1; // @[RegFile.scala 74:20:@37146.4]
  assign regs_207_clock = clock; // @[:@37155.4]
  assign regs_207_reset = io_reset; // @[:@37156.4 RegFile.scala 76:16:@37163.4]
  assign regs_207_io_in = 64'h0; // @[RegFile.scala 75:16:@37162.4]
  assign regs_207_io_reset = reset; // @[RegFile.scala 78:19:@37166.4]
  assign regs_207_io_enable = 1'h1; // @[RegFile.scala 74:20:@37160.4]
  assign regs_208_clock = clock; // @[:@37169.4]
  assign regs_208_reset = io_reset; // @[:@37170.4 RegFile.scala 76:16:@37177.4]
  assign regs_208_io_in = 64'h0; // @[RegFile.scala 75:16:@37176.4]
  assign regs_208_io_reset = reset; // @[RegFile.scala 78:19:@37180.4]
  assign regs_208_io_enable = 1'h1; // @[RegFile.scala 74:20:@37174.4]
  assign regs_209_clock = clock; // @[:@37183.4]
  assign regs_209_reset = io_reset; // @[:@37184.4 RegFile.scala 76:16:@37191.4]
  assign regs_209_io_in = 64'h0; // @[RegFile.scala 75:16:@37190.4]
  assign regs_209_io_reset = reset; // @[RegFile.scala 78:19:@37194.4]
  assign regs_209_io_enable = 1'h1; // @[RegFile.scala 74:20:@37188.4]
  assign regs_210_clock = clock; // @[:@37197.4]
  assign regs_210_reset = io_reset; // @[:@37198.4 RegFile.scala 76:16:@37205.4]
  assign regs_210_io_in = 64'h0; // @[RegFile.scala 75:16:@37204.4]
  assign regs_210_io_reset = reset; // @[RegFile.scala 78:19:@37208.4]
  assign regs_210_io_enable = 1'h1; // @[RegFile.scala 74:20:@37202.4]
  assign regs_211_clock = clock; // @[:@37211.4]
  assign regs_211_reset = io_reset; // @[:@37212.4 RegFile.scala 76:16:@37219.4]
  assign regs_211_io_in = 64'h0; // @[RegFile.scala 75:16:@37218.4]
  assign regs_211_io_reset = reset; // @[RegFile.scala 78:19:@37222.4]
  assign regs_211_io_enable = 1'h1; // @[RegFile.scala 74:20:@37216.4]
  assign regs_212_clock = clock; // @[:@37225.4]
  assign regs_212_reset = io_reset; // @[:@37226.4 RegFile.scala 76:16:@37233.4]
  assign regs_212_io_in = 64'h0; // @[RegFile.scala 75:16:@37232.4]
  assign regs_212_io_reset = reset; // @[RegFile.scala 78:19:@37236.4]
  assign regs_212_io_enable = 1'h1; // @[RegFile.scala 74:20:@37230.4]
  assign regs_213_clock = clock; // @[:@37239.4]
  assign regs_213_reset = io_reset; // @[:@37240.4 RegFile.scala 76:16:@37247.4]
  assign regs_213_io_in = 64'h0; // @[RegFile.scala 75:16:@37246.4]
  assign regs_213_io_reset = reset; // @[RegFile.scala 78:19:@37250.4]
  assign regs_213_io_enable = 1'h1; // @[RegFile.scala 74:20:@37244.4]
  assign regs_214_clock = clock; // @[:@37253.4]
  assign regs_214_reset = io_reset; // @[:@37254.4 RegFile.scala 76:16:@37261.4]
  assign regs_214_io_in = 64'h0; // @[RegFile.scala 75:16:@37260.4]
  assign regs_214_io_reset = reset; // @[RegFile.scala 78:19:@37264.4]
  assign regs_214_io_enable = 1'h1; // @[RegFile.scala 74:20:@37258.4]
  assign regs_215_clock = clock; // @[:@37267.4]
  assign regs_215_reset = io_reset; // @[:@37268.4 RegFile.scala 76:16:@37275.4]
  assign regs_215_io_in = 64'h0; // @[RegFile.scala 75:16:@37274.4]
  assign regs_215_io_reset = reset; // @[RegFile.scala 78:19:@37278.4]
  assign regs_215_io_enable = 1'h1; // @[RegFile.scala 74:20:@37272.4]
  assign regs_216_clock = clock; // @[:@37281.4]
  assign regs_216_reset = io_reset; // @[:@37282.4 RegFile.scala 76:16:@37289.4]
  assign regs_216_io_in = 64'h0; // @[RegFile.scala 75:16:@37288.4]
  assign regs_216_io_reset = reset; // @[RegFile.scala 78:19:@37292.4]
  assign regs_216_io_enable = 1'h1; // @[RegFile.scala 74:20:@37286.4]
  assign regs_217_clock = clock; // @[:@37295.4]
  assign regs_217_reset = io_reset; // @[:@37296.4 RegFile.scala 76:16:@37303.4]
  assign regs_217_io_in = 64'h0; // @[RegFile.scala 75:16:@37302.4]
  assign regs_217_io_reset = reset; // @[RegFile.scala 78:19:@37306.4]
  assign regs_217_io_enable = 1'h1; // @[RegFile.scala 74:20:@37300.4]
  assign regs_218_clock = clock; // @[:@37309.4]
  assign regs_218_reset = io_reset; // @[:@37310.4 RegFile.scala 76:16:@37317.4]
  assign regs_218_io_in = 64'h0; // @[RegFile.scala 75:16:@37316.4]
  assign regs_218_io_reset = reset; // @[RegFile.scala 78:19:@37320.4]
  assign regs_218_io_enable = 1'h1; // @[RegFile.scala 74:20:@37314.4]
  assign regs_219_clock = clock; // @[:@37323.4]
  assign regs_219_reset = io_reset; // @[:@37324.4 RegFile.scala 76:16:@37331.4]
  assign regs_219_io_in = 64'h0; // @[RegFile.scala 75:16:@37330.4]
  assign regs_219_io_reset = reset; // @[RegFile.scala 78:19:@37334.4]
  assign regs_219_io_enable = 1'h1; // @[RegFile.scala 74:20:@37328.4]
  assign regs_220_clock = clock; // @[:@37337.4]
  assign regs_220_reset = io_reset; // @[:@37338.4 RegFile.scala 76:16:@37345.4]
  assign regs_220_io_in = 64'h0; // @[RegFile.scala 75:16:@37344.4]
  assign regs_220_io_reset = reset; // @[RegFile.scala 78:19:@37348.4]
  assign regs_220_io_enable = 1'h1; // @[RegFile.scala 74:20:@37342.4]
  assign regs_221_clock = clock; // @[:@37351.4]
  assign regs_221_reset = io_reset; // @[:@37352.4 RegFile.scala 76:16:@37359.4]
  assign regs_221_io_in = 64'h0; // @[RegFile.scala 75:16:@37358.4]
  assign regs_221_io_reset = reset; // @[RegFile.scala 78:19:@37362.4]
  assign regs_221_io_enable = 1'h1; // @[RegFile.scala 74:20:@37356.4]
  assign regs_222_clock = clock; // @[:@37365.4]
  assign regs_222_reset = io_reset; // @[:@37366.4 RegFile.scala 76:16:@37373.4]
  assign regs_222_io_in = 64'h0; // @[RegFile.scala 75:16:@37372.4]
  assign regs_222_io_reset = reset; // @[RegFile.scala 78:19:@37376.4]
  assign regs_222_io_enable = 1'h1; // @[RegFile.scala 74:20:@37370.4]
  assign regs_223_clock = clock; // @[:@37379.4]
  assign regs_223_reset = io_reset; // @[:@37380.4 RegFile.scala 76:16:@37387.4]
  assign regs_223_io_in = 64'h0; // @[RegFile.scala 75:16:@37386.4]
  assign regs_223_io_reset = reset; // @[RegFile.scala 78:19:@37390.4]
  assign regs_223_io_enable = 1'h1; // @[RegFile.scala 74:20:@37384.4]
  assign regs_224_clock = clock; // @[:@37393.4]
  assign regs_224_reset = io_reset; // @[:@37394.4 RegFile.scala 76:16:@37401.4]
  assign regs_224_io_in = 64'h0; // @[RegFile.scala 75:16:@37400.4]
  assign regs_224_io_reset = reset; // @[RegFile.scala 78:19:@37404.4]
  assign regs_224_io_enable = 1'h1; // @[RegFile.scala 74:20:@37398.4]
  assign regs_225_clock = clock; // @[:@37407.4]
  assign regs_225_reset = io_reset; // @[:@37408.4 RegFile.scala 76:16:@37415.4]
  assign regs_225_io_in = 64'h0; // @[RegFile.scala 75:16:@37414.4]
  assign regs_225_io_reset = reset; // @[RegFile.scala 78:19:@37418.4]
  assign regs_225_io_enable = 1'h1; // @[RegFile.scala 74:20:@37412.4]
  assign regs_226_clock = clock; // @[:@37421.4]
  assign regs_226_reset = io_reset; // @[:@37422.4 RegFile.scala 76:16:@37429.4]
  assign regs_226_io_in = 64'h0; // @[RegFile.scala 75:16:@37428.4]
  assign regs_226_io_reset = reset; // @[RegFile.scala 78:19:@37432.4]
  assign regs_226_io_enable = 1'h1; // @[RegFile.scala 74:20:@37426.4]
  assign regs_227_clock = clock; // @[:@37435.4]
  assign regs_227_reset = io_reset; // @[:@37436.4 RegFile.scala 76:16:@37443.4]
  assign regs_227_io_in = 64'h0; // @[RegFile.scala 75:16:@37442.4]
  assign regs_227_io_reset = reset; // @[RegFile.scala 78:19:@37446.4]
  assign regs_227_io_enable = 1'h1; // @[RegFile.scala 74:20:@37440.4]
  assign regs_228_clock = clock; // @[:@37449.4]
  assign regs_228_reset = io_reset; // @[:@37450.4 RegFile.scala 76:16:@37457.4]
  assign regs_228_io_in = 64'h0; // @[RegFile.scala 75:16:@37456.4]
  assign regs_228_io_reset = reset; // @[RegFile.scala 78:19:@37460.4]
  assign regs_228_io_enable = 1'h1; // @[RegFile.scala 74:20:@37454.4]
  assign regs_229_clock = clock; // @[:@37463.4]
  assign regs_229_reset = io_reset; // @[:@37464.4 RegFile.scala 76:16:@37471.4]
  assign regs_229_io_in = 64'h0; // @[RegFile.scala 75:16:@37470.4]
  assign regs_229_io_reset = reset; // @[RegFile.scala 78:19:@37474.4]
  assign regs_229_io_enable = 1'h1; // @[RegFile.scala 74:20:@37468.4]
  assign regs_230_clock = clock; // @[:@37477.4]
  assign regs_230_reset = io_reset; // @[:@37478.4 RegFile.scala 76:16:@37485.4]
  assign regs_230_io_in = 64'h0; // @[RegFile.scala 75:16:@37484.4]
  assign regs_230_io_reset = reset; // @[RegFile.scala 78:19:@37488.4]
  assign regs_230_io_enable = 1'h1; // @[RegFile.scala 74:20:@37482.4]
  assign regs_231_clock = clock; // @[:@37491.4]
  assign regs_231_reset = io_reset; // @[:@37492.4 RegFile.scala 76:16:@37499.4]
  assign regs_231_io_in = 64'h0; // @[RegFile.scala 75:16:@37498.4]
  assign regs_231_io_reset = reset; // @[RegFile.scala 78:19:@37502.4]
  assign regs_231_io_enable = 1'h1; // @[RegFile.scala 74:20:@37496.4]
  assign regs_232_clock = clock; // @[:@37505.4]
  assign regs_232_reset = io_reset; // @[:@37506.4 RegFile.scala 76:16:@37513.4]
  assign regs_232_io_in = 64'h0; // @[RegFile.scala 75:16:@37512.4]
  assign regs_232_io_reset = reset; // @[RegFile.scala 78:19:@37516.4]
  assign regs_232_io_enable = 1'h1; // @[RegFile.scala 74:20:@37510.4]
  assign regs_233_clock = clock; // @[:@37519.4]
  assign regs_233_reset = io_reset; // @[:@37520.4 RegFile.scala 76:16:@37527.4]
  assign regs_233_io_in = 64'h0; // @[RegFile.scala 75:16:@37526.4]
  assign regs_233_io_reset = reset; // @[RegFile.scala 78:19:@37530.4]
  assign regs_233_io_enable = 1'h1; // @[RegFile.scala 74:20:@37524.4]
  assign regs_234_clock = clock; // @[:@37533.4]
  assign regs_234_reset = io_reset; // @[:@37534.4 RegFile.scala 76:16:@37541.4]
  assign regs_234_io_in = 64'h0; // @[RegFile.scala 75:16:@37540.4]
  assign regs_234_io_reset = reset; // @[RegFile.scala 78:19:@37544.4]
  assign regs_234_io_enable = 1'h1; // @[RegFile.scala 74:20:@37538.4]
  assign regs_235_clock = clock; // @[:@37547.4]
  assign regs_235_reset = io_reset; // @[:@37548.4 RegFile.scala 76:16:@37555.4]
  assign regs_235_io_in = 64'h0; // @[RegFile.scala 75:16:@37554.4]
  assign regs_235_io_reset = reset; // @[RegFile.scala 78:19:@37558.4]
  assign regs_235_io_enable = 1'h1; // @[RegFile.scala 74:20:@37552.4]
  assign regs_236_clock = clock; // @[:@37561.4]
  assign regs_236_reset = io_reset; // @[:@37562.4 RegFile.scala 76:16:@37569.4]
  assign regs_236_io_in = 64'h0; // @[RegFile.scala 75:16:@37568.4]
  assign regs_236_io_reset = reset; // @[RegFile.scala 78:19:@37572.4]
  assign regs_236_io_enable = 1'h1; // @[RegFile.scala 74:20:@37566.4]
  assign regs_237_clock = clock; // @[:@37575.4]
  assign regs_237_reset = io_reset; // @[:@37576.4 RegFile.scala 76:16:@37583.4]
  assign regs_237_io_in = 64'h0; // @[RegFile.scala 75:16:@37582.4]
  assign regs_237_io_reset = reset; // @[RegFile.scala 78:19:@37586.4]
  assign regs_237_io_enable = 1'h1; // @[RegFile.scala 74:20:@37580.4]
  assign regs_238_clock = clock; // @[:@37589.4]
  assign regs_238_reset = io_reset; // @[:@37590.4 RegFile.scala 76:16:@37597.4]
  assign regs_238_io_in = 64'h0; // @[RegFile.scala 75:16:@37596.4]
  assign regs_238_io_reset = reset; // @[RegFile.scala 78:19:@37600.4]
  assign regs_238_io_enable = 1'h1; // @[RegFile.scala 74:20:@37594.4]
  assign regs_239_clock = clock; // @[:@37603.4]
  assign regs_239_reset = io_reset; // @[:@37604.4 RegFile.scala 76:16:@37611.4]
  assign regs_239_io_in = 64'h0; // @[RegFile.scala 75:16:@37610.4]
  assign regs_239_io_reset = reset; // @[RegFile.scala 78:19:@37614.4]
  assign regs_239_io_enable = 1'h1; // @[RegFile.scala 74:20:@37608.4]
  assign regs_240_clock = clock; // @[:@37617.4]
  assign regs_240_reset = io_reset; // @[:@37618.4 RegFile.scala 76:16:@37625.4]
  assign regs_240_io_in = 64'h0; // @[RegFile.scala 75:16:@37624.4]
  assign regs_240_io_reset = reset; // @[RegFile.scala 78:19:@37628.4]
  assign regs_240_io_enable = 1'h1; // @[RegFile.scala 74:20:@37622.4]
  assign regs_241_clock = clock; // @[:@37631.4]
  assign regs_241_reset = io_reset; // @[:@37632.4 RegFile.scala 76:16:@37639.4]
  assign regs_241_io_in = 64'h0; // @[RegFile.scala 75:16:@37638.4]
  assign regs_241_io_reset = reset; // @[RegFile.scala 78:19:@37642.4]
  assign regs_241_io_enable = 1'h1; // @[RegFile.scala 74:20:@37636.4]
  assign regs_242_clock = clock; // @[:@37645.4]
  assign regs_242_reset = io_reset; // @[:@37646.4 RegFile.scala 76:16:@37653.4]
  assign regs_242_io_in = 64'h0; // @[RegFile.scala 75:16:@37652.4]
  assign regs_242_io_reset = reset; // @[RegFile.scala 78:19:@37656.4]
  assign regs_242_io_enable = 1'h1; // @[RegFile.scala 74:20:@37650.4]
  assign regs_243_clock = clock; // @[:@37659.4]
  assign regs_243_reset = io_reset; // @[:@37660.4 RegFile.scala 76:16:@37667.4]
  assign regs_243_io_in = 64'h0; // @[RegFile.scala 75:16:@37666.4]
  assign regs_243_io_reset = reset; // @[RegFile.scala 78:19:@37670.4]
  assign regs_243_io_enable = 1'h1; // @[RegFile.scala 74:20:@37664.4]
  assign regs_244_clock = clock; // @[:@37673.4]
  assign regs_244_reset = io_reset; // @[:@37674.4 RegFile.scala 76:16:@37681.4]
  assign regs_244_io_in = 64'h0; // @[RegFile.scala 75:16:@37680.4]
  assign regs_244_io_reset = reset; // @[RegFile.scala 78:19:@37684.4]
  assign regs_244_io_enable = 1'h1; // @[RegFile.scala 74:20:@37678.4]
  assign regs_245_clock = clock; // @[:@37687.4]
  assign regs_245_reset = io_reset; // @[:@37688.4 RegFile.scala 76:16:@37695.4]
  assign regs_245_io_in = 64'h0; // @[RegFile.scala 75:16:@37694.4]
  assign regs_245_io_reset = reset; // @[RegFile.scala 78:19:@37698.4]
  assign regs_245_io_enable = 1'h1; // @[RegFile.scala 74:20:@37692.4]
  assign regs_246_clock = clock; // @[:@37701.4]
  assign regs_246_reset = io_reset; // @[:@37702.4 RegFile.scala 76:16:@37709.4]
  assign regs_246_io_in = 64'h0; // @[RegFile.scala 75:16:@37708.4]
  assign regs_246_io_reset = reset; // @[RegFile.scala 78:19:@37712.4]
  assign regs_246_io_enable = 1'h1; // @[RegFile.scala 74:20:@37706.4]
  assign regs_247_clock = clock; // @[:@37715.4]
  assign regs_247_reset = io_reset; // @[:@37716.4 RegFile.scala 76:16:@37723.4]
  assign regs_247_io_in = 64'h0; // @[RegFile.scala 75:16:@37722.4]
  assign regs_247_io_reset = reset; // @[RegFile.scala 78:19:@37726.4]
  assign regs_247_io_enable = 1'h1; // @[RegFile.scala 74:20:@37720.4]
  assign regs_248_clock = clock; // @[:@37729.4]
  assign regs_248_reset = io_reset; // @[:@37730.4 RegFile.scala 76:16:@37737.4]
  assign regs_248_io_in = 64'h0; // @[RegFile.scala 75:16:@37736.4]
  assign regs_248_io_reset = reset; // @[RegFile.scala 78:19:@37740.4]
  assign regs_248_io_enable = 1'h1; // @[RegFile.scala 74:20:@37734.4]
  assign regs_249_clock = clock; // @[:@37743.4]
  assign regs_249_reset = io_reset; // @[:@37744.4 RegFile.scala 76:16:@37751.4]
  assign regs_249_io_in = 64'h0; // @[RegFile.scala 75:16:@37750.4]
  assign regs_249_io_reset = reset; // @[RegFile.scala 78:19:@37754.4]
  assign regs_249_io_enable = 1'h1; // @[RegFile.scala 74:20:@37748.4]
  assign regs_250_clock = clock; // @[:@37757.4]
  assign regs_250_reset = io_reset; // @[:@37758.4 RegFile.scala 76:16:@37765.4]
  assign regs_250_io_in = 64'h0; // @[RegFile.scala 75:16:@37764.4]
  assign regs_250_io_reset = reset; // @[RegFile.scala 78:19:@37768.4]
  assign regs_250_io_enable = 1'h1; // @[RegFile.scala 74:20:@37762.4]
  assign regs_251_clock = clock; // @[:@37771.4]
  assign regs_251_reset = io_reset; // @[:@37772.4 RegFile.scala 76:16:@37779.4]
  assign regs_251_io_in = 64'h0; // @[RegFile.scala 75:16:@37778.4]
  assign regs_251_io_reset = reset; // @[RegFile.scala 78:19:@37782.4]
  assign regs_251_io_enable = 1'h1; // @[RegFile.scala 74:20:@37776.4]
  assign regs_252_clock = clock; // @[:@37785.4]
  assign regs_252_reset = io_reset; // @[:@37786.4 RegFile.scala 76:16:@37793.4]
  assign regs_252_io_in = 64'h0; // @[RegFile.scala 75:16:@37792.4]
  assign regs_252_io_reset = reset; // @[RegFile.scala 78:19:@37796.4]
  assign regs_252_io_enable = 1'h1; // @[RegFile.scala 74:20:@37790.4]
  assign regs_253_clock = clock; // @[:@37799.4]
  assign regs_253_reset = io_reset; // @[:@37800.4 RegFile.scala 76:16:@37807.4]
  assign regs_253_io_in = 64'h0; // @[RegFile.scala 75:16:@37806.4]
  assign regs_253_io_reset = reset; // @[RegFile.scala 78:19:@37810.4]
  assign regs_253_io_enable = 1'h1; // @[RegFile.scala 74:20:@37804.4]
  assign regs_254_clock = clock; // @[:@37813.4]
  assign regs_254_reset = io_reset; // @[:@37814.4 RegFile.scala 76:16:@37821.4]
  assign regs_254_io_in = 64'h0; // @[RegFile.scala 75:16:@37820.4]
  assign regs_254_io_reset = reset; // @[RegFile.scala 78:19:@37824.4]
  assign regs_254_io_enable = 1'h1; // @[RegFile.scala 74:20:@37818.4]
  assign regs_255_clock = clock; // @[:@37827.4]
  assign regs_255_reset = io_reset; // @[:@37828.4 RegFile.scala 76:16:@37835.4]
  assign regs_255_io_in = 64'h0; // @[RegFile.scala 75:16:@37834.4]
  assign regs_255_io_reset = reset; // @[RegFile.scala 78:19:@37838.4]
  assign regs_255_io_enable = 1'h1; // @[RegFile.scala 74:20:@37832.4]
  assign regs_256_clock = clock; // @[:@37841.4]
  assign regs_256_reset = io_reset; // @[:@37842.4 RegFile.scala 76:16:@37849.4]
  assign regs_256_io_in = 64'h0; // @[RegFile.scala 75:16:@37848.4]
  assign regs_256_io_reset = reset; // @[RegFile.scala 78:19:@37852.4]
  assign regs_256_io_enable = 1'h1; // @[RegFile.scala 74:20:@37846.4]
  assign regs_257_clock = clock; // @[:@37855.4]
  assign regs_257_reset = io_reset; // @[:@37856.4 RegFile.scala 76:16:@37863.4]
  assign regs_257_io_in = 64'h0; // @[RegFile.scala 75:16:@37862.4]
  assign regs_257_io_reset = reset; // @[RegFile.scala 78:19:@37866.4]
  assign regs_257_io_enable = 1'h1; // @[RegFile.scala 74:20:@37860.4]
  assign regs_258_clock = clock; // @[:@37869.4]
  assign regs_258_reset = io_reset; // @[:@37870.4 RegFile.scala 76:16:@37877.4]
  assign regs_258_io_in = 64'h0; // @[RegFile.scala 75:16:@37876.4]
  assign regs_258_io_reset = reset; // @[RegFile.scala 78:19:@37880.4]
  assign regs_258_io_enable = 1'h1; // @[RegFile.scala 74:20:@37874.4]
  assign regs_259_clock = clock; // @[:@37883.4]
  assign regs_259_reset = io_reset; // @[:@37884.4 RegFile.scala 76:16:@37891.4]
  assign regs_259_io_in = 64'h0; // @[RegFile.scala 75:16:@37890.4]
  assign regs_259_io_reset = reset; // @[RegFile.scala 78:19:@37894.4]
  assign regs_259_io_enable = 1'h1; // @[RegFile.scala 74:20:@37888.4]
  assign regs_260_clock = clock; // @[:@37897.4]
  assign regs_260_reset = io_reset; // @[:@37898.4 RegFile.scala 76:16:@37905.4]
  assign regs_260_io_in = 64'h0; // @[RegFile.scala 75:16:@37904.4]
  assign regs_260_io_reset = reset; // @[RegFile.scala 78:19:@37908.4]
  assign regs_260_io_enable = 1'h1; // @[RegFile.scala 74:20:@37902.4]
  assign regs_261_clock = clock; // @[:@37911.4]
  assign regs_261_reset = io_reset; // @[:@37912.4 RegFile.scala 76:16:@37919.4]
  assign regs_261_io_in = 64'h0; // @[RegFile.scala 75:16:@37918.4]
  assign regs_261_io_reset = reset; // @[RegFile.scala 78:19:@37922.4]
  assign regs_261_io_enable = 1'h1; // @[RegFile.scala 74:20:@37916.4]
  assign regs_262_clock = clock; // @[:@37925.4]
  assign regs_262_reset = io_reset; // @[:@37926.4 RegFile.scala 76:16:@37933.4]
  assign regs_262_io_in = 64'h0; // @[RegFile.scala 75:16:@37932.4]
  assign regs_262_io_reset = reset; // @[RegFile.scala 78:19:@37936.4]
  assign regs_262_io_enable = 1'h1; // @[RegFile.scala 74:20:@37930.4]
  assign regs_263_clock = clock; // @[:@37939.4]
  assign regs_263_reset = io_reset; // @[:@37940.4 RegFile.scala 76:16:@37947.4]
  assign regs_263_io_in = 64'h0; // @[RegFile.scala 75:16:@37946.4]
  assign regs_263_io_reset = reset; // @[RegFile.scala 78:19:@37950.4]
  assign regs_263_io_enable = 1'h1; // @[RegFile.scala 74:20:@37944.4]
  assign regs_264_clock = clock; // @[:@37953.4]
  assign regs_264_reset = io_reset; // @[:@37954.4 RegFile.scala 76:16:@37961.4]
  assign regs_264_io_in = 64'h0; // @[RegFile.scala 75:16:@37960.4]
  assign regs_264_io_reset = reset; // @[RegFile.scala 78:19:@37964.4]
  assign regs_264_io_enable = 1'h1; // @[RegFile.scala 74:20:@37958.4]
  assign regs_265_clock = clock; // @[:@37967.4]
  assign regs_265_reset = io_reset; // @[:@37968.4 RegFile.scala 76:16:@37975.4]
  assign regs_265_io_in = 64'h0; // @[RegFile.scala 75:16:@37974.4]
  assign regs_265_io_reset = reset; // @[RegFile.scala 78:19:@37978.4]
  assign regs_265_io_enable = 1'h1; // @[RegFile.scala 74:20:@37972.4]
  assign regs_266_clock = clock; // @[:@37981.4]
  assign regs_266_reset = io_reset; // @[:@37982.4 RegFile.scala 76:16:@37989.4]
  assign regs_266_io_in = 64'h0; // @[RegFile.scala 75:16:@37988.4]
  assign regs_266_io_reset = reset; // @[RegFile.scala 78:19:@37992.4]
  assign regs_266_io_enable = 1'h1; // @[RegFile.scala 74:20:@37986.4]
  assign regs_267_clock = clock; // @[:@37995.4]
  assign regs_267_reset = io_reset; // @[:@37996.4 RegFile.scala 76:16:@38003.4]
  assign regs_267_io_in = 64'h0; // @[RegFile.scala 75:16:@38002.4]
  assign regs_267_io_reset = reset; // @[RegFile.scala 78:19:@38006.4]
  assign regs_267_io_enable = 1'h1; // @[RegFile.scala 74:20:@38000.4]
  assign regs_268_clock = clock; // @[:@38009.4]
  assign regs_268_reset = io_reset; // @[:@38010.4 RegFile.scala 76:16:@38017.4]
  assign regs_268_io_in = 64'h0; // @[RegFile.scala 75:16:@38016.4]
  assign regs_268_io_reset = reset; // @[RegFile.scala 78:19:@38020.4]
  assign regs_268_io_enable = 1'h1; // @[RegFile.scala 74:20:@38014.4]
  assign regs_269_clock = clock; // @[:@38023.4]
  assign regs_269_reset = io_reset; // @[:@38024.4 RegFile.scala 76:16:@38031.4]
  assign regs_269_io_in = 64'h0; // @[RegFile.scala 75:16:@38030.4]
  assign regs_269_io_reset = reset; // @[RegFile.scala 78:19:@38034.4]
  assign regs_269_io_enable = 1'h1; // @[RegFile.scala 74:20:@38028.4]
  assign regs_270_clock = clock; // @[:@38037.4]
  assign regs_270_reset = io_reset; // @[:@38038.4 RegFile.scala 76:16:@38045.4]
  assign regs_270_io_in = 64'h0; // @[RegFile.scala 75:16:@38044.4]
  assign regs_270_io_reset = reset; // @[RegFile.scala 78:19:@38048.4]
  assign regs_270_io_enable = 1'h1; // @[RegFile.scala 74:20:@38042.4]
  assign regs_271_clock = clock; // @[:@38051.4]
  assign regs_271_reset = io_reset; // @[:@38052.4 RegFile.scala 76:16:@38059.4]
  assign regs_271_io_in = 64'h0; // @[RegFile.scala 75:16:@38058.4]
  assign regs_271_io_reset = reset; // @[RegFile.scala 78:19:@38062.4]
  assign regs_271_io_enable = 1'h1; // @[RegFile.scala 74:20:@38056.4]
  assign regs_272_clock = clock; // @[:@38065.4]
  assign regs_272_reset = io_reset; // @[:@38066.4 RegFile.scala 76:16:@38073.4]
  assign regs_272_io_in = 64'h0; // @[RegFile.scala 75:16:@38072.4]
  assign regs_272_io_reset = reset; // @[RegFile.scala 78:19:@38076.4]
  assign regs_272_io_enable = 1'h1; // @[RegFile.scala 74:20:@38070.4]
  assign regs_273_clock = clock; // @[:@38079.4]
  assign regs_273_reset = io_reset; // @[:@38080.4 RegFile.scala 76:16:@38087.4]
  assign regs_273_io_in = 64'h0; // @[RegFile.scala 75:16:@38086.4]
  assign regs_273_io_reset = reset; // @[RegFile.scala 78:19:@38090.4]
  assign regs_273_io_enable = 1'h1; // @[RegFile.scala 74:20:@38084.4]
  assign regs_274_clock = clock; // @[:@38093.4]
  assign regs_274_reset = io_reset; // @[:@38094.4 RegFile.scala 76:16:@38101.4]
  assign regs_274_io_in = 64'h0; // @[RegFile.scala 75:16:@38100.4]
  assign regs_274_io_reset = reset; // @[RegFile.scala 78:19:@38104.4]
  assign regs_274_io_enable = 1'h1; // @[RegFile.scala 74:20:@38098.4]
  assign regs_275_clock = clock; // @[:@38107.4]
  assign regs_275_reset = io_reset; // @[:@38108.4 RegFile.scala 76:16:@38115.4]
  assign regs_275_io_in = 64'h0; // @[RegFile.scala 75:16:@38114.4]
  assign regs_275_io_reset = reset; // @[RegFile.scala 78:19:@38118.4]
  assign regs_275_io_enable = 1'h1; // @[RegFile.scala 74:20:@38112.4]
  assign regs_276_clock = clock; // @[:@38121.4]
  assign regs_276_reset = io_reset; // @[:@38122.4 RegFile.scala 76:16:@38129.4]
  assign regs_276_io_in = 64'h0; // @[RegFile.scala 75:16:@38128.4]
  assign regs_276_io_reset = reset; // @[RegFile.scala 78:19:@38132.4]
  assign regs_276_io_enable = 1'h1; // @[RegFile.scala 74:20:@38126.4]
  assign regs_277_clock = clock; // @[:@38135.4]
  assign regs_277_reset = io_reset; // @[:@38136.4 RegFile.scala 76:16:@38143.4]
  assign regs_277_io_in = 64'h0; // @[RegFile.scala 75:16:@38142.4]
  assign regs_277_io_reset = reset; // @[RegFile.scala 78:19:@38146.4]
  assign regs_277_io_enable = 1'h1; // @[RegFile.scala 74:20:@38140.4]
  assign regs_278_clock = clock; // @[:@38149.4]
  assign regs_278_reset = io_reset; // @[:@38150.4 RegFile.scala 76:16:@38157.4]
  assign regs_278_io_in = 64'h0; // @[RegFile.scala 75:16:@38156.4]
  assign regs_278_io_reset = reset; // @[RegFile.scala 78:19:@38160.4]
  assign regs_278_io_enable = 1'h1; // @[RegFile.scala 74:20:@38154.4]
  assign regs_279_clock = clock; // @[:@38163.4]
  assign regs_279_reset = io_reset; // @[:@38164.4 RegFile.scala 76:16:@38171.4]
  assign regs_279_io_in = 64'h0; // @[RegFile.scala 75:16:@38170.4]
  assign regs_279_io_reset = reset; // @[RegFile.scala 78:19:@38174.4]
  assign regs_279_io_enable = 1'h1; // @[RegFile.scala 74:20:@38168.4]
  assign regs_280_clock = clock; // @[:@38177.4]
  assign regs_280_reset = io_reset; // @[:@38178.4 RegFile.scala 76:16:@38185.4]
  assign regs_280_io_in = 64'h0; // @[RegFile.scala 75:16:@38184.4]
  assign regs_280_io_reset = reset; // @[RegFile.scala 78:19:@38188.4]
  assign regs_280_io_enable = 1'h1; // @[RegFile.scala 74:20:@38182.4]
  assign regs_281_clock = clock; // @[:@38191.4]
  assign regs_281_reset = io_reset; // @[:@38192.4 RegFile.scala 76:16:@38199.4]
  assign regs_281_io_in = 64'h0; // @[RegFile.scala 75:16:@38198.4]
  assign regs_281_io_reset = reset; // @[RegFile.scala 78:19:@38202.4]
  assign regs_281_io_enable = 1'h1; // @[RegFile.scala 74:20:@38196.4]
  assign regs_282_clock = clock; // @[:@38205.4]
  assign regs_282_reset = io_reset; // @[:@38206.4 RegFile.scala 76:16:@38213.4]
  assign regs_282_io_in = 64'h0; // @[RegFile.scala 75:16:@38212.4]
  assign regs_282_io_reset = reset; // @[RegFile.scala 78:19:@38216.4]
  assign regs_282_io_enable = 1'h1; // @[RegFile.scala 74:20:@38210.4]
  assign regs_283_clock = clock; // @[:@38219.4]
  assign regs_283_reset = io_reset; // @[:@38220.4 RegFile.scala 76:16:@38227.4]
  assign regs_283_io_in = 64'h0; // @[RegFile.scala 75:16:@38226.4]
  assign regs_283_io_reset = reset; // @[RegFile.scala 78:19:@38230.4]
  assign regs_283_io_enable = 1'h1; // @[RegFile.scala 74:20:@38224.4]
  assign regs_284_clock = clock; // @[:@38233.4]
  assign regs_284_reset = io_reset; // @[:@38234.4 RegFile.scala 76:16:@38241.4]
  assign regs_284_io_in = 64'h0; // @[RegFile.scala 75:16:@38240.4]
  assign regs_284_io_reset = reset; // @[RegFile.scala 78:19:@38244.4]
  assign regs_284_io_enable = 1'h1; // @[RegFile.scala 74:20:@38238.4]
  assign regs_285_clock = clock; // @[:@38247.4]
  assign regs_285_reset = io_reset; // @[:@38248.4 RegFile.scala 76:16:@38255.4]
  assign regs_285_io_in = 64'h0; // @[RegFile.scala 75:16:@38254.4]
  assign regs_285_io_reset = reset; // @[RegFile.scala 78:19:@38258.4]
  assign regs_285_io_enable = 1'h1; // @[RegFile.scala 74:20:@38252.4]
  assign regs_286_clock = clock; // @[:@38261.4]
  assign regs_286_reset = io_reset; // @[:@38262.4 RegFile.scala 76:16:@38269.4]
  assign regs_286_io_in = 64'h0; // @[RegFile.scala 75:16:@38268.4]
  assign regs_286_io_reset = reset; // @[RegFile.scala 78:19:@38272.4]
  assign regs_286_io_enable = 1'h1; // @[RegFile.scala 74:20:@38266.4]
  assign regs_287_clock = clock; // @[:@38275.4]
  assign regs_287_reset = io_reset; // @[:@38276.4 RegFile.scala 76:16:@38283.4]
  assign regs_287_io_in = 64'h0; // @[RegFile.scala 75:16:@38282.4]
  assign regs_287_io_reset = reset; // @[RegFile.scala 78:19:@38286.4]
  assign regs_287_io_enable = 1'h1; // @[RegFile.scala 74:20:@38280.4]
  assign regs_288_clock = clock; // @[:@38289.4]
  assign regs_288_reset = io_reset; // @[:@38290.4 RegFile.scala 76:16:@38297.4]
  assign regs_288_io_in = 64'h0; // @[RegFile.scala 75:16:@38296.4]
  assign regs_288_io_reset = reset; // @[RegFile.scala 78:19:@38300.4]
  assign regs_288_io_enable = 1'h1; // @[RegFile.scala 74:20:@38294.4]
  assign regs_289_clock = clock; // @[:@38303.4]
  assign regs_289_reset = io_reset; // @[:@38304.4 RegFile.scala 76:16:@38311.4]
  assign regs_289_io_in = 64'h0; // @[RegFile.scala 75:16:@38310.4]
  assign regs_289_io_reset = reset; // @[RegFile.scala 78:19:@38314.4]
  assign regs_289_io_enable = 1'h1; // @[RegFile.scala 74:20:@38308.4]
  assign regs_290_clock = clock; // @[:@38317.4]
  assign regs_290_reset = io_reset; // @[:@38318.4 RegFile.scala 76:16:@38325.4]
  assign regs_290_io_in = 64'h0; // @[RegFile.scala 75:16:@38324.4]
  assign regs_290_io_reset = reset; // @[RegFile.scala 78:19:@38328.4]
  assign regs_290_io_enable = 1'h1; // @[RegFile.scala 74:20:@38322.4]
  assign regs_291_clock = clock; // @[:@38331.4]
  assign regs_291_reset = io_reset; // @[:@38332.4 RegFile.scala 76:16:@38339.4]
  assign regs_291_io_in = 64'h0; // @[RegFile.scala 75:16:@38338.4]
  assign regs_291_io_reset = reset; // @[RegFile.scala 78:19:@38342.4]
  assign regs_291_io_enable = 1'h1; // @[RegFile.scala 74:20:@38336.4]
  assign regs_292_clock = clock; // @[:@38345.4]
  assign regs_292_reset = io_reset; // @[:@38346.4 RegFile.scala 76:16:@38353.4]
  assign regs_292_io_in = 64'h0; // @[RegFile.scala 75:16:@38352.4]
  assign regs_292_io_reset = reset; // @[RegFile.scala 78:19:@38356.4]
  assign regs_292_io_enable = 1'h1; // @[RegFile.scala 74:20:@38350.4]
  assign regs_293_clock = clock; // @[:@38359.4]
  assign regs_293_reset = io_reset; // @[:@38360.4 RegFile.scala 76:16:@38367.4]
  assign regs_293_io_in = 64'h0; // @[RegFile.scala 75:16:@38366.4]
  assign regs_293_io_reset = reset; // @[RegFile.scala 78:19:@38370.4]
  assign regs_293_io_enable = 1'h1; // @[RegFile.scala 74:20:@38364.4]
  assign regs_294_clock = clock; // @[:@38373.4]
  assign regs_294_reset = io_reset; // @[:@38374.4 RegFile.scala 76:16:@38381.4]
  assign regs_294_io_in = 64'h0; // @[RegFile.scala 75:16:@38380.4]
  assign regs_294_io_reset = reset; // @[RegFile.scala 78:19:@38384.4]
  assign regs_294_io_enable = 1'h1; // @[RegFile.scala 74:20:@38378.4]
  assign regs_295_clock = clock; // @[:@38387.4]
  assign regs_295_reset = io_reset; // @[:@38388.4 RegFile.scala 76:16:@38395.4]
  assign regs_295_io_in = 64'h0; // @[RegFile.scala 75:16:@38394.4]
  assign regs_295_io_reset = reset; // @[RegFile.scala 78:19:@38398.4]
  assign regs_295_io_enable = 1'h1; // @[RegFile.scala 74:20:@38392.4]
  assign regs_296_clock = clock; // @[:@38401.4]
  assign regs_296_reset = io_reset; // @[:@38402.4 RegFile.scala 76:16:@38409.4]
  assign regs_296_io_in = 64'h0; // @[RegFile.scala 75:16:@38408.4]
  assign regs_296_io_reset = reset; // @[RegFile.scala 78:19:@38412.4]
  assign regs_296_io_enable = 1'h1; // @[RegFile.scala 74:20:@38406.4]
  assign regs_297_clock = clock; // @[:@38415.4]
  assign regs_297_reset = io_reset; // @[:@38416.4 RegFile.scala 76:16:@38423.4]
  assign regs_297_io_in = 64'h0; // @[RegFile.scala 75:16:@38422.4]
  assign regs_297_io_reset = reset; // @[RegFile.scala 78:19:@38426.4]
  assign regs_297_io_enable = 1'h1; // @[RegFile.scala 74:20:@38420.4]
  assign regs_298_clock = clock; // @[:@38429.4]
  assign regs_298_reset = io_reset; // @[:@38430.4 RegFile.scala 76:16:@38437.4]
  assign regs_298_io_in = 64'h0; // @[RegFile.scala 75:16:@38436.4]
  assign regs_298_io_reset = reset; // @[RegFile.scala 78:19:@38440.4]
  assign regs_298_io_enable = 1'h1; // @[RegFile.scala 74:20:@38434.4]
  assign regs_299_clock = clock; // @[:@38443.4]
  assign regs_299_reset = io_reset; // @[:@38444.4 RegFile.scala 76:16:@38451.4]
  assign regs_299_io_in = 64'h0; // @[RegFile.scala 75:16:@38450.4]
  assign regs_299_io_reset = reset; // @[RegFile.scala 78:19:@38454.4]
  assign regs_299_io_enable = 1'h1; // @[RegFile.scala 74:20:@38448.4]
  assign regs_300_clock = clock; // @[:@38457.4]
  assign regs_300_reset = io_reset; // @[:@38458.4 RegFile.scala 76:16:@38465.4]
  assign regs_300_io_in = 64'h0; // @[RegFile.scala 75:16:@38464.4]
  assign regs_300_io_reset = reset; // @[RegFile.scala 78:19:@38468.4]
  assign regs_300_io_enable = 1'h1; // @[RegFile.scala 74:20:@38462.4]
  assign regs_301_clock = clock; // @[:@38471.4]
  assign regs_301_reset = io_reset; // @[:@38472.4 RegFile.scala 76:16:@38479.4]
  assign regs_301_io_in = 64'h0; // @[RegFile.scala 75:16:@38478.4]
  assign regs_301_io_reset = reset; // @[RegFile.scala 78:19:@38482.4]
  assign regs_301_io_enable = 1'h1; // @[RegFile.scala 74:20:@38476.4]
  assign regs_302_clock = clock; // @[:@38485.4]
  assign regs_302_reset = io_reset; // @[:@38486.4 RegFile.scala 76:16:@38493.4]
  assign regs_302_io_in = 64'h0; // @[RegFile.scala 75:16:@38492.4]
  assign regs_302_io_reset = reset; // @[RegFile.scala 78:19:@38496.4]
  assign regs_302_io_enable = 1'h1; // @[RegFile.scala 74:20:@38490.4]
  assign regs_303_clock = clock; // @[:@38499.4]
  assign regs_303_reset = io_reset; // @[:@38500.4 RegFile.scala 76:16:@38507.4]
  assign regs_303_io_in = 64'h0; // @[RegFile.scala 75:16:@38506.4]
  assign regs_303_io_reset = reset; // @[RegFile.scala 78:19:@38510.4]
  assign regs_303_io_enable = 1'h1; // @[RegFile.scala 74:20:@38504.4]
  assign regs_304_clock = clock; // @[:@38513.4]
  assign regs_304_reset = io_reset; // @[:@38514.4 RegFile.scala 76:16:@38521.4]
  assign regs_304_io_in = 64'h0; // @[RegFile.scala 75:16:@38520.4]
  assign regs_304_io_reset = reset; // @[RegFile.scala 78:19:@38524.4]
  assign regs_304_io_enable = 1'h1; // @[RegFile.scala 74:20:@38518.4]
  assign regs_305_clock = clock; // @[:@38527.4]
  assign regs_305_reset = io_reset; // @[:@38528.4 RegFile.scala 76:16:@38535.4]
  assign regs_305_io_in = 64'h0; // @[RegFile.scala 75:16:@38534.4]
  assign regs_305_io_reset = reset; // @[RegFile.scala 78:19:@38538.4]
  assign regs_305_io_enable = 1'h1; // @[RegFile.scala 74:20:@38532.4]
  assign regs_306_clock = clock; // @[:@38541.4]
  assign regs_306_reset = io_reset; // @[:@38542.4 RegFile.scala 76:16:@38549.4]
  assign regs_306_io_in = 64'h0; // @[RegFile.scala 75:16:@38548.4]
  assign regs_306_io_reset = reset; // @[RegFile.scala 78:19:@38552.4]
  assign regs_306_io_enable = 1'h1; // @[RegFile.scala 74:20:@38546.4]
  assign regs_307_clock = clock; // @[:@38555.4]
  assign regs_307_reset = io_reset; // @[:@38556.4 RegFile.scala 76:16:@38563.4]
  assign regs_307_io_in = 64'h0; // @[RegFile.scala 75:16:@38562.4]
  assign regs_307_io_reset = reset; // @[RegFile.scala 78:19:@38566.4]
  assign regs_307_io_enable = 1'h1; // @[RegFile.scala 74:20:@38560.4]
  assign regs_308_clock = clock; // @[:@38569.4]
  assign regs_308_reset = io_reset; // @[:@38570.4 RegFile.scala 76:16:@38577.4]
  assign regs_308_io_in = 64'h0; // @[RegFile.scala 75:16:@38576.4]
  assign regs_308_io_reset = reset; // @[RegFile.scala 78:19:@38580.4]
  assign regs_308_io_enable = 1'h1; // @[RegFile.scala 74:20:@38574.4]
  assign regs_309_clock = clock; // @[:@38583.4]
  assign regs_309_reset = io_reset; // @[:@38584.4 RegFile.scala 76:16:@38591.4]
  assign regs_309_io_in = 64'h0; // @[RegFile.scala 75:16:@38590.4]
  assign regs_309_io_reset = reset; // @[RegFile.scala 78:19:@38594.4]
  assign regs_309_io_enable = 1'h1; // @[RegFile.scala 74:20:@38588.4]
  assign regs_310_clock = clock; // @[:@38597.4]
  assign regs_310_reset = io_reset; // @[:@38598.4 RegFile.scala 76:16:@38605.4]
  assign regs_310_io_in = 64'h0; // @[RegFile.scala 75:16:@38604.4]
  assign regs_310_io_reset = reset; // @[RegFile.scala 78:19:@38608.4]
  assign regs_310_io_enable = 1'h1; // @[RegFile.scala 74:20:@38602.4]
  assign regs_311_clock = clock; // @[:@38611.4]
  assign regs_311_reset = io_reset; // @[:@38612.4 RegFile.scala 76:16:@38619.4]
  assign regs_311_io_in = 64'h0; // @[RegFile.scala 75:16:@38618.4]
  assign regs_311_io_reset = reset; // @[RegFile.scala 78:19:@38622.4]
  assign regs_311_io_enable = 1'h1; // @[RegFile.scala 74:20:@38616.4]
  assign regs_312_clock = clock; // @[:@38625.4]
  assign regs_312_reset = io_reset; // @[:@38626.4 RegFile.scala 76:16:@38633.4]
  assign regs_312_io_in = 64'h0; // @[RegFile.scala 75:16:@38632.4]
  assign regs_312_io_reset = reset; // @[RegFile.scala 78:19:@38636.4]
  assign regs_312_io_enable = 1'h1; // @[RegFile.scala 74:20:@38630.4]
  assign regs_313_clock = clock; // @[:@38639.4]
  assign regs_313_reset = io_reset; // @[:@38640.4 RegFile.scala 76:16:@38647.4]
  assign regs_313_io_in = 64'h0; // @[RegFile.scala 75:16:@38646.4]
  assign regs_313_io_reset = reset; // @[RegFile.scala 78:19:@38650.4]
  assign regs_313_io_enable = 1'h1; // @[RegFile.scala 74:20:@38644.4]
  assign regs_314_clock = clock; // @[:@38653.4]
  assign regs_314_reset = io_reset; // @[:@38654.4 RegFile.scala 76:16:@38661.4]
  assign regs_314_io_in = 64'h0; // @[RegFile.scala 75:16:@38660.4]
  assign regs_314_io_reset = reset; // @[RegFile.scala 78:19:@38664.4]
  assign regs_314_io_enable = 1'h1; // @[RegFile.scala 74:20:@38658.4]
  assign regs_315_clock = clock; // @[:@38667.4]
  assign regs_315_reset = io_reset; // @[:@38668.4 RegFile.scala 76:16:@38675.4]
  assign regs_315_io_in = 64'h0; // @[RegFile.scala 75:16:@38674.4]
  assign regs_315_io_reset = reset; // @[RegFile.scala 78:19:@38678.4]
  assign regs_315_io_enable = 1'h1; // @[RegFile.scala 74:20:@38672.4]
  assign regs_316_clock = clock; // @[:@38681.4]
  assign regs_316_reset = io_reset; // @[:@38682.4 RegFile.scala 76:16:@38689.4]
  assign regs_316_io_in = 64'h0; // @[RegFile.scala 75:16:@38688.4]
  assign regs_316_io_reset = reset; // @[RegFile.scala 78:19:@38692.4]
  assign regs_316_io_enable = 1'h1; // @[RegFile.scala 74:20:@38686.4]
  assign regs_317_clock = clock; // @[:@38695.4]
  assign regs_317_reset = io_reset; // @[:@38696.4 RegFile.scala 76:16:@38703.4]
  assign regs_317_io_in = 64'h0; // @[RegFile.scala 75:16:@38702.4]
  assign regs_317_io_reset = reset; // @[RegFile.scala 78:19:@38706.4]
  assign regs_317_io_enable = 1'h1; // @[RegFile.scala 74:20:@38700.4]
  assign regs_318_clock = clock; // @[:@38709.4]
  assign regs_318_reset = io_reset; // @[:@38710.4 RegFile.scala 76:16:@38717.4]
  assign regs_318_io_in = 64'h0; // @[RegFile.scala 75:16:@38716.4]
  assign regs_318_io_reset = reset; // @[RegFile.scala 78:19:@38720.4]
  assign regs_318_io_enable = 1'h1; // @[RegFile.scala 74:20:@38714.4]
  assign regs_319_clock = clock; // @[:@38723.4]
  assign regs_319_reset = io_reset; // @[:@38724.4 RegFile.scala 76:16:@38731.4]
  assign regs_319_io_in = 64'h0; // @[RegFile.scala 75:16:@38730.4]
  assign regs_319_io_reset = reset; // @[RegFile.scala 78:19:@38734.4]
  assign regs_319_io_enable = 1'h1; // @[RegFile.scala 74:20:@38728.4]
  assign regs_320_clock = clock; // @[:@38737.4]
  assign regs_320_reset = io_reset; // @[:@38738.4 RegFile.scala 76:16:@38745.4]
  assign regs_320_io_in = 64'h0; // @[RegFile.scala 75:16:@38744.4]
  assign regs_320_io_reset = reset; // @[RegFile.scala 78:19:@38748.4]
  assign regs_320_io_enable = 1'h1; // @[RegFile.scala 74:20:@38742.4]
  assign regs_321_clock = clock; // @[:@38751.4]
  assign regs_321_reset = io_reset; // @[:@38752.4 RegFile.scala 76:16:@38759.4]
  assign regs_321_io_in = 64'h0; // @[RegFile.scala 75:16:@38758.4]
  assign regs_321_io_reset = reset; // @[RegFile.scala 78:19:@38762.4]
  assign regs_321_io_enable = 1'h1; // @[RegFile.scala 74:20:@38756.4]
  assign regs_322_clock = clock; // @[:@38765.4]
  assign regs_322_reset = io_reset; // @[:@38766.4 RegFile.scala 76:16:@38773.4]
  assign regs_322_io_in = 64'h0; // @[RegFile.scala 75:16:@38772.4]
  assign regs_322_io_reset = reset; // @[RegFile.scala 78:19:@38776.4]
  assign regs_322_io_enable = 1'h1; // @[RegFile.scala 74:20:@38770.4]
  assign regs_323_clock = clock; // @[:@38779.4]
  assign regs_323_reset = io_reset; // @[:@38780.4 RegFile.scala 76:16:@38787.4]
  assign regs_323_io_in = 64'h0; // @[RegFile.scala 75:16:@38786.4]
  assign regs_323_io_reset = reset; // @[RegFile.scala 78:19:@38790.4]
  assign regs_323_io_enable = 1'h1; // @[RegFile.scala 74:20:@38784.4]
  assign regs_324_clock = clock; // @[:@38793.4]
  assign regs_324_reset = io_reset; // @[:@38794.4 RegFile.scala 76:16:@38801.4]
  assign regs_324_io_in = 64'h0; // @[RegFile.scala 75:16:@38800.4]
  assign regs_324_io_reset = reset; // @[RegFile.scala 78:19:@38804.4]
  assign regs_324_io_enable = 1'h1; // @[RegFile.scala 74:20:@38798.4]
  assign regs_325_clock = clock; // @[:@38807.4]
  assign regs_325_reset = io_reset; // @[:@38808.4 RegFile.scala 76:16:@38815.4]
  assign regs_325_io_in = 64'h0; // @[RegFile.scala 75:16:@38814.4]
  assign regs_325_io_reset = reset; // @[RegFile.scala 78:19:@38818.4]
  assign regs_325_io_enable = 1'h1; // @[RegFile.scala 74:20:@38812.4]
  assign regs_326_clock = clock; // @[:@38821.4]
  assign regs_326_reset = io_reset; // @[:@38822.4 RegFile.scala 76:16:@38829.4]
  assign regs_326_io_in = 64'h0; // @[RegFile.scala 75:16:@38828.4]
  assign regs_326_io_reset = reset; // @[RegFile.scala 78:19:@38832.4]
  assign regs_326_io_enable = 1'h1; // @[RegFile.scala 74:20:@38826.4]
  assign regs_327_clock = clock; // @[:@38835.4]
  assign regs_327_reset = io_reset; // @[:@38836.4 RegFile.scala 76:16:@38843.4]
  assign regs_327_io_in = 64'h0; // @[RegFile.scala 75:16:@38842.4]
  assign regs_327_io_reset = reset; // @[RegFile.scala 78:19:@38846.4]
  assign regs_327_io_enable = 1'h1; // @[RegFile.scala 74:20:@38840.4]
  assign regs_328_clock = clock; // @[:@38849.4]
  assign regs_328_reset = io_reset; // @[:@38850.4 RegFile.scala 76:16:@38857.4]
  assign regs_328_io_in = 64'h0; // @[RegFile.scala 75:16:@38856.4]
  assign regs_328_io_reset = reset; // @[RegFile.scala 78:19:@38860.4]
  assign regs_328_io_enable = 1'h1; // @[RegFile.scala 74:20:@38854.4]
  assign regs_329_clock = clock; // @[:@38863.4]
  assign regs_329_reset = io_reset; // @[:@38864.4 RegFile.scala 76:16:@38871.4]
  assign regs_329_io_in = 64'h0; // @[RegFile.scala 75:16:@38870.4]
  assign regs_329_io_reset = reset; // @[RegFile.scala 78:19:@38874.4]
  assign regs_329_io_enable = 1'h1; // @[RegFile.scala 74:20:@38868.4]
  assign regs_330_clock = clock; // @[:@38877.4]
  assign regs_330_reset = io_reset; // @[:@38878.4 RegFile.scala 76:16:@38885.4]
  assign regs_330_io_in = 64'h0; // @[RegFile.scala 75:16:@38884.4]
  assign regs_330_io_reset = reset; // @[RegFile.scala 78:19:@38888.4]
  assign regs_330_io_enable = 1'h1; // @[RegFile.scala 74:20:@38882.4]
  assign regs_331_clock = clock; // @[:@38891.4]
  assign regs_331_reset = io_reset; // @[:@38892.4 RegFile.scala 76:16:@38899.4]
  assign regs_331_io_in = 64'h0; // @[RegFile.scala 75:16:@38898.4]
  assign regs_331_io_reset = reset; // @[RegFile.scala 78:19:@38902.4]
  assign regs_331_io_enable = 1'h1; // @[RegFile.scala 74:20:@38896.4]
  assign regs_332_clock = clock; // @[:@38905.4]
  assign regs_332_reset = io_reset; // @[:@38906.4 RegFile.scala 76:16:@38913.4]
  assign regs_332_io_in = 64'h0; // @[RegFile.scala 75:16:@38912.4]
  assign regs_332_io_reset = reset; // @[RegFile.scala 78:19:@38916.4]
  assign regs_332_io_enable = 1'h1; // @[RegFile.scala 74:20:@38910.4]
  assign regs_333_clock = clock; // @[:@38919.4]
  assign regs_333_reset = io_reset; // @[:@38920.4 RegFile.scala 76:16:@38927.4]
  assign regs_333_io_in = 64'h0; // @[RegFile.scala 75:16:@38926.4]
  assign regs_333_io_reset = reset; // @[RegFile.scala 78:19:@38930.4]
  assign regs_333_io_enable = 1'h1; // @[RegFile.scala 74:20:@38924.4]
  assign regs_334_clock = clock; // @[:@38933.4]
  assign regs_334_reset = io_reset; // @[:@38934.4 RegFile.scala 76:16:@38941.4]
  assign regs_334_io_in = 64'h0; // @[RegFile.scala 75:16:@38940.4]
  assign regs_334_io_reset = reset; // @[RegFile.scala 78:19:@38944.4]
  assign regs_334_io_enable = 1'h1; // @[RegFile.scala 74:20:@38938.4]
  assign regs_335_clock = clock; // @[:@38947.4]
  assign regs_335_reset = io_reset; // @[:@38948.4 RegFile.scala 76:16:@38955.4]
  assign regs_335_io_in = 64'h0; // @[RegFile.scala 75:16:@38954.4]
  assign regs_335_io_reset = reset; // @[RegFile.scala 78:19:@38958.4]
  assign regs_335_io_enable = 1'h1; // @[RegFile.scala 74:20:@38952.4]
  assign regs_336_clock = clock; // @[:@38961.4]
  assign regs_336_reset = io_reset; // @[:@38962.4 RegFile.scala 76:16:@38969.4]
  assign regs_336_io_in = 64'h0; // @[RegFile.scala 75:16:@38968.4]
  assign regs_336_io_reset = reset; // @[RegFile.scala 78:19:@38972.4]
  assign regs_336_io_enable = 1'h1; // @[RegFile.scala 74:20:@38966.4]
  assign regs_337_clock = clock; // @[:@38975.4]
  assign regs_337_reset = io_reset; // @[:@38976.4 RegFile.scala 76:16:@38983.4]
  assign regs_337_io_in = 64'h0; // @[RegFile.scala 75:16:@38982.4]
  assign regs_337_io_reset = reset; // @[RegFile.scala 78:19:@38986.4]
  assign regs_337_io_enable = 1'h1; // @[RegFile.scala 74:20:@38980.4]
  assign regs_338_clock = clock; // @[:@38989.4]
  assign regs_338_reset = io_reset; // @[:@38990.4 RegFile.scala 76:16:@38997.4]
  assign regs_338_io_in = 64'h0; // @[RegFile.scala 75:16:@38996.4]
  assign regs_338_io_reset = reset; // @[RegFile.scala 78:19:@39000.4]
  assign regs_338_io_enable = 1'h1; // @[RegFile.scala 74:20:@38994.4]
  assign regs_339_clock = clock; // @[:@39003.4]
  assign regs_339_reset = io_reset; // @[:@39004.4 RegFile.scala 76:16:@39011.4]
  assign regs_339_io_in = 64'h0; // @[RegFile.scala 75:16:@39010.4]
  assign regs_339_io_reset = reset; // @[RegFile.scala 78:19:@39014.4]
  assign regs_339_io_enable = 1'h1; // @[RegFile.scala 74:20:@39008.4]
  assign regs_340_clock = clock; // @[:@39017.4]
  assign regs_340_reset = io_reset; // @[:@39018.4 RegFile.scala 76:16:@39025.4]
  assign regs_340_io_in = 64'h0; // @[RegFile.scala 75:16:@39024.4]
  assign regs_340_io_reset = reset; // @[RegFile.scala 78:19:@39028.4]
  assign regs_340_io_enable = 1'h1; // @[RegFile.scala 74:20:@39022.4]
  assign regs_341_clock = clock; // @[:@39031.4]
  assign regs_341_reset = io_reset; // @[:@39032.4 RegFile.scala 76:16:@39039.4]
  assign regs_341_io_in = 64'h0; // @[RegFile.scala 75:16:@39038.4]
  assign regs_341_io_reset = reset; // @[RegFile.scala 78:19:@39042.4]
  assign regs_341_io_enable = 1'h1; // @[RegFile.scala 74:20:@39036.4]
  assign regs_342_clock = clock; // @[:@39045.4]
  assign regs_342_reset = io_reset; // @[:@39046.4 RegFile.scala 76:16:@39053.4]
  assign regs_342_io_in = 64'h0; // @[RegFile.scala 75:16:@39052.4]
  assign regs_342_io_reset = reset; // @[RegFile.scala 78:19:@39056.4]
  assign regs_342_io_enable = 1'h1; // @[RegFile.scala 74:20:@39050.4]
  assign regs_343_clock = clock; // @[:@39059.4]
  assign regs_343_reset = io_reset; // @[:@39060.4 RegFile.scala 76:16:@39067.4]
  assign regs_343_io_in = 64'h0; // @[RegFile.scala 75:16:@39066.4]
  assign regs_343_io_reset = reset; // @[RegFile.scala 78:19:@39070.4]
  assign regs_343_io_enable = 1'h1; // @[RegFile.scala 74:20:@39064.4]
  assign regs_344_clock = clock; // @[:@39073.4]
  assign regs_344_reset = io_reset; // @[:@39074.4 RegFile.scala 76:16:@39081.4]
  assign regs_344_io_in = 64'h0; // @[RegFile.scala 75:16:@39080.4]
  assign regs_344_io_reset = reset; // @[RegFile.scala 78:19:@39084.4]
  assign regs_344_io_enable = 1'h1; // @[RegFile.scala 74:20:@39078.4]
  assign regs_345_clock = clock; // @[:@39087.4]
  assign regs_345_reset = io_reset; // @[:@39088.4 RegFile.scala 76:16:@39095.4]
  assign regs_345_io_in = 64'h0; // @[RegFile.scala 75:16:@39094.4]
  assign regs_345_io_reset = reset; // @[RegFile.scala 78:19:@39098.4]
  assign regs_345_io_enable = 1'h1; // @[RegFile.scala 74:20:@39092.4]
  assign regs_346_clock = clock; // @[:@39101.4]
  assign regs_346_reset = io_reset; // @[:@39102.4 RegFile.scala 76:16:@39109.4]
  assign regs_346_io_in = 64'h0; // @[RegFile.scala 75:16:@39108.4]
  assign regs_346_io_reset = reset; // @[RegFile.scala 78:19:@39112.4]
  assign regs_346_io_enable = 1'h1; // @[RegFile.scala 74:20:@39106.4]
  assign regs_347_clock = clock; // @[:@39115.4]
  assign regs_347_reset = io_reset; // @[:@39116.4 RegFile.scala 76:16:@39123.4]
  assign regs_347_io_in = 64'h0; // @[RegFile.scala 75:16:@39122.4]
  assign regs_347_io_reset = reset; // @[RegFile.scala 78:19:@39126.4]
  assign regs_347_io_enable = 1'h1; // @[RegFile.scala 74:20:@39120.4]
  assign regs_348_clock = clock; // @[:@39129.4]
  assign regs_348_reset = io_reset; // @[:@39130.4 RegFile.scala 76:16:@39137.4]
  assign regs_348_io_in = 64'h0; // @[RegFile.scala 75:16:@39136.4]
  assign regs_348_io_reset = reset; // @[RegFile.scala 78:19:@39140.4]
  assign regs_348_io_enable = 1'h1; // @[RegFile.scala 74:20:@39134.4]
  assign regs_349_clock = clock; // @[:@39143.4]
  assign regs_349_reset = io_reset; // @[:@39144.4 RegFile.scala 76:16:@39151.4]
  assign regs_349_io_in = 64'h0; // @[RegFile.scala 75:16:@39150.4]
  assign regs_349_io_reset = reset; // @[RegFile.scala 78:19:@39154.4]
  assign regs_349_io_enable = 1'h1; // @[RegFile.scala 74:20:@39148.4]
  assign regs_350_clock = clock; // @[:@39157.4]
  assign regs_350_reset = io_reset; // @[:@39158.4 RegFile.scala 76:16:@39165.4]
  assign regs_350_io_in = 64'h0; // @[RegFile.scala 75:16:@39164.4]
  assign regs_350_io_reset = reset; // @[RegFile.scala 78:19:@39168.4]
  assign regs_350_io_enable = 1'h1; // @[RegFile.scala 74:20:@39162.4]
  assign regs_351_clock = clock; // @[:@39171.4]
  assign regs_351_reset = io_reset; // @[:@39172.4 RegFile.scala 76:16:@39179.4]
  assign regs_351_io_in = 64'h0; // @[RegFile.scala 75:16:@39178.4]
  assign regs_351_io_reset = reset; // @[RegFile.scala 78:19:@39182.4]
  assign regs_351_io_enable = 1'h1; // @[RegFile.scala 74:20:@39176.4]
  assign regs_352_clock = clock; // @[:@39185.4]
  assign regs_352_reset = io_reset; // @[:@39186.4 RegFile.scala 76:16:@39193.4]
  assign regs_352_io_in = 64'h0; // @[RegFile.scala 75:16:@39192.4]
  assign regs_352_io_reset = reset; // @[RegFile.scala 78:19:@39196.4]
  assign regs_352_io_enable = 1'h1; // @[RegFile.scala 74:20:@39190.4]
  assign regs_353_clock = clock; // @[:@39199.4]
  assign regs_353_reset = io_reset; // @[:@39200.4 RegFile.scala 76:16:@39207.4]
  assign regs_353_io_in = 64'h0; // @[RegFile.scala 75:16:@39206.4]
  assign regs_353_io_reset = reset; // @[RegFile.scala 78:19:@39210.4]
  assign regs_353_io_enable = 1'h1; // @[RegFile.scala 74:20:@39204.4]
  assign regs_354_clock = clock; // @[:@39213.4]
  assign regs_354_reset = io_reset; // @[:@39214.4 RegFile.scala 76:16:@39221.4]
  assign regs_354_io_in = 64'h0; // @[RegFile.scala 75:16:@39220.4]
  assign regs_354_io_reset = reset; // @[RegFile.scala 78:19:@39224.4]
  assign regs_354_io_enable = 1'h1; // @[RegFile.scala 74:20:@39218.4]
  assign regs_355_clock = clock; // @[:@39227.4]
  assign regs_355_reset = io_reset; // @[:@39228.4 RegFile.scala 76:16:@39235.4]
  assign regs_355_io_in = 64'h0; // @[RegFile.scala 75:16:@39234.4]
  assign regs_355_io_reset = reset; // @[RegFile.scala 78:19:@39238.4]
  assign regs_355_io_enable = 1'h1; // @[RegFile.scala 74:20:@39232.4]
  assign regs_356_clock = clock; // @[:@39241.4]
  assign regs_356_reset = io_reset; // @[:@39242.4 RegFile.scala 76:16:@39249.4]
  assign regs_356_io_in = 64'h0; // @[RegFile.scala 75:16:@39248.4]
  assign regs_356_io_reset = reset; // @[RegFile.scala 78:19:@39252.4]
  assign regs_356_io_enable = 1'h1; // @[RegFile.scala 74:20:@39246.4]
  assign regs_357_clock = clock; // @[:@39255.4]
  assign regs_357_reset = io_reset; // @[:@39256.4 RegFile.scala 76:16:@39263.4]
  assign regs_357_io_in = 64'h0; // @[RegFile.scala 75:16:@39262.4]
  assign regs_357_io_reset = reset; // @[RegFile.scala 78:19:@39266.4]
  assign regs_357_io_enable = 1'h1; // @[RegFile.scala 74:20:@39260.4]
  assign regs_358_clock = clock; // @[:@39269.4]
  assign regs_358_reset = io_reset; // @[:@39270.4 RegFile.scala 76:16:@39277.4]
  assign regs_358_io_in = 64'h0; // @[RegFile.scala 75:16:@39276.4]
  assign regs_358_io_reset = reset; // @[RegFile.scala 78:19:@39280.4]
  assign regs_358_io_enable = 1'h1; // @[RegFile.scala 74:20:@39274.4]
  assign regs_359_clock = clock; // @[:@39283.4]
  assign regs_359_reset = io_reset; // @[:@39284.4 RegFile.scala 76:16:@39291.4]
  assign regs_359_io_in = 64'h0; // @[RegFile.scala 75:16:@39290.4]
  assign regs_359_io_reset = reset; // @[RegFile.scala 78:19:@39294.4]
  assign regs_359_io_enable = 1'h1; // @[RegFile.scala 74:20:@39288.4]
  assign regs_360_clock = clock; // @[:@39297.4]
  assign regs_360_reset = io_reset; // @[:@39298.4 RegFile.scala 76:16:@39305.4]
  assign regs_360_io_in = 64'h0; // @[RegFile.scala 75:16:@39304.4]
  assign regs_360_io_reset = reset; // @[RegFile.scala 78:19:@39308.4]
  assign regs_360_io_enable = 1'h1; // @[RegFile.scala 74:20:@39302.4]
  assign regs_361_clock = clock; // @[:@39311.4]
  assign regs_361_reset = io_reset; // @[:@39312.4 RegFile.scala 76:16:@39319.4]
  assign regs_361_io_in = 64'h0; // @[RegFile.scala 75:16:@39318.4]
  assign regs_361_io_reset = reset; // @[RegFile.scala 78:19:@39322.4]
  assign regs_361_io_enable = 1'h1; // @[RegFile.scala 74:20:@39316.4]
  assign regs_362_clock = clock; // @[:@39325.4]
  assign regs_362_reset = io_reset; // @[:@39326.4 RegFile.scala 76:16:@39333.4]
  assign regs_362_io_in = 64'h0; // @[RegFile.scala 75:16:@39332.4]
  assign regs_362_io_reset = reset; // @[RegFile.scala 78:19:@39336.4]
  assign regs_362_io_enable = 1'h1; // @[RegFile.scala 74:20:@39330.4]
  assign regs_363_clock = clock; // @[:@39339.4]
  assign regs_363_reset = io_reset; // @[:@39340.4 RegFile.scala 76:16:@39347.4]
  assign regs_363_io_in = 64'h0; // @[RegFile.scala 75:16:@39346.4]
  assign regs_363_io_reset = reset; // @[RegFile.scala 78:19:@39350.4]
  assign regs_363_io_enable = 1'h1; // @[RegFile.scala 74:20:@39344.4]
  assign regs_364_clock = clock; // @[:@39353.4]
  assign regs_364_reset = io_reset; // @[:@39354.4 RegFile.scala 76:16:@39361.4]
  assign regs_364_io_in = 64'h0; // @[RegFile.scala 75:16:@39360.4]
  assign regs_364_io_reset = reset; // @[RegFile.scala 78:19:@39364.4]
  assign regs_364_io_enable = 1'h1; // @[RegFile.scala 74:20:@39358.4]
  assign regs_365_clock = clock; // @[:@39367.4]
  assign regs_365_reset = io_reset; // @[:@39368.4 RegFile.scala 76:16:@39375.4]
  assign regs_365_io_in = 64'h0; // @[RegFile.scala 75:16:@39374.4]
  assign regs_365_io_reset = reset; // @[RegFile.scala 78:19:@39378.4]
  assign regs_365_io_enable = 1'h1; // @[RegFile.scala 74:20:@39372.4]
  assign regs_366_clock = clock; // @[:@39381.4]
  assign regs_366_reset = io_reset; // @[:@39382.4 RegFile.scala 76:16:@39389.4]
  assign regs_366_io_in = 64'h0; // @[RegFile.scala 75:16:@39388.4]
  assign regs_366_io_reset = reset; // @[RegFile.scala 78:19:@39392.4]
  assign regs_366_io_enable = 1'h1; // @[RegFile.scala 74:20:@39386.4]
  assign regs_367_clock = clock; // @[:@39395.4]
  assign regs_367_reset = io_reset; // @[:@39396.4 RegFile.scala 76:16:@39403.4]
  assign regs_367_io_in = 64'h0; // @[RegFile.scala 75:16:@39402.4]
  assign regs_367_io_reset = reset; // @[RegFile.scala 78:19:@39406.4]
  assign regs_367_io_enable = 1'h1; // @[RegFile.scala 74:20:@39400.4]
  assign regs_368_clock = clock; // @[:@39409.4]
  assign regs_368_reset = io_reset; // @[:@39410.4 RegFile.scala 76:16:@39417.4]
  assign regs_368_io_in = 64'h0; // @[RegFile.scala 75:16:@39416.4]
  assign regs_368_io_reset = reset; // @[RegFile.scala 78:19:@39420.4]
  assign regs_368_io_enable = 1'h1; // @[RegFile.scala 74:20:@39414.4]
  assign regs_369_clock = clock; // @[:@39423.4]
  assign regs_369_reset = io_reset; // @[:@39424.4 RegFile.scala 76:16:@39431.4]
  assign regs_369_io_in = 64'h0; // @[RegFile.scala 75:16:@39430.4]
  assign regs_369_io_reset = reset; // @[RegFile.scala 78:19:@39434.4]
  assign regs_369_io_enable = 1'h1; // @[RegFile.scala 74:20:@39428.4]
  assign regs_370_clock = clock; // @[:@39437.4]
  assign regs_370_reset = io_reset; // @[:@39438.4 RegFile.scala 76:16:@39445.4]
  assign regs_370_io_in = 64'h0; // @[RegFile.scala 75:16:@39444.4]
  assign regs_370_io_reset = reset; // @[RegFile.scala 78:19:@39448.4]
  assign regs_370_io_enable = 1'h1; // @[RegFile.scala 74:20:@39442.4]
  assign regs_371_clock = clock; // @[:@39451.4]
  assign regs_371_reset = io_reset; // @[:@39452.4 RegFile.scala 76:16:@39459.4]
  assign regs_371_io_in = 64'h0; // @[RegFile.scala 75:16:@39458.4]
  assign regs_371_io_reset = reset; // @[RegFile.scala 78:19:@39462.4]
  assign regs_371_io_enable = 1'h1; // @[RegFile.scala 74:20:@39456.4]
  assign regs_372_clock = clock; // @[:@39465.4]
  assign regs_372_reset = io_reset; // @[:@39466.4 RegFile.scala 76:16:@39473.4]
  assign regs_372_io_in = 64'h0; // @[RegFile.scala 75:16:@39472.4]
  assign regs_372_io_reset = reset; // @[RegFile.scala 78:19:@39476.4]
  assign regs_372_io_enable = 1'h1; // @[RegFile.scala 74:20:@39470.4]
  assign regs_373_clock = clock; // @[:@39479.4]
  assign regs_373_reset = io_reset; // @[:@39480.4 RegFile.scala 76:16:@39487.4]
  assign regs_373_io_in = 64'h0; // @[RegFile.scala 75:16:@39486.4]
  assign regs_373_io_reset = reset; // @[RegFile.scala 78:19:@39490.4]
  assign regs_373_io_enable = 1'h1; // @[RegFile.scala 74:20:@39484.4]
  assign regs_374_clock = clock; // @[:@39493.4]
  assign regs_374_reset = io_reset; // @[:@39494.4 RegFile.scala 76:16:@39501.4]
  assign regs_374_io_in = 64'h0; // @[RegFile.scala 75:16:@39500.4]
  assign regs_374_io_reset = reset; // @[RegFile.scala 78:19:@39504.4]
  assign regs_374_io_enable = 1'h1; // @[RegFile.scala 74:20:@39498.4]
  assign regs_375_clock = clock; // @[:@39507.4]
  assign regs_375_reset = io_reset; // @[:@39508.4 RegFile.scala 76:16:@39515.4]
  assign regs_375_io_in = 64'h0; // @[RegFile.scala 75:16:@39514.4]
  assign regs_375_io_reset = reset; // @[RegFile.scala 78:19:@39518.4]
  assign regs_375_io_enable = 1'h1; // @[RegFile.scala 74:20:@39512.4]
  assign regs_376_clock = clock; // @[:@39521.4]
  assign regs_376_reset = io_reset; // @[:@39522.4 RegFile.scala 76:16:@39529.4]
  assign regs_376_io_in = 64'h0; // @[RegFile.scala 75:16:@39528.4]
  assign regs_376_io_reset = reset; // @[RegFile.scala 78:19:@39532.4]
  assign regs_376_io_enable = 1'h1; // @[RegFile.scala 74:20:@39526.4]
  assign regs_377_clock = clock; // @[:@39535.4]
  assign regs_377_reset = io_reset; // @[:@39536.4 RegFile.scala 76:16:@39543.4]
  assign regs_377_io_in = 64'h0; // @[RegFile.scala 75:16:@39542.4]
  assign regs_377_io_reset = reset; // @[RegFile.scala 78:19:@39546.4]
  assign regs_377_io_enable = 1'h1; // @[RegFile.scala 74:20:@39540.4]
  assign regs_378_clock = clock; // @[:@39549.4]
  assign regs_378_reset = io_reset; // @[:@39550.4 RegFile.scala 76:16:@39557.4]
  assign regs_378_io_in = 64'h0; // @[RegFile.scala 75:16:@39556.4]
  assign regs_378_io_reset = reset; // @[RegFile.scala 78:19:@39560.4]
  assign regs_378_io_enable = 1'h1; // @[RegFile.scala 74:20:@39554.4]
  assign regs_379_clock = clock; // @[:@39563.4]
  assign regs_379_reset = io_reset; // @[:@39564.4 RegFile.scala 76:16:@39571.4]
  assign regs_379_io_in = 64'h0; // @[RegFile.scala 75:16:@39570.4]
  assign regs_379_io_reset = reset; // @[RegFile.scala 78:19:@39574.4]
  assign regs_379_io_enable = 1'h1; // @[RegFile.scala 74:20:@39568.4]
  assign regs_380_clock = clock; // @[:@39577.4]
  assign regs_380_reset = io_reset; // @[:@39578.4 RegFile.scala 76:16:@39585.4]
  assign regs_380_io_in = 64'h0; // @[RegFile.scala 75:16:@39584.4]
  assign regs_380_io_reset = reset; // @[RegFile.scala 78:19:@39588.4]
  assign regs_380_io_enable = 1'h1; // @[RegFile.scala 74:20:@39582.4]
  assign regs_381_clock = clock; // @[:@39591.4]
  assign regs_381_reset = io_reset; // @[:@39592.4 RegFile.scala 76:16:@39599.4]
  assign regs_381_io_in = 64'h0; // @[RegFile.scala 75:16:@39598.4]
  assign regs_381_io_reset = reset; // @[RegFile.scala 78:19:@39602.4]
  assign regs_381_io_enable = 1'h1; // @[RegFile.scala 74:20:@39596.4]
  assign regs_382_clock = clock; // @[:@39605.4]
  assign regs_382_reset = io_reset; // @[:@39606.4 RegFile.scala 76:16:@39613.4]
  assign regs_382_io_in = 64'h0; // @[RegFile.scala 75:16:@39612.4]
  assign regs_382_io_reset = reset; // @[RegFile.scala 78:19:@39616.4]
  assign regs_382_io_enable = 1'h1; // @[RegFile.scala 74:20:@39610.4]
  assign regs_383_clock = clock; // @[:@39619.4]
  assign regs_383_reset = io_reset; // @[:@39620.4 RegFile.scala 76:16:@39627.4]
  assign regs_383_io_in = 64'h0; // @[RegFile.scala 75:16:@39626.4]
  assign regs_383_io_reset = reset; // @[RegFile.scala 78:19:@39630.4]
  assign regs_383_io_enable = 1'h1; // @[RegFile.scala 74:20:@39624.4]
  assign regs_384_clock = clock; // @[:@39633.4]
  assign regs_384_reset = io_reset; // @[:@39634.4 RegFile.scala 76:16:@39641.4]
  assign regs_384_io_in = 64'h0; // @[RegFile.scala 75:16:@39640.4]
  assign regs_384_io_reset = reset; // @[RegFile.scala 78:19:@39644.4]
  assign regs_384_io_enable = 1'h1; // @[RegFile.scala 74:20:@39638.4]
  assign regs_385_clock = clock; // @[:@39647.4]
  assign regs_385_reset = io_reset; // @[:@39648.4 RegFile.scala 76:16:@39655.4]
  assign regs_385_io_in = 64'h0; // @[RegFile.scala 75:16:@39654.4]
  assign regs_385_io_reset = reset; // @[RegFile.scala 78:19:@39658.4]
  assign regs_385_io_enable = 1'h1; // @[RegFile.scala 74:20:@39652.4]
  assign regs_386_clock = clock; // @[:@39661.4]
  assign regs_386_reset = io_reset; // @[:@39662.4 RegFile.scala 76:16:@39669.4]
  assign regs_386_io_in = 64'h0; // @[RegFile.scala 75:16:@39668.4]
  assign regs_386_io_reset = reset; // @[RegFile.scala 78:19:@39672.4]
  assign regs_386_io_enable = 1'h1; // @[RegFile.scala 74:20:@39666.4]
  assign regs_387_clock = clock; // @[:@39675.4]
  assign regs_387_reset = io_reset; // @[:@39676.4 RegFile.scala 76:16:@39683.4]
  assign regs_387_io_in = 64'h0; // @[RegFile.scala 75:16:@39682.4]
  assign regs_387_io_reset = reset; // @[RegFile.scala 78:19:@39686.4]
  assign regs_387_io_enable = 1'h1; // @[RegFile.scala 74:20:@39680.4]
  assign regs_388_clock = clock; // @[:@39689.4]
  assign regs_388_reset = io_reset; // @[:@39690.4 RegFile.scala 76:16:@39697.4]
  assign regs_388_io_in = 64'h0; // @[RegFile.scala 75:16:@39696.4]
  assign regs_388_io_reset = reset; // @[RegFile.scala 78:19:@39700.4]
  assign regs_388_io_enable = 1'h1; // @[RegFile.scala 74:20:@39694.4]
  assign regs_389_clock = clock; // @[:@39703.4]
  assign regs_389_reset = io_reset; // @[:@39704.4 RegFile.scala 76:16:@39711.4]
  assign regs_389_io_in = 64'h0; // @[RegFile.scala 75:16:@39710.4]
  assign regs_389_io_reset = reset; // @[RegFile.scala 78:19:@39714.4]
  assign regs_389_io_enable = 1'h1; // @[RegFile.scala 74:20:@39708.4]
  assign regs_390_clock = clock; // @[:@39717.4]
  assign regs_390_reset = io_reset; // @[:@39718.4 RegFile.scala 76:16:@39725.4]
  assign regs_390_io_in = 64'h0; // @[RegFile.scala 75:16:@39724.4]
  assign regs_390_io_reset = reset; // @[RegFile.scala 78:19:@39728.4]
  assign regs_390_io_enable = 1'h1; // @[RegFile.scala 74:20:@39722.4]
  assign regs_391_clock = clock; // @[:@39731.4]
  assign regs_391_reset = io_reset; // @[:@39732.4 RegFile.scala 76:16:@39739.4]
  assign regs_391_io_in = 64'h0; // @[RegFile.scala 75:16:@39738.4]
  assign regs_391_io_reset = reset; // @[RegFile.scala 78:19:@39742.4]
  assign regs_391_io_enable = 1'h1; // @[RegFile.scala 74:20:@39736.4]
  assign regs_392_clock = clock; // @[:@39745.4]
  assign regs_392_reset = io_reset; // @[:@39746.4 RegFile.scala 76:16:@39753.4]
  assign regs_392_io_in = 64'h0; // @[RegFile.scala 75:16:@39752.4]
  assign regs_392_io_reset = reset; // @[RegFile.scala 78:19:@39756.4]
  assign regs_392_io_enable = 1'h1; // @[RegFile.scala 74:20:@39750.4]
  assign regs_393_clock = clock; // @[:@39759.4]
  assign regs_393_reset = io_reset; // @[:@39760.4 RegFile.scala 76:16:@39767.4]
  assign regs_393_io_in = 64'h0; // @[RegFile.scala 75:16:@39766.4]
  assign regs_393_io_reset = reset; // @[RegFile.scala 78:19:@39770.4]
  assign regs_393_io_enable = 1'h1; // @[RegFile.scala 74:20:@39764.4]
  assign regs_394_clock = clock; // @[:@39773.4]
  assign regs_394_reset = io_reset; // @[:@39774.4 RegFile.scala 76:16:@39781.4]
  assign regs_394_io_in = 64'h0; // @[RegFile.scala 75:16:@39780.4]
  assign regs_394_io_reset = reset; // @[RegFile.scala 78:19:@39784.4]
  assign regs_394_io_enable = 1'h1; // @[RegFile.scala 74:20:@39778.4]
  assign regs_395_clock = clock; // @[:@39787.4]
  assign regs_395_reset = io_reset; // @[:@39788.4 RegFile.scala 76:16:@39795.4]
  assign regs_395_io_in = 64'h0; // @[RegFile.scala 75:16:@39794.4]
  assign regs_395_io_reset = reset; // @[RegFile.scala 78:19:@39798.4]
  assign regs_395_io_enable = 1'h1; // @[RegFile.scala 74:20:@39792.4]
  assign regs_396_clock = clock; // @[:@39801.4]
  assign regs_396_reset = io_reset; // @[:@39802.4 RegFile.scala 76:16:@39809.4]
  assign regs_396_io_in = 64'h0; // @[RegFile.scala 75:16:@39808.4]
  assign regs_396_io_reset = reset; // @[RegFile.scala 78:19:@39812.4]
  assign regs_396_io_enable = 1'h1; // @[RegFile.scala 74:20:@39806.4]
  assign regs_397_clock = clock; // @[:@39815.4]
  assign regs_397_reset = io_reset; // @[:@39816.4 RegFile.scala 76:16:@39823.4]
  assign regs_397_io_in = 64'h0; // @[RegFile.scala 75:16:@39822.4]
  assign regs_397_io_reset = reset; // @[RegFile.scala 78:19:@39826.4]
  assign regs_397_io_enable = 1'h1; // @[RegFile.scala 74:20:@39820.4]
  assign regs_398_clock = clock; // @[:@39829.4]
  assign regs_398_reset = io_reset; // @[:@39830.4 RegFile.scala 76:16:@39837.4]
  assign regs_398_io_in = 64'h0; // @[RegFile.scala 75:16:@39836.4]
  assign regs_398_io_reset = reset; // @[RegFile.scala 78:19:@39840.4]
  assign regs_398_io_enable = 1'h1; // @[RegFile.scala 74:20:@39834.4]
  assign regs_399_clock = clock; // @[:@39843.4]
  assign regs_399_reset = io_reset; // @[:@39844.4 RegFile.scala 76:16:@39851.4]
  assign regs_399_io_in = 64'h0; // @[RegFile.scala 75:16:@39850.4]
  assign regs_399_io_reset = reset; // @[RegFile.scala 78:19:@39854.4]
  assign regs_399_io_enable = 1'h1; // @[RegFile.scala 74:20:@39848.4]
  assign regs_400_clock = clock; // @[:@39857.4]
  assign regs_400_reset = io_reset; // @[:@39858.4 RegFile.scala 76:16:@39865.4]
  assign regs_400_io_in = 64'h0; // @[RegFile.scala 75:16:@39864.4]
  assign regs_400_io_reset = reset; // @[RegFile.scala 78:19:@39868.4]
  assign regs_400_io_enable = 1'h1; // @[RegFile.scala 74:20:@39862.4]
  assign regs_401_clock = clock; // @[:@39871.4]
  assign regs_401_reset = io_reset; // @[:@39872.4 RegFile.scala 76:16:@39879.4]
  assign regs_401_io_in = 64'h0; // @[RegFile.scala 75:16:@39878.4]
  assign regs_401_io_reset = reset; // @[RegFile.scala 78:19:@39882.4]
  assign regs_401_io_enable = 1'h1; // @[RegFile.scala 74:20:@39876.4]
  assign regs_402_clock = clock; // @[:@39885.4]
  assign regs_402_reset = io_reset; // @[:@39886.4 RegFile.scala 76:16:@39893.4]
  assign regs_402_io_in = 64'h0; // @[RegFile.scala 75:16:@39892.4]
  assign regs_402_io_reset = reset; // @[RegFile.scala 78:19:@39896.4]
  assign regs_402_io_enable = 1'h1; // @[RegFile.scala 74:20:@39890.4]
  assign regs_403_clock = clock; // @[:@39899.4]
  assign regs_403_reset = io_reset; // @[:@39900.4 RegFile.scala 76:16:@39907.4]
  assign regs_403_io_in = 64'h0; // @[RegFile.scala 75:16:@39906.4]
  assign regs_403_io_reset = reset; // @[RegFile.scala 78:19:@39910.4]
  assign regs_403_io_enable = 1'h1; // @[RegFile.scala 74:20:@39904.4]
  assign regs_404_clock = clock; // @[:@39913.4]
  assign regs_404_reset = io_reset; // @[:@39914.4 RegFile.scala 76:16:@39921.4]
  assign regs_404_io_in = 64'h0; // @[RegFile.scala 75:16:@39920.4]
  assign regs_404_io_reset = reset; // @[RegFile.scala 78:19:@39924.4]
  assign regs_404_io_enable = 1'h1; // @[RegFile.scala 74:20:@39918.4]
  assign regs_405_clock = clock; // @[:@39927.4]
  assign regs_405_reset = io_reset; // @[:@39928.4 RegFile.scala 76:16:@39935.4]
  assign regs_405_io_in = 64'h0; // @[RegFile.scala 75:16:@39934.4]
  assign regs_405_io_reset = reset; // @[RegFile.scala 78:19:@39938.4]
  assign regs_405_io_enable = 1'h1; // @[RegFile.scala 74:20:@39932.4]
  assign regs_406_clock = clock; // @[:@39941.4]
  assign regs_406_reset = io_reset; // @[:@39942.4 RegFile.scala 76:16:@39949.4]
  assign regs_406_io_in = 64'h0; // @[RegFile.scala 75:16:@39948.4]
  assign regs_406_io_reset = reset; // @[RegFile.scala 78:19:@39952.4]
  assign regs_406_io_enable = 1'h1; // @[RegFile.scala 74:20:@39946.4]
  assign regs_407_clock = clock; // @[:@39955.4]
  assign regs_407_reset = io_reset; // @[:@39956.4 RegFile.scala 76:16:@39963.4]
  assign regs_407_io_in = 64'h0; // @[RegFile.scala 75:16:@39962.4]
  assign regs_407_io_reset = reset; // @[RegFile.scala 78:19:@39966.4]
  assign regs_407_io_enable = 1'h1; // @[RegFile.scala 74:20:@39960.4]
  assign regs_408_clock = clock; // @[:@39969.4]
  assign regs_408_reset = io_reset; // @[:@39970.4 RegFile.scala 76:16:@39977.4]
  assign regs_408_io_in = 64'h0; // @[RegFile.scala 75:16:@39976.4]
  assign regs_408_io_reset = reset; // @[RegFile.scala 78:19:@39980.4]
  assign regs_408_io_enable = 1'h1; // @[RegFile.scala 74:20:@39974.4]
  assign regs_409_clock = clock; // @[:@39983.4]
  assign regs_409_reset = io_reset; // @[:@39984.4 RegFile.scala 76:16:@39991.4]
  assign regs_409_io_in = 64'h0; // @[RegFile.scala 75:16:@39990.4]
  assign regs_409_io_reset = reset; // @[RegFile.scala 78:19:@39994.4]
  assign regs_409_io_enable = 1'h1; // @[RegFile.scala 74:20:@39988.4]
  assign regs_410_clock = clock; // @[:@39997.4]
  assign regs_410_reset = io_reset; // @[:@39998.4 RegFile.scala 76:16:@40005.4]
  assign regs_410_io_in = 64'h0; // @[RegFile.scala 75:16:@40004.4]
  assign regs_410_io_reset = reset; // @[RegFile.scala 78:19:@40008.4]
  assign regs_410_io_enable = 1'h1; // @[RegFile.scala 74:20:@40002.4]
  assign regs_411_clock = clock; // @[:@40011.4]
  assign regs_411_reset = io_reset; // @[:@40012.4 RegFile.scala 76:16:@40019.4]
  assign regs_411_io_in = 64'h0; // @[RegFile.scala 75:16:@40018.4]
  assign regs_411_io_reset = reset; // @[RegFile.scala 78:19:@40022.4]
  assign regs_411_io_enable = 1'h1; // @[RegFile.scala 74:20:@40016.4]
  assign regs_412_clock = clock; // @[:@40025.4]
  assign regs_412_reset = io_reset; // @[:@40026.4 RegFile.scala 76:16:@40033.4]
  assign regs_412_io_in = 64'h0; // @[RegFile.scala 75:16:@40032.4]
  assign regs_412_io_reset = reset; // @[RegFile.scala 78:19:@40036.4]
  assign regs_412_io_enable = 1'h1; // @[RegFile.scala 74:20:@40030.4]
  assign regs_413_clock = clock; // @[:@40039.4]
  assign regs_413_reset = io_reset; // @[:@40040.4 RegFile.scala 76:16:@40047.4]
  assign regs_413_io_in = 64'h0; // @[RegFile.scala 75:16:@40046.4]
  assign regs_413_io_reset = reset; // @[RegFile.scala 78:19:@40050.4]
  assign regs_413_io_enable = 1'h1; // @[RegFile.scala 74:20:@40044.4]
  assign regs_414_clock = clock; // @[:@40053.4]
  assign regs_414_reset = io_reset; // @[:@40054.4 RegFile.scala 76:16:@40061.4]
  assign regs_414_io_in = 64'h0; // @[RegFile.scala 75:16:@40060.4]
  assign regs_414_io_reset = reset; // @[RegFile.scala 78:19:@40064.4]
  assign regs_414_io_enable = 1'h1; // @[RegFile.scala 74:20:@40058.4]
  assign regs_415_clock = clock; // @[:@40067.4]
  assign regs_415_reset = io_reset; // @[:@40068.4 RegFile.scala 76:16:@40075.4]
  assign regs_415_io_in = 64'h0; // @[RegFile.scala 75:16:@40074.4]
  assign regs_415_io_reset = reset; // @[RegFile.scala 78:19:@40078.4]
  assign regs_415_io_enable = 1'h1; // @[RegFile.scala 74:20:@40072.4]
  assign regs_416_clock = clock; // @[:@40081.4]
  assign regs_416_reset = io_reset; // @[:@40082.4 RegFile.scala 76:16:@40089.4]
  assign regs_416_io_in = 64'h0; // @[RegFile.scala 75:16:@40088.4]
  assign regs_416_io_reset = reset; // @[RegFile.scala 78:19:@40092.4]
  assign regs_416_io_enable = 1'h1; // @[RegFile.scala 74:20:@40086.4]
  assign regs_417_clock = clock; // @[:@40095.4]
  assign regs_417_reset = io_reset; // @[:@40096.4 RegFile.scala 76:16:@40103.4]
  assign regs_417_io_in = 64'h0; // @[RegFile.scala 75:16:@40102.4]
  assign regs_417_io_reset = reset; // @[RegFile.scala 78:19:@40106.4]
  assign regs_417_io_enable = 1'h1; // @[RegFile.scala 74:20:@40100.4]
  assign regs_418_clock = clock; // @[:@40109.4]
  assign regs_418_reset = io_reset; // @[:@40110.4 RegFile.scala 76:16:@40117.4]
  assign regs_418_io_in = 64'h0; // @[RegFile.scala 75:16:@40116.4]
  assign regs_418_io_reset = reset; // @[RegFile.scala 78:19:@40120.4]
  assign regs_418_io_enable = 1'h1; // @[RegFile.scala 74:20:@40114.4]
  assign regs_419_clock = clock; // @[:@40123.4]
  assign regs_419_reset = io_reset; // @[:@40124.4 RegFile.scala 76:16:@40131.4]
  assign regs_419_io_in = 64'h0; // @[RegFile.scala 75:16:@40130.4]
  assign regs_419_io_reset = reset; // @[RegFile.scala 78:19:@40134.4]
  assign regs_419_io_enable = 1'h1; // @[RegFile.scala 74:20:@40128.4]
  assign regs_420_clock = clock; // @[:@40137.4]
  assign regs_420_reset = io_reset; // @[:@40138.4 RegFile.scala 76:16:@40145.4]
  assign regs_420_io_in = 64'h0; // @[RegFile.scala 75:16:@40144.4]
  assign regs_420_io_reset = reset; // @[RegFile.scala 78:19:@40148.4]
  assign regs_420_io_enable = 1'h1; // @[RegFile.scala 74:20:@40142.4]
  assign regs_421_clock = clock; // @[:@40151.4]
  assign regs_421_reset = io_reset; // @[:@40152.4 RegFile.scala 76:16:@40159.4]
  assign regs_421_io_in = 64'h0; // @[RegFile.scala 75:16:@40158.4]
  assign regs_421_io_reset = reset; // @[RegFile.scala 78:19:@40162.4]
  assign regs_421_io_enable = 1'h1; // @[RegFile.scala 74:20:@40156.4]
  assign regs_422_clock = clock; // @[:@40165.4]
  assign regs_422_reset = io_reset; // @[:@40166.4 RegFile.scala 76:16:@40173.4]
  assign regs_422_io_in = 64'h0; // @[RegFile.scala 75:16:@40172.4]
  assign regs_422_io_reset = reset; // @[RegFile.scala 78:19:@40176.4]
  assign regs_422_io_enable = 1'h1; // @[RegFile.scala 74:20:@40170.4]
  assign regs_423_clock = clock; // @[:@40179.4]
  assign regs_423_reset = io_reset; // @[:@40180.4 RegFile.scala 76:16:@40187.4]
  assign regs_423_io_in = 64'h0; // @[RegFile.scala 75:16:@40186.4]
  assign regs_423_io_reset = reset; // @[RegFile.scala 78:19:@40190.4]
  assign regs_423_io_enable = 1'h1; // @[RegFile.scala 74:20:@40184.4]
  assign regs_424_clock = clock; // @[:@40193.4]
  assign regs_424_reset = io_reset; // @[:@40194.4 RegFile.scala 76:16:@40201.4]
  assign regs_424_io_in = 64'h0; // @[RegFile.scala 75:16:@40200.4]
  assign regs_424_io_reset = reset; // @[RegFile.scala 78:19:@40204.4]
  assign regs_424_io_enable = 1'h1; // @[RegFile.scala 74:20:@40198.4]
  assign regs_425_clock = clock; // @[:@40207.4]
  assign regs_425_reset = io_reset; // @[:@40208.4 RegFile.scala 76:16:@40215.4]
  assign regs_425_io_in = 64'h0; // @[RegFile.scala 75:16:@40214.4]
  assign regs_425_io_reset = reset; // @[RegFile.scala 78:19:@40218.4]
  assign regs_425_io_enable = 1'h1; // @[RegFile.scala 74:20:@40212.4]
  assign regs_426_clock = clock; // @[:@40221.4]
  assign regs_426_reset = io_reset; // @[:@40222.4 RegFile.scala 76:16:@40229.4]
  assign regs_426_io_in = 64'h0; // @[RegFile.scala 75:16:@40228.4]
  assign regs_426_io_reset = reset; // @[RegFile.scala 78:19:@40232.4]
  assign regs_426_io_enable = 1'h1; // @[RegFile.scala 74:20:@40226.4]
  assign regs_427_clock = clock; // @[:@40235.4]
  assign regs_427_reset = io_reset; // @[:@40236.4 RegFile.scala 76:16:@40243.4]
  assign regs_427_io_in = 64'h0; // @[RegFile.scala 75:16:@40242.4]
  assign regs_427_io_reset = reset; // @[RegFile.scala 78:19:@40246.4]
  assign regs_427_io_enable = 1'h1; // @[RegFile.scala 74:20:@40240.4]
  assign regs_428_clock = clock; // @[:@40249.4]
  assign regs_428_reset = io_reset; // @[:@40250.4 RegFile.scala 76:16:@40257.4]
  assign regs_428_io_in = 64'h0; // @[RegFile.scala 75:16:@40256.4]
  assign regs_428_io_reset = reset; // @[RegFile.scala 78:19:@40260.4]
  assign regs_428_io_enable = 1'h1; // @[RegFile.scala 74:20:@40254.4]
  assign regs_429_clock = clock; // @[:@40263.4]
  assign regs_429_reset = io_reset; // @[:@40264.4 RegFile.scala 76:16:@40271.4]
  assign regs_429_io_in = 64'h0; // @[RegFile.scala 75:16:@40270.4]
  assign regs_429_io_reset = reset; // @[RegFile.scala 78:19:@40274.4]
  assign regs_429_io_enable = 1'h1; // @[RegFile.scala 74:20:@40268.4]
  assign regs_430_clock = clock; // @[:@40277.4]
  assign regs_430_reset = io_reset; // @[:@40278.4 RegFile.scala 76:16:@40285.4]
  assign regs_430_io_in = 64'h0; // @[RegFile.scala 75:16:@40284.4]
  assign regs_430_io_reset = reset; // @[RegFile.scala 78:19:@40288.4]
  assign regs_430_io_enable = 1'h1; // @[RegFile.scala 74:20:@40282.4]
  assign regs_431_clock = clock; // @[:@40291.4]
  assign regs_431_reset = io_reset; // @[:@40292.4 RegFile.scala 76:16:@40299.4]
  assign regs_431_io_in = 64'h0; // @[RegFile.scala 75:16:@40298.4]
  assign regs_431_io_reset = reset; // @[RegFile.scala 78:19:@40302.4]
  assign regs_431_io_enable = 1'h1; // @[RegFile.scala 74:20:@40296.4]
  assign regs_432_clock = clock; // @[:@40305.4]
  assign regs_432_reset = io_reset; // @[:@40306.4 RegFile.scala 76:16:@40313.4]
  assign regs_432_io_in = 64'h0; // @[RegFile.scala 75:16:@40312.4]
  assign regs_432_io_reset = reset; // @[RegFile.scala 78:19:@40316.4]
  assign regs_432_io_enable = 1'h1; // @[RegFile.scala 74:20:@40310.4]
  assign regs_433_clock = clock; // @[:@40319.4]
  assign regs_433_reset = io_reset; // @[:@40320.4 RegFile.scala 76:16:@40327.4]
  assign regs_433_io_in = 64'h0; // @[RegFile.scala 75:16:@40326.4]
  assign regs_433_io_reset = reset; // @[RegFile.scala 78:19:@40330.4]
  assign regs_433_io_enable = 1'h1; // @[RegFile.scala 74:20:@40324.4]
  assign regs_434_clock = clock; // @[:@40333.4]
  assign regs_434_reset = io_reset; // @[:@40334.4 RegFile.scala 76:16:@40341.4]
  assign regs_434_io_in = 64'h0; // @[RegFile.scala 75:16:@40340.4]
  assign regs_434_io_reset = reset; // @[RegFile.scala 78:19:@40344.4]
  assign regs_434_io_enable = 1'h1; // @[RegFile.scala 74:20:@40338.4]
  assign regs_435_clock = clock; // @[:@40347.4]
  assign regs_435_reset = io_reset; // @[:@40348.4 RegFile.scala 76:16:@40355.4]
  assign regs_435_io_in = 64'h0; // @[RegFile.scala 75:16:@40354.4]
  assign regs_435_io_reset = reset; // @[RegFile.scala 78:19:@40358.4]
  assign regs_435_io_enable = 1'h1; // @[RegFile.scala 74:20:@40352.4]
  assign regs_436_clock = clock; // @[:@40361.4]
  assign regs_436_reset = io_reset; // @[:@40362.4 RegFile.scala 76:16:@40369.4]
  assign regs_436_io_in = 64'h0; // @[RegFile.scala 75:16:@40368.4]
  assign regs_436_io_reset = reset; // @[RegFile.scala 78:19:@40372.4]
  assign regs_436_io_enable = 1'h1; // @[RegFile.scala 74:20:@40366.4]
  assign regs_437_clock = clock; // @[:@40375.4]
  assign regs_437_reset = io_reset; // @[:@40376.4 RegFile.scala 76:16:@40383.4]
  assign regs_437_io_in = 64'h0; // @[RegFile.scala 75:16:@40382.4]
  assign regs_437_io_reset = reset; // @[RegFile.scala 78:19:@40386.4]
  assign regs_437_io_enable = 1'h1; // @[RegFile.scala 74:20:@40380.4]
  assign regs_438_clock = clock; // @[:@40389.4]
  assign regs_438_reset = io_reset; // @[:@40390.4 RegFile.scala 76:16:@40397.4]
  assign regs_438_io_in = 64'h0; // @[RegFile.scala 75:16:@40396.4]
  assign regs_438_io_reset = reset; // @[RegFile.scala 78:19:@40400.4]
  assign regs_438_io_enable = 1'h1; // @[RegFile.scala 74:20:@40394.4]
  assign regs_439_clock = clock; // @[:@40403.4]
  assign regs_439_reset = io_reset; // @[:@40404.4 RegFile.scala 76:16:@40411.4]
  assign regs_439_io_in = 64'h0; // @[RegFile.scala 75:16:@40410.4]
  assign regs_439_io_reset = reset; // @[RegFile.scala 78:19:@40414.4]
  assign regs_439_io_enable = 1'h1; // @[RegFile.scala 74:20:@40408.4]
  assign regs_440_clock = clock; // @[:@40417.4]
  assign regs_440_reset = io_reset; // @[:@40418.4 RegFile.scala 76:16:@40425.4]
  assign regs_440_io_in = 64'h0; // @[RegFile.scala 75:16:@40424.4]
  assign regs_440_io_reset = reset; // @[RegFile.scala 78:19:@40428.4]
  assign regs_440_io_enable = 1'h1; // @[RegFile.scala 74:20:@40422.4]
  assign regs_441_clock = clock; // @[:@40431.4]
  assign regs_441_reset = io_reset; // @[:@40432.4 RegFile.scala 76:16:@40439.4]
  assign regs_441_io_in = 64'h0; // @[RegFile.scala 75:16:@40438.4]
  assign regs_441_io_reset = reset; // @[RegFile.scala 78:19:@40442.4]
  assign regs_441_io_enable = 1'h1; // @[RegFile.scala 74:20:@40436.4]
  assign regs_442_clock = clock; // @[:@40445.4]
  assign regs_442_reset = io_reset; // @[:@40446.4 RegFile.scala 76:16:@40453.4]
  assign regs_442_io_in = 64'h0; // @[RegFile.scala 75:16:@40452.4]
  assign regs_442_io_reset = reset; // @[RegFile.scala 78:19:@40456.4]
  assign regs_442_io_enable = 1'h1; // @[RegFile.scala 74:20:@40450.4]
  assign regs_443_clock = clock; // @[:@40459.4]
  assign regs_443_reset = io_reset; // @[:@40460.4 RegFile.scala 76:16:@40467.4]
  assign regs_443_io_in = 64'h0; // @[RegFile.scala 75:16:@40466.4]
  assign regs_443_io_reset = reset; // @[RegFile.scala 78:19:@40470.4]
  assign regs_443_io_enable = 1'h1; // @[RegFile.scala 74:20:@40464.4]
  assign regs_444_clock = clock; // @[:@40473.4]
  assign regs_444_reset = io_reset; // @[:@40474.4 RegFile.scala 76:16:@40481.4]
  assign regs_444_io_in = 64'h0; // @[RegFile.scala 75:16:@40480.4]
  assign regs_444_io_reset = reset; // @[RegFile.scala 78:19:@40484.4]
  assign regs_444_io_enable = 1'h1; // @[RegFile.scala 74:20:@40478.4]
  assign regs_445_clock = clock; // @[:@40487.4]
  assign regs_445_reset = io_reset; // @[:@40488.4 RegFile.scala 76:16:@40495.4]
  assign regs_445_io_in = 64'h0; // @[RegFile.scala 75:16:@40494.4]
  assign regs_445_io_reset = reset; // @[RegFile.scala 78:19:@40498.4]
  assign regs_445_io_enable = 1'h1; // @[RegFile.scala 74:20:@40492.4]
  assign regs_446_clock = clock; // @[:@40501.4]
  assign regs_446_reset = io_reset; // @[:@40502.4 RegFile.scala 76:16:@40509.4]
  assign regs_446_io_in = 64'h0; // @[RegFile.scala 75:16:@40508.4]
  assign regs_446_io_reset = reset; // @[RegFile.scala 78:19:@40512.4]
  assign regs_446_io_enable = 1'h1; // @[RegFile.scala 74:20:@40506.4]
  assign regs_447_clock = clock; // @[:@40515.4]
  assign regs_447_reset = io_reset; // @[:@40516.4 RegFile.scala 76:16:@40523.4]
  assign regs_447_io_in = 64'h0; // @[RegFile.scala 75:16:@40522.4]
  assign regs_447_io_reset = reset; // @[RegFile.scala 78:19:@40526.4]
  assign regs_447_io_enable = 1'h1; // @[RegFile.scala 74:20:@40520.4]
  assign regs_448_clock = clock; // @[:@40529.4]
  assign regs_448_reset = io_reset; // @[:@40530.4 RegFile.scala 76:16:@40537.4]
  assign regs_448_io_in = 64'h0; // @[RegFile.scala 75:16:@40536.4]
  assign regs_448_io_reset = reset; // @[RegFile.scala 78:19:@40540.4]
  assign regs_448_io_enable = 1'h1; // @[RegFile.scala 74:20:@40534.4]
  assign regs_449_clock = clock; // @[:@40543.4]
  assign regs_449_reset = io_reset; // @[:@40544.4 RegFile.scala 76:16:@40551.4]
  assign regs_449_io_in = 64'h0; // @[RegFile.scala 75:16:@40550.4]
  assign regs_449_io_reset = reset; // @[RegFile.scala 78:19:@40554.4]
  assign regs_449_io_enable = 1'h1; // @[RegFile.scala 74:20:@40548.4]
  assign regs_450_clock = clock; // @[:@40557.4]
  assign regs_450_reset = io_reset; // @[:@40558.4 RegFile.scala 76:16:@40565.4]
  assign regs_450_io_in = 64'h0; // @[RegFile.scala 75:16:@40564.4]
  assign regs_450_io_reset = reset; // @[RegFile.scala 78:19:@40568.4]
  assign regs_450_io_enable = 1'h1; // @[RegFile.scala 74:20:@40562.4]
  assign regs_451_clock = clock; // @[:@40571.4]
  assign regs_451_reset = io_reset; // @[:@40572.4 RegFile.scala 76:16:@40579.4]
  assign regs_451_io_in = 64'h0; // @[RegFile.scala 75:16:@40578.4]
  assign regs_451_io_reset = reset; // @[RegFile.scala 78:19:@40582.4]
  assign regs_451_io_enable = 1'h1; // @[RegFile.scala 74:20:@40576.4]
  assign regs_452_clock = clock; // @[:@40585.4]
  assign regs_452_reset = io_reset; // @[:@40586.4 RegFile.scala 76:16:@40593.4]
  assign regs_452_io_in = 64'h0; // @[RegFile.scala 75:16:@40592.4]
  assign regs_452_io_reset = reset; // @[RegFile.scala 78:19:@40596.4]
  assign regs_452_io_enable = 1'h1; // @[RegFile.scala 74:20:@40590.4]
  assign regs_453_clock = clock; // @[:@40599.4]
  assign regs_453_reset = io_reset; // @[:@40600.4 RegFile.scala 76:16:@40607.4]
  assign regs_453_io_in = 64'h0; // @[RegFile.scala 75:16:@40606.4]
  assign regs_453_io_reset = reset; // @[RegFile.scala 78:19:@40610.4]
  assign regs_453_io_enable = 1'h1; // @[RegFile.scala 74:20:@40604.4]
  assign regs_454_clock = clock; // @[:@40613.4]
  assign regs_454_reset = io_reset; // @[:@40614.4 RegFile.scala 76:16:@40621.4]
  assign regs_454_io_in = 64'h0; // @[RegFile.scala 75:16:@40620.4]
  assign regs_454_io_reset = reset; // @[RegFile.scala 78:19:@40624.4]
  assign regs_454_io_enable = 1'h1; // @[RegFile.scala 74:20:@40618.4]
  assign regs_455_clock = clock; // @[:@40627.4]
  assign regs_455_reset = io_reset; // @[:@40628.4 RegFile.scala 76:16:@40635.4]
  assign regs_455_io_in = 64'h0; // @[RegFile.scala 75:16:@40634.4]
  assign regs_455_io_reset = reset; // @[RegFile.scala 78:19:@40638.4]
  assign regs_455_io_enable = 1'h1; // @[RegFile.scala 74:20:@40632.4]
  assign regs_456_clock = clock; // @[:@40641.4]
  assign regs_456_reset = io_reset; // @[:@40642.4 RegFile.scala 76:16:@40649.4]
  assign regs_456_io_in = 64'h0; // @[RegFile.scala 75:16:@40648.4]
  assign regs_456_io_reset = reset; // @[RegFile.scala 78:19:@40652.4]
  assign regs_456_io_enable = 1'h1; // @[RegFile.scala 74:20:@40646.4]
  assign regs_457_clock = clock; // @[:@40655.4]
  assign regs_457_reset = io_reset; // @[:@40656.4 RegFile.scala 76:16:@40663.4]
  assign regs_457_io_in = 64'h0; // @[RegFile.scala 75:16:@40662.4]
  assign regs_457_io_reset = reset; // @[RegFile.scala 78:19:@40666.4]
  assign regs_457_io_enable = 1'h1; // @[RegFile.scala 74:20:@40660.4]
  assign regs_458_clock = clock; // @[:@40669.4]
  assign regs_458_reset = io_reset; // @[:@40670.4 RegFile.scala 76:16:@40677.4]
  assign regs_458_io_in = 64'h0; // @[RegFile.scala 75:16:@40676.4]
  assign regs_458_io_reset = reset; // @[RegFile.scala 78:19:@40680.4]
  assign regs_458_io_enable = 1'h1; // @[RegFile.scala 74:20:@40674.4]
  assign regs_459_clock = clock; // @[:@40683.4]
  assign regs_459_reset = io_reset; // @[:@40684.4 RegFile.scala 76:16:@40691.4]
  assign regs_459_io_in = 64'h0; // @[RegFile.scala 75:16:@40690.4]
  assign regs_459_io_reset = reset; // @[RegFile.scala 78:19:@40694.4]
  assign regs_459_io_enable = 1'h1; // @[RegFile.scala 74:20:@40688.4]
  assign regs_460_clock = clock; // @[:@40697.4]
  assign regs_460_reset = io_reset; // @[:@40698.4 RegFile.scala 76:16:@40705.4]
  assign regs_460_io_in = 64'h0; // @[RegFile.scala 75:16:@40704.4]
  assign regs_460_io_reset = reset; // @[RegFile.scala 78:19:@40708.4]
  assign regs_460_io_enable = 1'h1; // @[RegFile.scala 74:20:@40702.4]
  assign regs_461_clock = clock; // @[:@40711.4]
  assign regs_461_reset = io_reset; // @[:@40712.4 RegFile.scala 76:16:@40719.4]
  assign regs_461_io_in = 64'h0; // @[RegFile.scala 75:16:@40718.4]
  assign regs_461_io_reset = reset; // @[RegFile.scala 78:19:@40722.4]
  assign regs_461_io_enable = 1'h1; // @[RegFile.scala 74:20:@40716.4]
  assign regs_462_clock = clock; // @[:@40725.4]
  assign regs_462_reset = io_reset; // @[:@40726.4 RegFile.scala 76:16:@40733.4]
  assign regs_462_io_in = 64'h0; // @[RegFile.scala 75:16:@40732.4]
  assign regs_462_io_reset = reset; // @[RegFile.scala 78:19:@40736.4]
  assign regs_462_io_enable = 1'h1; // @[RegFile.scala 74:20:@40730.4]
  assign regs_463_clock = clock; // @[:@40739.4]
  assign regs_463_reset = io_reset; // @[:@40740.4 RegFile.scala 76:16:@40747.4]
  assign regs_463_io_in = 64'h0; // @[RegFile.scala 75:16:@40746.4]
  assign regs_463_io_reset = reset; // @[RegFile.scala 78:19:@40750.4]
  assign regs_463_io_enable = 1'h1; // @[RegFile.scala 74:20:@40744.4]
  assign regs_464_clock = clock; // @[:@40753.4]
  assign regs_464_reset = io_reset; // @[:@40754.4 RegFile.scala 76:16:@40761.4]
  assign regs_464_io_in = 64'h0; // @[RegFile.scala 75:16:@40760.4]
  assign regs_464_io_reset = reset; // @[RegFile.scala 78:19:@40764.4]
  assign regs_464_io_enable = 1'h1; // @[RegFile.scala 74:20:@40758.4]
  assign regs_465_clock = clock; // @[:@40767.4]
  assign regs_465_reset = io_reset; // @[:@40768.4 RegFile.scala 76:16:@40775.4]
  assign regs_465_io_in = 64'h0; // @[RegFile.scala 75:16:@40774.4]
  assign regs_465_io_reset = reset; // @[RegFile.scala 78:19:@40778.4]
  assign regs_465_io_enable = 1'h1; // @[RegFile.scala 74:20:@40772.4]
  assign regs_466_clock = clock; // @[:@40781.4]
  assign regs_466_reset = io_reset; // @[:@40782.4 RegFile.scala 76:16:@40789.4]
  assign regs_466_io_in = 64'h0; // @[RegFile.scala 75:16:@40788.4]
  assign regs_466_io_reset = reset; // @[RegFile.scala 78:19:@40792.4]
  assign regs_466_io_enable = 1'h1; // @[RegFile.scala 74:20:@40786.4]
  assign regs_467_clock = clock; // @[:@40795.4]
  assign regs_467_reset = io_reset; // @[:@40796.4 RegFile.scala 76:16:@40803.4]
  assign regs_467_io_in = 64'h0; // @[RegFile.scala 75:16:@40802.4]
  assign regs_467_io_reset = reset; // @[RegFile.scala 78:19:@40806.4]
  assign regs_467_io_enable = 1'h1; // @[RegFile.scala 74:20:@40800.4]
  assign regs_468_clock = clock; // @[:@40809.4]
  assign regs_468_reset = io_reset; // @[:@40810.4 RegFile.scala 76:16:@40817.4]
  assign regs_468_io_in = 64'h0; // @[RegFile.scala 75:16:@40816.4]
  assign regs_468_io_reset = reset; // @[RegFile.scala 78:19:@40820.4]
  assign regs_468_io_enable = 1'h1; // @[RegFile.scala 74:20:@40814.4]
  assign regs_469_clock = clock; // @[:@40823.4]
  assign regs_469_reset = io_reset; // @[:@40824.4 RegFile.scala 76:16:@40831.4]
  assign regs_469_io_in = 64'h0; // @[RegFile.scala 75:16:@40830.4]
  assign regs_469_io_reset = reset; // @[RegFile.scala 78:19:@40834.4]
  assign regs_469_io_enable = 1'h1; // @[RegFile.scala 74:20:@40828.4]
  assign regs_470_clock = clock; // @[:@40837.4]
  assign regs_470_reset = io_reset; // @[:@40838.4 RegFile.scala 76:16:@40845.4]
  assign regs_470_io_in = 64'h0; // @[RegFile.scala 75:16:@40844.4]
  assign regs_470_io_reset = reset; // @[RegFile.scala 78:19:@40848.4]
  assign regs_470_io_enable = 1'h1; // @[RegFile.scala 74:20:@40842.4]
  assign regs_471_clock = clock; // @[:@40851.4]
  assign regs_471_reset = io_reset; // @[:@40852.4 RegFile.scala 76:16:@40859.4]
  assign regs_471_io_in = 64'h0; // @[RegFile.scala 75:16:@40858.4]
  assign regs_471_io_reset = reset; // @[RegFile.scala 78:19:@40862.4]
  assign regs_471_io_enable = 1'h1; // @[RegFile.scala 74:20:@40856.4]
  assign regs_472_clock = clock; // @[:@40865.4]
  assign regs_472_reset = io_reset; // @[:@40866.4 RegFile.scala 76:16:@40873.4]
  assign regs_472_io_in = 64'h0; // @[RegFile.scala 75:16:@40872.4]
  assign regs_472_io_reset = reset; // @[RegFile.scala 78:19:@40876.4]
  assign regs_472_io_enable = 1'h1; // @[RegFile.scala 74:20:@40870.4]
  assign regs_473_clock = clock; // @[:@40879.4]
  assign regs_473_reset = io_reset; // @[:@40880.4 RegFile.scala 76:16:@40887.4]
  assign regs_473_io_in = 64'h0; // @[RegFile.scala 75:16:@40886.4]
  assign regs_473_io_reset = reset; // @[RegFile.scala 78:19:@40890.4]
  assign regs_473_io_enable = 1'h1; // @[RegFile.scala 74:20:@40884.4]
  assign regs_474_clock = clock; // @[:@40893.4]
  assign regs_474_reset = io_reset; // @[:@40894.4 RegFile.scala 76:16:@40901.4]
  assign regs_474_io_in = 64'h0; // @[RegFile.scala 75:16:@40900.4]
  assign regs_474_io_reset = reset; // @[RegFile.scala 78:19:@40904.4]
  assign regs_474_io_enable = 1'h1; // @[RegFile.scala 74:20:@40898.4]
  assign regs_475_clock = clock; // @[:@40907.4]
  assign regs_475_reset = io_reset; // @[:@40908.4 RegFile.scala 76:16:@40915.4]
  assign regs_475_io_in = 64'h0; // @[RegFile.scala 75:16:@40914.4]
  assign regs_475_io_reset = reset; // @[RegFile.scala 78:19:@40918.4]
  assign regs_475_io_enable = 1'h1; // @[RegFile.scala 74:20:@40912.4]
  assign regs_476_clock = clock; // @[:@40921.4]
  assign regs_476_reset = io_reset; // @[:@40922.4 RegFile.scala 76:16:@40929.4]
  assign regs_476_io_in = 64'h0; // @[RegFile.scala 75:16:@40928.4]
  assign regs_476_io_reset = reset; // @[RegFile.scala 78:19:@40932.4]
  assign regs_476_io_enable = 1'h1; // @[RegFile.scala 74:20:@40926.4]
  assign regs_477_clock = clock; // @[:@40935.4]
  assign regs_477_reset = io_reset; // @[:@40936.4 RegFile.scala 76:16:@40943.4]
  assign regs_477_io_in = 64'h0; // @[RegFile.scala 75:16:@40942.4]
  assign regs_477_io_reset = reset; // @[RegFile.scala 78:19:@40946.4]
  assign regs_477_io_enable = 1'h1; // @[RegFile.scala 74:20:@40940.4]
  assign regs_478_clock = clock; // @[:@40949.4]
  assign regs_478_reset = io_reset; // @[:@40950.4 RegFile.scala 76:16:@40957.4]
  assign regs_478_io_in = 64'h0; // @[RegFile.scala 75:16:@40956.4]
  assign regs_478_io_reset = reset; // @[RegFile.scala 78:19:@40960.4]
  assign regs_478_io_enable = 1'h1; // @[RegFile.scala 74:20:@40954.4]
  assign regs_479_clock = clock; // @[:@40963.4]
  assign regs_479_reset = io_reset; // @[:@40964.4 RegFile.scala 76:16:@40971.4]
  assign regs_479_io_in = 64'h0; // @[RegFile.scala 75:16:@40970.4]
  assign regs_479_io_reset = reset; // @[RegFile.scala 78:19:@40974.4]
  assign regs_479_io_enable = 1'h1; // @[RegFile.scala 74:20:@40968.4]
  assign regs_480_clock = clock; // @[:@40977.4]
  assign regs_480_reset = io_reset; // @[:@40978.4 RegFile.scala 76:16:@40985.4]
  assign regs_480_io_in = 64'h0; // @[RegFile.scala 75:16:@40984.4]
  assign regs_480_io_reset = reset; // @[RegFile.scala 78:19:@40988.4]
  assign regs_480_io_enable = 1'h1; // @[RegFile.scala 74:20:@40982.4]
  assign regs_481_clock = clock; // @[:@40991.4]
  assign regs_481_reset = io_reset; // @[:@40992.4 RegFile.scala 76:16:@40999.4]
  assign regs_481_io_in = 64'h0; // @[RegFile.scala 75:16:@40998.4]
  assign regs_481_io_reset = reset; // @[RegFile.scala 78:19:@41002.4]
  assign regs_481_io_enable = 1'h1; // @[RegFile.scala 74:20:@40996.4]
  assign regs_482_clock = clock; // @[:@41005.4]
  assign regs_482_reset = io_reset; // @[:@41006.4 RegFile.scala 76:16:@41013.4]
  assign regs_482_io_in = 64'h0; // @[RegFile.scala 75:16:@41012.4]
  assign regs_482_io_reset = reset; // @[RegFile.scala 78:19:@41016.4]
  assign regs_482_io_enable = 1'h1; // @[RegFile.scala 74:20:@41010.4]
  assign regs_483_clock = clock; // @[:@41019.4]
  assign regs_483_reset = io_reset; // @[:@41020.4 RegFile.scala 76:16:@41027.4]
  assign regs_483_io_in = 64'h0; // @[RegFile.scala 75:16:@41026.4]
  assign regs_483_io_reset = reset; // @[RegFile.scala 78:19:@41030.4]
  assign regs_483_io_enable = 1'h1; // @[RegFile.scala 74:20:@41024.4]
  assign regs_484_clock = clock; // @[:@41033.4]
  assign regs_484_reset = io_reset; // @[:@41034.4 RegFile.scala 76:16:@41041.4]
  assign regs_484_io_in = 64'h0; // @[RegFile.scala 75:16:@41040.4]
  assign regs_484_io_reset = reset; // @[RegFile.scala 78:19:@41044.4]
  assign regs_484_io_enable = 1'h1; // @[RegFile.scala 74:20:@41038.4]
  assign regs_485_clock = clock; // @[:@41047.4]
  assign regs_485_reset = io_reset; // @[:@41048.4 RegFile.scala 76:16:@41055.4]
  assign regs_485_io_in = 64'h0; // @[RegFile.scala 75:16:@41054.4]
  assign regs_485_io_reset = reset; // @[RegFile.scala 78:19:@41058.4]
  assign regs_485_io_enable = 1'h1; // @[RegFile.scala 74:20:@41052.4]
  assign regs_486_clock = clock; // @[:@41061.4]
  assign regs_486_reset = io_reset; // @[:@41062.4 RegFile.scala 76:16:@41069.4]
  assign regs_486_io_in = 64'h0; // @[RegFile.scala 75:16:@41068.4]
  assign regs_486_io_reset = reset; // @[RegFile.scala 78:19:@41072.4]
  assign regs_486_io_enable = 1'h1; // @[RegFile.scala 74:20:@41066.4]
  assign regs_487_clock = clock; // @[:@41075.4]
  assign regs_487_reset = io_reset; // @[:@41076.4 RegFile.scala 76:16:@41083.4]
  assign regs_487_io_in = 64'h0; // @[RegFile.scala 75:16:@41082.4]
  assign regs_487_io_reset = reset; // @[RegFile.scala 78:19:@41086.4]
  assign regs_487_io_enable = 1'h1; // @[RegFile.scala 74:20:@41080.4]
  assign regs_488_clock = clock; // @[:@41089.4]
  assign regs_488_reset = io_reset; // @[:@41090.4 RegFile.scala 76:16:@41097.4]
  assign regs_488_io_in = 64'h0; // @[RegFile.scala 75:16:@41096.4]
  assign regs_488_io_reset = reset; // @[RegFile.scala 78:19:@41100.4]
  assign regs_488_io_enable = 1'h1; // @[RegFile.scala 74:20:@41094.4]
  assign regs_489_clock = clock; // @[:@41103.4]
  assign regs_489_reset = io_reset; // @[:@41104.4 RegFile.scala 76:16:@41111.4]
  assign regs_489_io_in = 64'h0; // @[RegFile.scala 75:16:@41110.4]
  assign regs_489_io_reset = reset; // @[RegFile.scala 78:19:@41114.4]
  assign regs_489_io_enable = 1'h1; // @[RegFile.scala 74:20:@41108.4]
  assign regs_490_clock = clock; // @[:@41117.4]
  assign regs_490_reset = io_reset; // @[:@41118.4 RegFile.scala 76:16:@41125.4]
  assign regs_490_io_in = 64'h0; // @[RegFile.scala 75:16:@41124.4]
  assign regs_490_io_reset = reset; // @[RegFile.scala 78:19:@41128.4]
  assign regs_490_io_enable = 1'h1; // @[RegFile.scala 74:20:@41122.4]
  assign regs_491_clock = clock; // @[:@41131.4]
  assign regs_491_reset = io_reset; // @[:@41132.4 RegFile.scala 76:16:@41139.4]
  assign regs_491_io_in = 64'h0; // @[RegFile.scala 75:16:@41138.4]
  assign regs_491_io_reset = reset; // @[RegFile.scala 78:19:@41142.4]
  assign regs_491_io_enable = 1'h1; // @[RegFile.scala 74:20:@41136.4]
  assign regs_492_clock = clock; // @[:@41145.4]
  assign regs_492_reset = io_reset; // @[:@41146.4 RegFile.scala 76:16:@41153.4]
  assign regs_492_io_in = 64'h0; // @[RegFile.scala 75:16:@41152.4]
  assign regs_492_io_reset = reset; // @[RegFile.scala 78:19:@41156.4]
  assign regs_492_io_enable = 1'h1; // @[RegFile.scala 74:20:@41150.4]
  assign regs_493_clock = clock; // @[:@41159.4]
  assign regs_493_reset = io_reset; // @[:@41160.4 RegFile.scala 76:16:@41167.4]
  assign regs_493_io_in = 64'h0; // @[RegFile.scala 75:16:@41166.4]
  assign regs_493_io_reset = reset; // @[RegFile.scala 78:19:@41170.4]
  assign regs_493_io_enable = 1'h1; // @[RegFile.scala 74:20:@41164.4]
  assign regs_494_clock = clock; // @[:@41173.4]
  assign regs_494_reset = io_reset; // @[:@41174.4 RegFile.scala 76:16:@41181.4]
  assign regs_494_io_in = 64'h0; // @[RegFile.scala 75:16:@41180.4]
  assign regs_494_io_reset = reset; // @[RegFile.scala 78:19:@41184.4]
  assign regs_494_io_enable = 1'h1; // @[RegFile.scala 74:20:@41178.4]
  assign regs_495_clock = clock; // @[:@41187.4]
  assign regs_495_reset = io_reset; // @[:@41188.4 RegFile.scala 76:16:@41195.4]
  assign regs_495_io_in = 64'h0; // @[RegFile.scala 75:16:@41194.4]
  assign regs_495_io_reset = reset; // @[RegFile.scala 78:19:@41198.4]
  assign regs_495_io_enable = 1'h1; // @[RegFile.scala 74:20:@41192.4]
  assign regs_496_clock = clock; // @[:@41201.4]
  assign regs_496_reset = io_reset; // @[:@41202.4 RegFile.scala 76:16:@41209.4]
  assign regs_496_io_in = 64'h0; // @[RegFile.scala 75:16:@41208.4]
  assign regs_496_io_reset = reset; // @[RegFile.scala 78:19:@41212.4]
  assign regs_496_io_enable = 1'h1; // @[RegFile.scala 74:20:@41206.4]
  assign regs_497_clock = clock; // @[:@41215.4]
  assign regs_497_reset = io_reset; // @[:@41216.4 RegFile.scala 76:16:@41223.4]
  assign regs_497_io_in = 64'h0; // @[RegFile.scala 75:16:@41222.4]
  assign regs_497_io_reset = reset; // @[RegFile.scala 78:19:@41226.4]
  assign regs_497_io_enable = 1'h1; // @[RegFile.scala 74:20:@41220.4]
  assign regs_498_clock = clock; // @[:@41229.4]
  assign regs_498_reset = io_reset; // @[:@41230.4 RegFile.scala 76:16:@41237.4]
  assign regs_498_io_in = 64'h0; // @[RegFile.scala 75:16:@41236.4]
  assign regs_498_io_reset = reset; // @[RegFile.scala 78:19:@41240.4]
  assign regs_498_io_enable = 1'h1; // @[RegFile.scala 74:20:@41234.4]
  assign regs_499_clock = clock; // @[:@41243.4]
  assign regs_499_reset = io_reset; // @[:@41244.4 RegFile.scala 76:16:@41251.4]
  assign regs_499_io_in = 64'h0; // @[RegFile.scala 75:16:@41250.4]
  assign regs_499_io_reset = reset; // @[RegFile.scala 78:19:@41254.4]
  assign regs_499_io_enable = 1'h1; // @[RegFile.scala 74:20:@41248.4]
  assign regs_500_clock = clock; // @[:@41257.4]
  assign regs_500_reset = io_reset; // @[:@41258.4 RegFile.scala 76:16:@41265.4]
  assign regs_500_io_in = 64'h0; // @[RegFile.scala 75:16:@41264.4]
  assign regs_500_io_reset = reset; // @[RegFile.scala 78:19:@41268.4]
  assign regs_500_io_enable = 1'h1; // @[RegFile.scala 74:20:@41262.4]
  assign regs_501_clock = clock; // @[:@41271.4]
  assign regs_501_reset = io_reset; // @[:@41272.4 RegFile.scala 76:16:@41279.4]
  assign regs_501_io_in = 64'h0; // @[RegFile.scala 75:16:@41278.4]
  assign regs_501_io_reset = reset; // @[RegFile.scala 78:19:@41282.4]
  assign regs_501_io_enable = 1'h1; // @[RegFile.scala 74:20:@41276.4]
  assign regs_502_clock = clock; // @[:@41285.4]
  assign regs_502_reset = io_reset; // @[:@41286.4 RegFile.scala 76:16:@41293.4]
  assign regs_502_io_in = 64'h0; // @[RegFile.scala 75:16:@41292.4]
  assign regs_502_io_reset = reset; // @[RegFile.scala 78:19:@41296.4]
  assign regs_502_io_enable = 1'h1; // @[RegFile.scala 74:20:@41290.4]
  assign rport_io_ins_0 = regs_0_io_out; // @[RegFile.scala 97:16:@41805.4]
  assign rport_io_ins_1 = regs_1_io_out; // @[RegFile.scala 97:16:@41806.4]
  assign rport_io_ins_2 = regs_2_io_out; // @[RegFile.scala 97:16:@41807.4]
  assign rport_io_ins_3 = regs_3_io_out; // @[RegFile.scala 97:16:@41808.4]
  assign rport_io_ins_4 = regs_4_io_out; // @[RegFile.scala 97:16:@41809.4]
  assign rport_io_ins_5 = regs_5_io_out; // @[RegFile.scala 97:16:@41810.4]
  assign rport_io_ins_6 = regs_6_io_out; // @[RegFile.scala 97:16:@41811.4]
  assign rport_io_ins_7 = regs_7_io_out; // @[RegFile.scala 97:16:@41812.4]
  assign rport_io_ins_8 = regs_8_io_out; // @[RegFile.scala 97:16:@41813.4]
  assign rport_io_ins_9 = regs_9_io_out; // @[RegFile.scala 97:16:@41814.4]
  assign rport_io_ins_10 = regs_10_io_out; // @[RegFile.scala 97:16:@41815.4]
  assign rport_io_ins_11 = regs_11_io_out; // @[RegFile.scala 97:16:@41816.4]
  assign rport_io_ins_12 = regs_12_io_out; // @[RegFile.scala 97:16:@41817.4]
  assign rport_io_ins_13 = regs_13_io_out; // @[RegFile.scala 97:16:@41818.4]
  assign rport_io_ins_14 = regs_14_io_out; // @[RegFile.scala 97:16:@41819.4]
  assign rport_io_ins_15 = regs_15_io_out; // @[RegFile.scala 97:16:@41820.4]
  assign rport_io_ins_16 = regs_16_io_out; // @[RegFile.scala 97:16:@41821.4]
  assign rport_io_ins_17 = regs_17_io_out; // @[RegFile.scala 97:16:@41822.4]
  assign rport_io_ins_18 = regs_18_io_out; // @[RegFile.scala 97:16:@41823.4]
  assign rport_io_ins_19 = regs_19_io_out; // @[RegFile.scala 97:16:@41824.4]
  assign rport_io_ins_20 = regs_20_io_out; // @[RegFile.scala 97:16:@41825.4]
  assign rport_io_ins_21 = regs_21_io_out; // @[RegFile.scala 97:16:@41826.4]
  assign rport_io_ins_22 = regs_22_io_out; // @[RegFile.scala 97:16:@41827.4]
  assign rport_io_ins_23 = regs_23_io_out; // @[RegFile.scala 97:16:@41828.4]
  assign rport_io_ins_24 = regs_24_io_out; // @[RegFile.scala 97:16:@41829.4]
  assign rport_io_ins_25 = regs_25_io_out; // @[RegFile.scala 97:16:@41830.4]
  assign rport_io_ins_26 = regs_26_io_out; // @[RegFile.scala 97:16:@41831.4]
  assign rport_io_ins_27 = regs_27_io_out; // @[RegFile.scala 97:16:@41832.4]
  assign rport_io_ins_28 = regs_28_io_out; // @[RegFile.scala 97:16:@41833.4]
  assign rport_io_ins_29 = regs_29_io_out; // @[RegFile.scala 97:16:@41834.4]
  assign rport_io_ins_30 = regs_30_io_out; // @[RegFile.scala 97:16:@41835.4]
  assign rport_io_ins_31 = regs_31_io_out; // @[RegFile.scala 97:16:@41836.4]
  assign rport_io_ins_32 = regs_32_io_out; // @[RegFile.scala 97:16:@41837.4]
  assign rport_io_ins_33 = regs_33_io_out; // @[RegFile.scala 97:16:@41838.4]
  assign rport_io_ins_34 = regs_34_io_out; // @[RegFile.scala 97:16:@41839.4]
  assign rport_io_ins_35 = regs_35_io_out; // @[RegFile.scala 97:16:@41840.4]
  assign rport_io_ins_36 = regs_36_io_out; // @[RegFile.scala 97:16:@41841.4]
  assign rport_io_ins_37 = regs_37_io_out; // @[RegFile.scala 97:16:@41842.4]
  assign rport_io_ins_38 = regs_38_io_out; // @[RegFile.scala 97:16:@41843.4]
  assign rport_io_ins_39 = regs_39_io_out; // @[RegFile.scala 97:16:@41844.4]
  assign rport_io_ins_40 = regs_40_io_out; // @[RegFile.scala 97:16:@41845.4]
  assign rport_io_ins_41 = regs_41_io_out; // @[RegFile.scala 97:16:@41846.4]
  assign rport_io_ins_42 = regs_42_io_out; // @[RegFile.scala 97:16:@41847.4]
  assign rport_io_ins_43 = regs_43_io_out; // @[RegFile.scala 97:16:@41848.4]
  assign rport_io_ins_44 = regs_44_io_out; // @[RegFile.scala 97:16:@41849.4]
  assign rport_io_ins_45 = regs_45_io_out; // @[RegFile.scala 97:16:@41850.4]
  assign rport_io_ins_46 = regs_46_io_out; // @[RegFile.scala 97:16:@41851.4]
  assign rport_io_ins_47 = regs_47_io_out; // @[RegFile.scala 97:16:@41852.4]
  assign rport_io_ins_48 = regs_48_io_out; // @[RegFile.scala 97:16:@41853.4]
  assign rport_io_ins_49 = regs_49_io_out; // @[RegFile.scala 97:16:@41854.4]
  assign rport_io_ins_50 = regs_50_io_out; // @[RegFile.scala 97:16:@41855.4]
  assign rport_io_ins_51 = regs_51_io_out; // @[RegFile.scala 97:16:@41856.4]
  assign rport_io_ins_52 = regs_52_io_out; // @[RegFile.scala 97:16:@41857.4]
  assign rport_io_ins_53 = regs_53_io_out; // @[RegFile.scala 97:16:@41858.4]
  assign rport_io_ins_54 = regs_54_io_out; // @[RegFile.scala 97:16:@41859.4]
  assign rport_io_ins_55 = regs_55_io_out; // @[RegFile.scala 97:16:@41860.4]
  assign rport_io_ins_56 = regs_56_io_out; // @[RegFile.scala 97:16:@41861.4]
  assign rport_io_ins_57 = regs_57_io_out; // @[RegFile.scala 97:16:@41862.4]
  assign rport_io_ins_58 = regs_58_io_out; // @[RegFile.scala 97:16:@41863.4]
  assign rport_io_ins_59 = regs_59_io_out; // @[RegFile.scala 97:16:@41864.4]
  assign rport_io_ins_60 = regs_60_io_out; // @[RegFile.scala 97:16:@41865.4]
  assign rport_io_ins_61 = regs_61_io_out; // @[RegFile.scala 97:16:@41866.4]
  assign rport_io_ins_62 = regs_62_io_out; // @[RegFile.scala 97:16:@41867.4]
  assign rport_io_ins_63 = regs_63_io_out; // @[RegFile.scala 97:16:@41868.4]
  assign rport_io_ins_64 = regs_64_io_out; // @[RegFile.scala 97:16:@41869.4]
  assign rport_io_ins_65 = regs_65_io_out; // @[RegFile.scala 97:16:@41870.4]
  assign rport_io_ins_66 = regs_66_io_out; // @[RegFile.scala 97:16:@41871.4]
  assign rport_io_ins_67 = regs_67_io_out; // @[RegFile.scala 97:16:@41872.4]
  assign rport_io_ins_68 = regs_68_io_out; // @[RegFile.scala 97:16:@41873.4]
  assign rport_io_ins_69 = regs_69_io_out; // @[RegFile.scala 97:16:@41874.4]
  assign rport_io_ins_70 = regs_70_io_out; // @[RegFile.scala 97:16:@41875.4]
  assign rport_io_ins_71 = regs_71_io_out; // @[RegFile.scala 97:16:@41876.4]
  assign rport_io_ins_72 = regs_72_io_out; // @[RegFile.scala 97:16:@41877.4]
  assign rport_io_ins_73 = regs_73_io_out; // @[RegFile.scala 97:16:@41878.4]
  assign rport_io_ins_74 = regs_74_io_out; // @[RegFile.scala 97:16:@41879.4]
  assign rport_io_ins_75 = regs_75_io_out; // @[RegFile.scala 97:16:@41880.4]
  assign rport_io_ins_76 = regs_76_io_out; // @[RegFile.scala 97:16:@41881.4]
  assign rport_io_ins_77 = regs_77_io_out; // @[RegFile.scala 97:16:@41882.4]
  assign rport_io_ins_78 = regs_78_io_out; // @[RegFile.scala 97:16:@41883.4]
  assign rport_io_ins_79 = regs_79_io_out; // @[RegFile.scala 97:16:@41884.4]
  assign rport_io_ins_80 = regs_80_io_out; // @[RegFile.scala 97:16:@41885.4]
  assign rport_io_ins_81 = regs_81_io_out; // @[RegFile.scala 97:16:@41886.4]
  assign rport_io_ins_82 = regs_82_io_out; // @[RegFile.scala 97:16:@41887.4]
  assign rport_io_ins_83 = regs_83_io_out; // @[RegFile.scala 97:16:@41888.4]
  assign rport_io_ins_84 = regs_84_io_out; // @[RegFile.scala 97:16:@41889.4]
  assign rport_io_ins_85 = regs_85_io_out; // @[RegFile.scala 97:16:@41890.4]
  assign rport_io_ins_86 = regs_86_io_out; // @[RegFile.scala 97:16:@41891.4]
  assign rport_io_ins_87 = regs_87_io_out; // @[RegFile.scala 97:16:@41892.4]
  assign rport_io_ins_88 = regs_88_io_out; // @[RegFile.scala 97:16:@41893.4]
  assign rport_io_ins_89 = regs_89_io_out; // @[RegFile.scala 97:16:@41894.4]
  assign rport_io_ins_90 = regs_90_io_out; // @[RegFile.scala 97:16:@41895.4]
  assign rport_io_ins_91 = regs_91_io_out; // @[RegFile.scala 97:16:@41896.4]
  assign rport_io_ins_92 = regs_92_io_out; // @[RegFile.scala 97:16:@41897.4]
  assign rport_io_ins_93 = regs_93_io_out; // @[RegFile.scala 97:16:@41898.4]
  assign rport_io_ins_94 = regs_94_io_out; // @[RegFile.scala 97:16:@41899.4]
  assign rport_io_ins_95 = regs_95_io_out; // @[RegFile.scala 97:16:@41900.4]
  assign rport_io_ins_96 = regs_96_io_out; // @[RegFile.scala 97:16:@41901.4]
  assign rport_io_ins_97 = regs_97_io_out; // @[RegFile.scala 97:16:@41902.4]
  assign rport_io_ins_98 = regs_98_io_out; // @[RegFile.scala 97:16:@41903.4]
  assign rport_io_ins_99 = regs_99_io_out; // @[RegFile.scala 97:16:@41904.4]
  assign rport_io_ins_100 = regs_100_io_out; // @[RegFile.scala 97:16:@41905.4]
  assign rport_io_ins_101 = regs_101_io_out; // @[RegFile.scala 97:16:@41906.4]
  assign rport_io_ins_102 = regs_102_io_out; // @[RegFile.scala 97:16:@41907.4]
  assign rport_io_ins_103 = regs_103_io_out; // @[RegFile.scala 97:16:@41908.4]
  assign rport_io_ins_104 = regs_104_io_out; // @[RegFile.scala 97:16:@41909.4]
  assign rport_io_ins_105 = regs_105_io_out; // @[RegFile.scala 97:16:@41910.4]
  assign rport_io_ins_106 = regs_106_io_out; // @[RegFile.scala 97:16:@41911.4]
  assign rport_io_ins_107 = regs_107_io_out; // @[RegFile.scala 97:16:@41912.4]
  assign rport_io_ins_108 = regs_108_io_out; // @[RegFile.scala 97:16:@41913.4]
  assign rport_io_ins_109 = regs_109_io_out; // @[RegFile.scala 97:16:@41914.4]
  assign rport_io_ins_110 = regs_110_io_out; // @[RegFile.scala 97:16:@41915.4]
  assign rport_io_ins_111 = regs_111_io_out; // @[RegFile.scala 97:16:@41916.4]
  assign rport_io_ins_112 = regs_112_io_out; // @[RegFile.scala 97:16:@41917.4]
  assign rport_io_ins_113 = regs_113_io_out; // @[RegFile.scala 97:16:@41918.4]
  assign rport_io_ins_114 = regs_114_io_out; // @[RegFile.scala 97:16:@41919.4]
  assign rport_io_ins_115 = regs_115_io_out; // @[RegFile.scala 97:16:@41920.4]
  assign rport_io_ins_116 = regs_116_io_out; // @[RegFile.scala 97:16:@41921.4]
  assign rport_io_ins_117 = regs_117_io_out; // @[RegFile.scala 97:16:@41922.4]
  assign rport_io_ins_118 = regs_118_io_out; // @[RegFile.scala 97:16:@41923.4]
  assign rport_io_ins_119 = regs_119_io_out; // @[RegFile.scala 97:16:@41924.4]
  assign rport_io_ins_120 = regs_120_io_out; // @[RegFile.scala 97:16:@41925.4]
  assign rport_io_ins_121 = regs_121_io_out; // @[RegFile.scala 97:16:@41926.4]
  assign rport_io_ins_122 = regs_122_io_out; // @[RegFile.scala 97:16:@41927.4]
  assign rport_io_ins_123 = regs_123_io_out; // @[RegFile.scala 97:16:@41928.4]
  assign rport_io_ins_124 = regs_124_io_out; // @[RegFile.scala 97:16:@41929.4]
  assign rport_io_ins_125 = regs_125_io_out; // @[RegFile.scala 97:16:@41930.4]
  assign rport_io_ins_126 = regs_126_io_out; // @[RegFile.scala 97:16:@41931.4]
  assign rport_io_ins_127 = regs_127_io_out; // @[RegFile.scala 97:16:@41932.4]
  assign rport_io_ins_128 = regs_128_io_out; // @[RegFile.scala 97:16:@41933.4]
  assign rport_io_ins_129 = regs_129_io_out; // @[RegFile.scala 97:16:@41934.4]
  assign rport_io_ins_130 = regs_130_io_out; // @[RegFile.scala 97:16:@41935.4]
  assign rport_io_ins_131 = regs_131_io_out; // @[RegFile.scala 97:16:@41936.4]
  assign rport_io_ins_132 = regs_132_io_out; // @[RegFile.scala 97:16:@41937.4]
  assign rport_io_ins_133 = regs_133_io_out; // @[RegFile.scala 97:16:@41938.4]
  assign rport_io_ins_134 = regs_134_io_out; // @[RegFile.scala 97:16:@41939.4]
  assign rport_io_ins_135 = regs_135_io_out; // @[RegFile.scala 97:16:@41940.4]
  assign rport_io_ins_136 = regs_136_io_out; // @[RegFile.scala 97:16:@41941.4]
  assign rport_io_ins_137 = regs_137_io_out; // @[RegFile.scala 97:16:@41942.4]
  assign rport_io_ins_138 = regs_138_io_out; // @[RegFile.scala 97:16:@41943.4]
  assign rport_io_ins_139 = regs_139_io_out; // @[RegFile.scala 97:16:@41944.4]
  assign rport_io_ins_140 = regs_140_io_out; // @[RegFile.scala 97:16:@41945.4]
  assign rport_io_ins_141 = regs_141_io_out; // @[RegFile.scala 97:16:@41946.4]
  assign rport_io_ins_142 = regs_142_io_out; // @[RegFile.scala 97:16:@41947.4]
  assign rport_io_ins_143 = regs_143_io_out; // @[RegFile.scala 97:16:@41948.4]
  assign rport_io_ins_144 = regs_144_io_out; // @[RegFile.scala 97:16:@41949.4]
  assign rport_io_ins_145 = regs_145_io_out; // @[RegFile.scala 97:16:@41950.4]
  assign rport_io_ins_146 = regs_146_io_out; // @[RegFile.scala 97:16:@41951.4]
  assign rport_io_ins_147 = regs_147_io_out; // @[RegFile.scala 97:16:@41952.4]
  assign rport_io_ins_148 = regs_148_io_out; // @[RegFile.scala 97:16:@41953.4]
  assign rport_io_ins_149 = regs_149_io_out; // @[RegFile.scala 97:16:@41954.4]
  assign rport_io_ins_150 = regs_150_io_out; // @[RegFile.scala 97:16:@41955.4]
  assign rport_io_ins_151 = regs_151_io_out; // @[RegFile.scala 97:16:@41956.4]
  assign rport_io_ins_152 = regs_152_io_out; // @[RegFile.scala 97:16:@41957.4]
  assign rport_io_ins_153 = regs_153_io_out; // @[RegFile.scala 97:16:@41958.4]
  assign rport_io_ins_154 = regs_154_io_out; // @[RegFile.scala 97:16:@41959.4]
  assign rport_io_ins_155 = regs_155_io_out; // @[RegFile.scala 97:16:@41960.4]
  assign rport_io_ins_156 = regs_156_io_out; // @[RegFile.scala 97:16:@41961.4]
  assign rport_io_ins_157 = regs_157_io_out; // @[RegFile.scala 97:16:@41962.4]
  assign rport_io_ins_158 = regs_158_io_out; // @[RegFile.scala 97:16:@41963.4]
  assign rport_io_ins_159 = regs_159_io_out; // @[RegFile.scala 97:16:@41964.4]
  assign rport_io_ins_160 = regs_160_io_out; // @[RegFile.scala 97:16:@41965.4]
  assign rport_io_ins_161 = regs_161_io_out; // @[RegFile.scala 97:16:@41966.4]
  assign rport_io_ins_162 = regs_162_io_out; // @[RegFile.scala 97:16:@41967.4]
  assign rport_io_ins_163 = regs_163_io_out; // @[RegFile.scala 97:16:@41968.4]
  assign rport_io_ins_164 = regs_164_io_out; // @[RegFile.scala 97:16:@41969.4]
  assign rport_io_ins_165 = regs_165_io_out; // @[RegFile.scala 97:16:@41970.4]
  assign rport_io_ins_166 = regs_166_io_out; // @[RegFile.scala 97:16:@41971.4]
  assign rport_io_ins_167 = regs_167_io_out; // @[RegFile.scala 97:16:@41972.4]
  assign rport_io_ins_168 = regs_168_io_out; // @[RegFile.scala 97:16:@41973.4]
  assign rport_io_ins_169 = regs_169_io_out; // @[RegFile.scala 97:16:@41974.4]
  assign rport_io_ins_170 = regs_170_io_out; // @[RegFile.scala 97:16:@41975.4]
  assign rport_io_ins_171 = regs_171_io_out; // @[RegFile.scala 97:16:@41976.4]
  assign rport_io_ins_172 = regs_172_io_out; // @[RegFile.scala 97:16:@41977.4]
  assign rport_io_ins_173 = regs_173_io_out; // @[RegFile.scala 97:16:@41978.4]
  assign rport_io_ins_174 = regs_174_io_out; // @[RegFile.scala 97:16:@41979.4]
  assign rport_io_ins_175 = regs_175_io_out; // @[RegFile.scala 97:16:@41980.4]
  assign rport_io_ins_176 = regs_176_io_out; // @[RegFile.scala 97:16:@41981.4]
  assign rport_io_ins_177 = regs_177_io_out; // @[RegFile.scala 97:16:@41982.4]
  assign rport_io_ins_178 = regs_178_io_out; // @[RegFile.scala 97:16:@41983.4]
  assign rport_io_ins_179 = regs_179_io_out; // @[RegFile.scala 97:16:@41984.4]
  assign rport_io_ins_180 = regs_180_io_out; // @[RegFile.scala 97:16:@41985.4]
  assign rport_io_ins_181 = regs_181_io_out; // @[RegFile.scala 97:16:@41986.4]
  assign rport_io_ins_182 = regs_182_io_out; // @[RegFile.scala 97:16:@41987.4]
  assign rport_io_ins_183 = regs_183_io_out; // @[RegFile.scala 97:16:@41988.4]
  assign rport_io_ins_184 = regs_184_io_out; // @[RegFile.scala 97:16:@41989.4]
  assign rport_io_ins_185 = regs_185_io_out; // @[RegFile.scala 97:16:@41990.4]
  assign rport_io_ins_186 = regs_186_io_out; // @[RegFile.scala 97:16:@41991.4]
  assign rport_io_ins_187 = regs_187_io_out; // @[RegFile.scala 97:16:@41992.4]
  assign rport_io_ins_188 = regs_188_io_out; // @[RegFile.scala 97:16:@41993.4]
  assign rport_io_ins_189 = regs_189_io_out; // @[RegFile.scala 97:16:@41994.4]
  assign rport_io_ins_190 = regs_190_io_out; // @[RegFile.scala 97:16:@41995.4]
  assign rport_io_ins_191 = regs_191_io_out; // @[RegFile.scala 97:16:@41996.4]
  assign rport_io_ins_192 = regs_192_io_out; // @[RegFile.scala 97:16:@41997.4]
  assign rport_io_ins_193 = regs_193_io_out; // @[RegFile.scala 97:16:@41998.4]
  assign rport_io_ins_194 = regs_194_io_out; // @[RegFile.scala 97:16:@41999.4]
  assign rport_io_ins_195 = regs_195_io_out; // @[RegFile.scala 97:16:@42000.4]
  assign rport_io_ins_196 = regs_196_io_out; // @[RegFile.scala 97:16:@42001.4]
  assign rport_io_ins_197 = regs_197_io_out; // @[RegFile.scala 97:16:@42002.4]
  assign rport_io_ins_198 = regs_198_io_out; // @[RegFile.scala 97:16:@42003.4]
  assign rport_io_ins_199 = regs_199_io_out; // @[RegFile.scala 97:16:@42004.4]
  assign rport_io_ins_200 = regs_200_io_out; // @[RegFile.scala 97:16:@42005.4]
  assign rport_io_ins_201 = regs_201_io_out; // @[RegFile.scala 97:16:@42006.4]
  assign rport_io_ins_202 = regs_202_io_out; // @[RegFile.scala 97:16:@42007.4]
  assign rport_io_ins_203 = regs_203_io_out; // @[RegFile.scala 97:16:@42008.4]
  assign rport_io_ins_204 = regs_204_io_out; // @[RegFile.scala 97:16:@42009.4]
  assign rport_io_ins_205 = regs_205_io_out; // @[RegFile.scala 97:16:@42010.4]
  assign rport_io_ins_206 = regs_206_io_out; // @[RegFile.scala 97:16:@42011.4]
  assign rport_io_ins_207 = regs_207_io_out; // @[RegFile.scala 97:16:@42012.4]
  assign rport_io_ins_208 = regs_208_io_out; // @[RegFile.scala 97:16:@42013.4]
  assign rport_io_ins_209 = regs_209_io_out; // @[RegFile.scala 97:16:@42014.4]
  assign rport_io_ins_210 = regs_210_io_out; // @[RegFile.scala 97:16:@42015.4]
  assign rport_io_ins_211 = regs_211_io_out; // @[RegFile.scala 97:16:@42016.4]
  assign rport_io_ins_212 = regs_212_io_out; // @[RegFile.scala 97:16:@42017.4]
  assign rport_io_ins_213 = regs_213_io_out; // @[RegFile.scala 97:16:@42018.4]
  assign rport_io_ins_214 = regs_214_io_out; // @[RegFile.scala 97:16:@42019.4]
  assign rport_io_ins_215 = regs_215_io_out; // @[RegFile.scala 97:16:@42020.4]
  assign rport_io_ins_216 = regs_216_io_out; // @[RegFile.scala 97:16:@42021.4]
  assign rport_io_ins_217 = regs_217_io_out; // @[RegFile.scala 97:16:@42022.4]
  assign rport_io_ins_218 = regs_218_io_out; // @[RegFile.scala 97:16:@42023.4]
  assign rport_io_ins_219 = regs_219_io_out; // @[RegFile.scala 97:16:@42024.4]
  assign rport_io_ins_220 = regs_220_io_out; // @[RegFile.scala 97:16:@42025.4]
  assign rport_io_ins_221 = regs_221_io_out; // @[RegFile.scala 97:16:@42026.4]
  assign rport_io_ins_222 = regs_222_io_out; // @[RegFile.scala 97:16:@42027.4]
  assign rport_io_ins_223 = regs_223_io_out; // @[RegFile.scala 97:16:@42028.4]
  assign rport_io_ins_224 = regs_224_io_out; // @[RegFile.scala 97:16:@42029.4]
  assign rport_io_ins_225 = regs_225_io_out; // @[RegFile.scala 97:16:@42030.4]
  assign rport_io_ins_226 = regs_226_io_out; // @[RegFile.scala 97:16:@42031.4]
  assign rport_io_ins_227 = regs_227_io_out; // @[RegFile.scala 97:16:@42032.4]
  assign rport_io_ins_228 = regs_228_io_out; // @[RegFile.scala 97:16:@42033.4]
  assign rport_io_ins_229 = regs_229_io_out; // @[RegFile.scala 97:16:@42034.4]
  assign rport_io_ins_230 = regs_230_io_out; // @[RegFile.scala 97:16:@42035.4]
  assign rport_io_ins_231 = regs_231_io_out; // @[RegFile.scala 97:16:@42036.4]
  assign rport_io_ins_232 = regs_232_io_out; // @[RegFile.scala 97:16:@42037.4]
  assign rport_io_ins_233 = regs_233_io_out; // @[RegFile.scala 97:16:@42038.4]
  assign rport_io_ins_234 = regs_234_io_out; // @[RegFile.scala 97:16:@42039.4]
  assign rport_io_ins_235 = regs_235_io_out; // @[RegFile.scala 97:16:@42040.4]
  assign rport_io_ins_236 = regs_236_io_out; // @[RegFile.scala 97:16:@42041.4]
  assign rport_io_ins_237 = regs_237_io_out; // @[RegFile.scala 97:16:@42042.4]
  assign rport_io_ins_238 = regs_238_io_out; // @[RegFile.scala 97:16:@42043.4]
  assign rport_io_ins_239 = regs_239_io_out; // @[RegFile.scala 97:16:@42044.4]
  assign rport_io_ins_240 = regs_240_io_out; // @[RegFile.scala 97:16:@42045.4]
  assign rport_io_ins_241 = regs_241_io_out; // @[RegFile.scala 97:16:@42046.4]
  assign rport_io_ins_242 = regs_242_io_out; // @[RegFile.scala 97:16:@42047.4]
  assign rport_io_ins_243 = regs_243_io_out; // @[RegFile.scala 97:16:@42048.4]
  assign rport_io_ins_244 = regs_244_io_out; // @[RegFile.scala 97:16:@42049.4]
  assign rport_io_ins_245 = regs_245_io_out; // @[RegFile.scala 97:16:@42050.4]
  assign rport_io_ins_246 = regs_246_io_out; // @[RegFile.scala 97:16:@42051.4]
  assign rport_io_ins_247 = regs_247_io_out; // @[RegFile.scala 97:16:@42052.4]
  assign rport_io_ins_248 = regs_248_io_out; // @[RegFile.scala 97:16:@42053.4]
  assign rport_io_ins_249 = regs_249_io_out; // @[RegFile.scala 97:16:@42054.4]
  assign rport_io_ins_250 = regs_250_io_out; // @[RegFile.scala 97:16:@42055.4]
  assign rport_io_ins_251 = regs_251_io_out; // @[RegFile.scala 97:16:@42056.4]
  assign rport_io_ins_252 = regs_252_io_out; // @[RegFile.scala 97:16:@42057.4]
  assign rport_io_ins_253 = regs_253_io_out; // @[RegFile.scala 97:16:@42058.4]
  assign rport_io_ins_254 = regs_254_io_out; // @[RegFile.scala 97:16:@42059.4]
  assign rport_io_ins_255 = regs_255_io_out; // @[RegFile.scala 97:16:@42060.4]
  assign rport_io_ins_256 = regs_256_io_out; // @[RegFile.scala 97:16:@42061.4]
  assign rport_io_ins_257 = regs_257_io_out; // @[RegFile.scala 97:16:@42062.4]
  assign rport_io_ins_258 = regs_258_io_out; // @[RegFile.scala 97:16:@42063.4]
  assign rport_io_ins_259 = regs_259_io_out; // @[RegFile.scala 97:16:@42064.4]
  assign rport_io_ins_260 = regs_260_io_out; // @[RegFile.scala 97:16:@42065.4]
  assign rport_io_ins_261 = regs_261_io_out; // @[RegFile.scala 97:16:@42066.4]
  assign rport_io_ins_262 = regs_262_io_out; // @[RegFile.scala 97:16:@42067.4]
  assign rport_io_ins_263 = regs_263_io_out; // @[RegFile.scala 97:16:@42068.4]
  assign rport_io_ins_264 = regs_264_io_out; // @[RegFile.scala 97:16:@42069.4]
  assign rport_io_ins_265 = regs_265_io_out; // @[RegFile.scala 97:16:@42070.4]
  assign rport_io_ins_266 = regs_266_io_out; // @[RegFile.scala 97:16:@42071.4]
  assign rport_io_ins_267 = regs_267_io_out; // @[RegFile.scala 97:16:@42072.4]
  assign rport_io_ins_268 = regs_268_io_out; // @[RegFile.scala 97:16:@42073.4]
  assign rport_io_ins_269 = regs_269_io_out; // @[RegFile.scala 97:16:@42074.4]
  assign rport_io_ins_270 = regs_270_io_out; // @[RegFile.scala 97:16:@42075.4]
  assign rport_io_ins_271 = regs_271_io_out; // @[RegFile.scala 97:16:@42076.4]
  assign rport_io_ins_272 = regs_272_io_out; // @[RegFile.scala 97:16:@42077.4]
  assign rport_io_ins_273 = regs_273_io_out; // @[RegFile.scala 97:16:@42078.4]
  assign rport_io_ins_274 = regs_274_io_out; // @[RegFile.scala 97:16:@42079.4]
  assign rport_io_ins_275 = regs_275_io_out; // @[RegFile.scala 97:16:@42080.4]
  assign rport_io_ins_276 = regs_276_io_out; // @[RegFile.scala 97:16:@42081.4]
  assign rport_io_ins_277 = regs_277_io_out; // @[RegFile.scala 97:16:@42082.4]
  assign rport_io_ins_278 = regs_278_io_out; // @[RegFile.scala 97:16:@42083.4]
  assign rport_io_ins_279 = regs_279_io_out; // @[RegFile.scala 97:16:@42084.4]
  assign rport_io_ins_280 = regs_280_io_out; // @[RegFile.scala 97:16:@42085.4]
  assign rport_io_ins_281 = regs_281_io_out; // @[RegFile.scala 97:16:@42086.4]
  assign rport_io_ins_282 = regs_282_io_out; // @[RegFile.scala 97:16:@42087.4]
  assign rport_io_ins_283 = regs_283_io_out; // @[RegFile.scala 97:16:@42088.4]
  assign rport_io_ins_284 = regs_284_io_out; // @[RegFile.scala 97:16:@42089.4]
  assign rport_io_ins_285 = regs_285_io_out; // @[RegFile.scala 97:16:@42090.4]
  assign rport_io_ins_286 = regs_286_io_out; // @[RegFile.scala 97:16:@42091.4]
  assign rport_io_ins_287 = regs_287_io_out; // @[RegFile.scala 97:16:@42092.4]
  assign rport_io_ins_288 = regs_288_io_out; // @[RegFile.scala 97:16:@42093.4]
  assign rport_io_ins_289 = regs_289_io_out; // @[RegFile.scala 97:16:@42094.4]
  assign rport_io_ins_290 = regs_290_io_out; // @[RegFile.scala 97:16:@42095.4]
  assign rport_io_ins_291 = regs_291_io_out; // @[RegFile.scala 97:16:@42096.4]
  assign rport_io_ins_292 = regs_292_io_out; // @[RegFile.scala 97:16:@42097.4]
  assign rport_io_ins_293 = regs_293_io_out; // @[RegFile.scala 97:16:@42098.4]
  assign rport_io_ins_294 = regs_294_io_out; // @[RegFile.scala 97:16:@42099.4]
  assign rport_io_ins_295 = regs_295_io_out; // @[RegFile.scala 97:16:@42100.4]
  assign rport_io_ins_296 = regs_296_io_out; // @[RegFile.scala 97:16:@42101.4]
  assign rport_io_ins_297 = regs_297_io_out; // @[RegFile.scala 97:16:@42102.4]
  assign rport_io_ins_298 = regs_298_io_out; // @[RegFile.scala 97:16:@42103.4]
  assign rport_io_ins_299 = regs_299_io_out; // @[RegFile.scala 97:16:@42104.4]
  assign rport_io_ins_300 = regs_300_io_out; // @[RegFile.scala 97:16:@42105.4]
  assign rport_io_ins_301 = regs_301_io_out; // @[RegFile.scala 97:16:@42106.4]
  assign rport_io_ins_302 = regs_302_io_out; // @[RegFile.scala 97:16:@42107.4]
  assign rport_io_ins_303 = regs_303_io_out; // @[RegFile.scala 97:16:@42108.4]
  assign rport_io_ins_304 = regs_304_io_out; // @[RegFile.scala 97:16:@42109.4]
  assign rport_io_ins_305 = regs_305_io_out; // @[RegFile.scala 97:16:@42110.4]
  assign rport_io_ins_306 = regs_306_io_out; // @[RegFile.scala 97:16:@42111.4]
  assign rport_io_ins_307 = regs_307_io_out; // @[RegFile.scala 97:16:@42112.4]
  assign rport_io_ins_308 = regs_308_io_out; // @[RegFile.scala 97:16:@42113.4]
  assign rport_io_ins_309 = regs_309_io_out; // @[RegFile.scala 97:16:@42114.4]
  assign rport_io_ins_310 = regs_310_io_out; // @[RegFile.scala 97:16:@42115.4]
  assign rport_io_ins_311 = regs_311_io_out; // @[RegFile.scala 97:16:@42116.4]
  assign rport_io_ins_312 = regs_312_io_out; // @[RegFile.scala 97:16:@42117.4]
  assign rport_io_ins_313 = regs_313_io_out; // @[RegFile.scala 97:16:@42118.4]
  assign rport_io_ins_314 = regs_314_io_out; // @[RegFile.scala 97:16:@42119.4]
  assign rport_io_ins_315 = regs_315_io_out; // @[RegFile.scala 97:16:@42120.4]
  assign rport_io_ins_316 = regs_316_io_out; // @[RegFile.scala 97:16:@42121.4]
  assign rport_io_ins_317 = regs_317_io_out; // @[RegFile.scala 97:16:@42122.4]
  assign rport_io_ins_318 = regs_318_io_out; // @[RegFile.scala 97:16:@42123.4]
  assign rport_io_ins_319 = regs_319_io_out; // @[RegFile.scala 97:16:@42124.4]
  assign rport_io_ins_320 = regs_320_io_out; // @[RegFile.scala 97:16:@42125.4]
  assign rport_io_ins_321 = regs_321_io_out; // @[RegFile.scala 97:16:@42126.4]
  assign rport_io_ins_322 = regs_322_io_out; // @[RegFile.scala 97:16:@42127.4]
  assign rport_io_ins_323 = regs_323_io_out; // @[RegFile.scala 97:16:@42128.4]
  assign rport_io_ins_324 = regs_324_io_out; // @[RegFile.scala 97:16:@42129.4]
  assign rport_io_ins_325 = regs_325_io_out; // @[RegFile.scala 97:16:@42130.4]
  assign rport_io_ins_326 = regs_326_io_out; // @[RegFile.scala 97:16:@42131.4]
  assign rport_io_ins_327 = regs_327_io_out; // @[RegFile.scala 97:16:@42132.4]
  assign rport_io_ins_328 = regs_328_io_out; // @[RegFile.scala 97:16:@42133.4]
  assign rport_io_ins_329 = regs_329_io_out; // @[RegFile.scala 97:16:@42134.4]
  assign rport_io_ins_330 = regs_330_io_out; // @[RegFile.scala 97:16:@42135.4]
  assign rport_io_ins_331 = regs_331_io_out; // @[RegFile.scala 97:16:@42136.4]
  assign rport_io_ins_332 = regs_332_io_out; // @[RegFile.scala 97:16:@42137.4]
  assign rport_io_ins_333 = regs_333_io_out; // @[RegFile.scala 97:16:@42138.4]
  assign rport_io_ins_334 = regs_334_io_out; // @[RegFile.scala 97:16:@42139.4]
  assign rport_io_ins_335 = regs_335_io_out; // @[RegFile.scala 97:16:@42140.4]
  assign rport_io_ins_336 = regs_336_io_out; // @[RegFile.scala 97:16:@42141.4]
  assign rport_io_ins_337 = regs_337_io_out; // @[RegFile.scala 97:16:@42142.4]
  assign rport_io_ins_338 = regs_338_io_out; // @[RegFile.scala 97:16:@42143.4]
  assign rport_io_ins_339 = regs_339_io_out; // @[RegFile.scala 97:16:@42144.4]
  assign rport_io_ins_340 = regs_340_io_out; // @[RegFile.scala 97:16:@42145.4]
  assign rport_io_ins_341 = regs_341_io_out; // @[RegFile.scala 97:16:@42146.4]
  assign rport_io_ins_342 = regs_342_io_out; // @[RegFile.scala 97:16:@42147.4]
  assign rport_io_ins_343 = regs_343_io_out; // @[RegFile.scala 97:16:@42148.4]
  assign rport_io_ins_344 = regs_344_io_out; // @[RegFile.scala 97:16:@42149.4]
  assign rport_io_ins_345 = regs_345_io_out; // @[RegFile.scala 97:16:@42150.4]
  assign rport_io_ins_346 = regs_346_io_out; // @[RegFile.scala 97:16:@42151.4]
  assign rport_io_ins_347 = regs_347_io_out; // @[RegFile.scala 97:16:@42152.4]
  assign rport_io_ins_348 = regs_348_io_out; // @[RegFile.scala 97:16:@42153.4]
  assign rport_io_ins_349 = regs_349_io_out; // @[RegFile.scala 97:16:@42154.4]
  assign rport_io_ins_350 = regs_350_io_out; // @[RegFile.scala 97:16:@42155.4]
  assign rport_io_ins_351 = regs_351_io_out; // @[RegFile.scala 97:16:@42156.4]
  assign rport_io_ins_352 = regs_352_io_out; // @[RegFile.scala 97:16:@42157.4]
  assign rport_io_ins_353 = regs_353_io_out; // @[RegFile.scala 97:16:@42158.4]
  assign rport_io_ins_354 = regs_354_io_out; // @[RegFile.scala 97:16:@42159.4]
  assign rport_io_ins_355 = regs_355_io_out; // @[RegFile.scala 97:16:@42160.4]
  assign rport_io_ins_356 = regs_356_io_out; // @[RegFile.scala 97:16:@42161.4]
  assign rport_io_ins_357 = regs_357_io_out; // @[RegFile.scala 97:16:@42162.4]
  assign rport_io_ins_358 = regs_358_io_out; // @[RegFile.scala 97:16:@42163.4]
  assign rport_io_ins_359 = regs_359_io_out; // @[RegFile.scala 97:16:@42164.4]
  assign rport_io_ins_360 = regs_360_io_out; // @[RegFile.scala 97:16:@42165.4]
  assign rport_io_ins_361 = regs_361_io_out; // @[RegFile.scala 97:16:@42166.4]
  assign rport_io_ins_362 = regs_362_io_out; // @[RegFile.scala 97:16:@42167.4]
  assign rport_io_ins_363 = regs_363_io_out; // @[RegFile.scala 97:16:@42168.4]
  assign rport_io_ins_364 = regs_364_io_out; // @[RegFile.scala 97:16:@42169.4]
  assign rport_io_ins_365 = regs_365_io_out; // @[RegFile.scala 97:16:@42170.4]
  assign rport_io_ins_366 = regs_366_io_out; // @[RegFile.scala 97:16:@42171.4]
  assign rport_io_ins_367 = regs_367_io_out; // @[RegFile.scala 97:16:@42172.4]
  assign rport_io_ins_368 = regs_368_io_out; // @[RegFile.scala 97:16:@42173.4]
  assign rport_io_ins_369 = regs_369_io_out; // @[RegFile.scala 97:16:@42174.4]
  assign rport_io_ins_370 = regs_370_io_out; // @[RegFile.scala 97:16:@42175.4]
  assign rport_io_ins_371 = regs_371_io_out; // @[RegFile.scala 97:16:@42176.4]
  assign rport_io_ins_372 = regs_372_io_out; // @[RegFile.scala 97:16:@42177.4]
  assign rport_io_ins_373 = regs_373_io_out; // @[RegFile.scala 97:16:@42178.4]
  assign rport_io_ins_374 = regs_374_io_out; // @[RegFile.scala 97:16:@42179.4]
  assign rport_io_ins_375 = regs_375_io_out; // @[RegFile.scala 97:16:@42180.4]
  assign rport_io_ins_376 = regs_376_io_out; // @[RegFile.scala 97:16:@42181.4]
  assign rport_io_ins_377 = regs_377_io_out; // @[RegFile.scala 97:16:@42182.4]
  assign rport_io_ins_378 = regs_378_io_out; // @[RegFile.scala 97:16:@42183.4]
  assign rport_io_ins_379 = regs_379_io_out; // @[RegFile.scala 97:16:@42184.4]
  assign rport_io_ins_380 = regs_380_io_out; // @[RegFile.scala 97:16:@42185.4]
  assign rport_io_ins_381 = regs_381_io_out; // @[RegFile.scala 97:16:@42186.4]
  assign rport_io_ins_382 = regs_382_io_out; // @[RegFile.scala 97:16:@42187.4]
  assign rport_io_ins_383 = regs_383_io_out; // @[RegFile.scala 97:16:@42188.4]
  assign rport_io_ins_384 = regs_384_io_out; // @[RegFile.scala 97:16:@42189.4]
  assign rport_io_ins_385 = regs_385_io_out; // @[RegFile.scala 97:16:@42190.4]
  assign rport_io_ins_386 = regs_386_io_out; // @[RegFile.scala 97:16:@42191.4]
  assign rport_io_ins_387 = regs_387_io_out; // @[RegFile.scala 97:16:@42192.4]
  assign rport_io_ins_388 = regs_388_io_out; // @[RegFile.scala 97:16:@42193.4]
  assign rport_io_ins_389 = regs_389_io_out; // @[RegFile.scala 97:16:@42194.4]
  assign rport_io_ins_390 = regs_390_io_out; // @[RegFile.scala 97:16:@42195.4]
  assign rport_io_ins_391 = regs_391_io_out; // @[RegFile.scala 97:16:@42196.4]
  assign rport_io_ins_392 = regs_392_io_out; // @[RegFile.scala 97:16:@42197.4]
  assign rport_io_ins_393 = regs_393_io_out; // @[RegFile.scala 97:16:@42198.4]
  assign rport_io_ins_394 = regs_394_io_out; // @[RegFile.scala 97:16:@42199.4]
  assign rport_io_ins_395 = regs_395_io_out; // @[RegFile.scala 97:16:@42200.4]
  assign rport_io_ins_396 = regs_396_io_out; // @[RegFile.scala 97:16:@42201.4]
  assign rport_io_ins_397 = regs_397_io_out; // @[RegFile.scala 97:16:@42202.4]
  assign rport_io_ins_398 = regs_398_io_out; // @[RegFile.scala 97:16:@42203.4]
  assign rport_io_ins_399 = regs_399_io_out; // @[RegFile.scala 97:16:@42204.4]
  assign rport_io_ins_400 = regs_400_io_out; // @[RegFile.scala 97:16:@42205.4]
  assign rport_io_ins_401 = regs_401_io_out; // @[RegFile.scala 97:16:@42206.4]
  assign rport_io_ins_402 = regs_402_io_out; // @[RegFile.scala 97:16:@42207.4]
  assign rport_io_ins_403 = regs_403_io_out; // @[RegFile.scala 97:16:@42208.4]
  assign rport_io_ins_404 = regs_404_io_out; // @[RegFile.scala 97:16:@42209.4]
  assign rport_io_ins_405 = regs_405_io_out; // @[RegFile.scala 97:16:@42210.4]
  assign rport_io_ins_406 = regs_406_io_out; // @[RegFile.scala 97:16:@42211.4]
  assign rport_io_ins_407 = regs_407_io_out; // @[RegFile.scala 97:16:@42212.4]
  assign rport_io_ins_408 = regs_408_io_out; // @[RegFile.scala 97:16:@42213.4]
  assign rport_io_ins_409 = regs_409_io_out; // @[RegFile.scala 97:16:@42214.4]
  assign rport_io_ins_410 = regs_410_io_out; // @[RegFile.scala 97:16:@42215.4]
  assign rport_io_ins_411 = regs_411_io_out; // @[RegFile.scala 97:16:@42216.4]
  assign rport_io_ins_412 = regs_412_io_out; // @[RegFile.scala 97:16:@42217.4]
  assign rport_io_ins_413 = regs_413_io_out; // @[RegFile.scala 97:16:@42218.4]
  assign rport_io_ins_414 = regs_414_io_out; // @[RegFile.scala 97:16:@42219.4]
  assign rport_io_ins_415 = regs_415_io_out; // @[RegFile.scala 97:16:@42220.4]
  assign rport_io_ins_416 = regs_416_io_out; // @[RegFile.scala 97:16:@42221.4]
  assign rport_io_ins_417 = regs_417_io_out; // @[RegFile.scala 97:16:@42222.4]
  assign rport_io_ins_418 = regs_418_io_out; // @[RegFile.scala 97:16:@42223.4]
  assign rport_io_ins_419 = regs_419_io_out; // @[RegFile.scala 97:16:@42224.4]
  assign rport_io_ins_420 = regs_420_io_out; // @[RegFile.scala 97:16:@42225.4]
  assign rport_io_ins_421 = regs_421_io_out; // @[RegFile.scala 97:16:@42226.4]
  assign rport_io_ins_422 = regs_422_io_out; // @[RegFile.scala 97:16:@42227.4]
  assign rport_io_ins_423 = regs_423_io_out; // @[RegFile.scala 97:16:@42228.4]
  assign rport_io_ins_424 = regs_424_io_out; // @[RegFile.scala 97:16:@42229.4]
  assign rport_io_ins_425 = regs_425_io_out; // @[RegFile.scala 97:16:@42230.4]
  assign rport_io_ins_426 = regs_426_io_out; // @[RegFile.scala 97:16:@42231.4]
  assign rport_io_ins_427 = regs_427_io_out; // @[RegFile.scala 97:16:@42232.4]
  assign rport_io_ins_428 = regs_428_io_out; // @[RegFile.scala 97:16:@42233.4]
  assign rport_io_ins_429 = regs_429_io_out; // @[RegFile.scala 97:16:@42234.4]
  assign rport_io_ins_430 = regs_430_io_out; // @[RegFile.scala 97:16:@42235.4]
  assign rport_io_ins_431 = regs_431_io_out; // @[RegFile.scala 97:16:@42236.4]
  assign rport_io_ins_432 = regs_432_io_out; // @[RegFile.scala 97:16:@42237.4]
  assign rport_io_ins_433 = regs_433_io_out; // @[RegFile.scala 97:16:@42238.4]
  assign rport_io_ins_434 = regs_434_io_out; // @[RegFile.scala 97:16:@42239.4]
  assign rport_io_ins_435 = regs_435_io_out; // @[RegFile.scala 97:16:@42240.4]
  assign rport_io_ins_436 = regs_436_io_out; // @[RegFile.scala 97:16:@42241.4]
  assign rport_io_ins_437 = regs_437_io_out; // @[RegFile.scala 97:16:@42242.4]
  assign rport_io_ins_438 = regs_438_io_out; // @[RegFile.scala 97:16:@42243.4]
  assign rport_io_ins_439 = regs_439_io_out; // @[RegFile.scala 97:16:@42244.4]
  assign rport_io_ins_440 = regs_440_io_out; // @[RegFile.scala 97:16:@42245.4]
  assign rport_io_ins_441 = regs_441_io_out; // @[RegFile.scala 97:16:@42246.4]
  assign rport_io_ins_442 = regs_442_io_out; // @[RegFile.scala 97:16:@42247.4]
  assign rport_io_ins_443 = regs_443_io_out; // @[RegFile.scala 97:16:@42248.4]
  assign rport_io_ins_444 = regs_444_io_out; // @[RegFile.scala 97:16:@42249.4]
  assign rport_io_ins_445 = regs_445_io_out; // @[RegFile.scala 97:16:@42250.4]
  assign rport_io_ins_446 = regs_446_io_out; // @[RegFile.scala 97:16:@42251.4]
  assign rport_io_ins_447 = regs_447_io_out; // @[RegFile.scala 97:16:@42252.4]
  assign rport_io_ins_448 = regs_448_io_out; // @[RegFile.scala 97:16:@42253.4]
  assign rport_io_ins_449 = regs_449_io_out; // @[RegFile.scala 97:16:@42254.4]
  assign rport_io_ins_450 = regs_450_io_out; // @[RegFile.scala 97:16:@42255.4]
  assign rport_io_ins_451 = regs_451_io_out; // @[RegFile.scala 97:16:@42256.4]
  assign rport_io_ins_452 = regs_452_io_out; // @[RegFile.scala 97:16:@42257.4]
  assign rport_io_ins_453 = regs_453_io_out; // @[RegFile.scala 97:16:@42258.4]
  assign rport_io_ins_454 = regs_454_io_out; // @[RegFile.scala 97:16:@42259.4]
  assign rport_io_ins_455 = regs_455_io_out; // @[RegFile.scala 97:16:@42260.4]
  assign rport_io_ins_456 = regs_456_io_out; // @[RegFile.scala 97:16:@42261.4]
  assign rport_io_ins_457 = regs_457_io_out; // @[RegFile.scala 97:16:@42262.4]
  assign rport_io_ins_458 = regs_458_io_out; // @[RegFile.scala 97:16:@42263.4]
  assign rport_io_ins_459 = regs_459_io_out; // @[RegFile.scala 97:16:@42264.4]
  assign rport_io_ins_460 = regs_460_io_out; // @[RegFile.scala 97:16:@42265.4]
  assign rport_io_ins_461 = regs_461_io_out; // @[RegFile.scala 97:16:@42266.4]
  assign rport_io_ins_462 = regs_462_io_out; // @[RegFile.scala 97:16:@42267.4]
  assign rport_io_ins_463 = regs_463_io_out; // @[RegFile.scala 97:16:@42268.4]
  assign rport_io_ins_464 = regs_464_io_out; // @[RegFile.scala 97:16:@42269.4]
  assign rport_io_ins_465 = regs_465_io_out; // @[RegFile.scala 97:16:@42270.4]
  assign rport_io_ins_466 = regs_466_io_out; // @[RegFile.scala 97:16:@42271.4]
  assign rport_io_ins_467 = regs_467_io_out; // @[RegFile.scala 97:16:@42272.4]
  assign rport_io_ins_468 = regs_468_io_out; // @[RegFile.scala 97:16:@42273.4]
  assign rport_io_ins_469 = regs_469_io_out; // @[RegFile.scala 97:16:@42274.4]
  assign rport_io_ins_470 = regs_470_io_out; // @[RegFile.scala 97:16:@42275.4]
  assign rport_io_ins_471 = regs_471_io_out; // @[RegFile.scala 97:16:@42276.4]
  assign rport_io_ins_472 = regs_472_io_out; // @[RegFile.scala 97:16:@42277.4]
  assign rport_io_ins_473 = regs_473_io_out; // @[RegFile.scala 97:16:@42278.4]
  assign rport_io_ins_474 = regs_474_io_out; // @[RegFile.scala 97:16:@42279.4]
  assign rport_io_ins_475 = regs_475_io_out; // @[RegFile.scala 97:16:@42280.4]
  assign rport_io_ins_476 = regs_476_io_out; // @[RegFile.scala 97:16:@42281.4]
  assign rport_io_ins_477 = regs_477_io_out; // @[RegFile.scala 97:16:@42282.4]
  assign rport_io_ins_478 = regs_478_io_out; // @[RegFile.scala 97:16:@42283.4]
  assign rport_io_ins_479 = regs_479_io_out; // @[RegFile.scala 97:16:@42284.4]
  assign rport_io_ins_480 = regs_480_io_out; // @[RegFile.scala 97:16:@42285.4]
  assign rport_io_ins_481 = regs_481_io_out; // @[RegFile.scala 97:16:@42286.4]
  assign rport_io_ins_482 = regs_482_io_out; // @[RegFile.scala 97:16:@42287.4]
  assign rport_io_ins_483 = regs_483_io_out; // @[RegFile.scala 97:16:@42288.4]
  assign rport_io_ins_484 = regs_484_io_out; // @[RegFile.scala 97:16:@42289.4]
  assign rport_io_ins_485 = regs_485_io_out; // @[RegFile.scala 97:16:@42290.4]
  assign rport_io_ins_486 = regs_486_io_out; // @[RegFile.scala 97:16:@42291.4]
  assign rport_io_ins_487 = regs_487_io_out; // @[RegFile.scala 97:16:@42292.4]
  assign rport_io_ins_488 = regs_488_io_out; // @[RegFile.scala 97:16:@42293.4]
  assign rport_io_ins_489 = regs_489_io_out; // @[RegFile.scala 97:16:@42294.4]
  assign rport_io_ins_490 = regs_490_io_out; // @[RegFile.scala 97:16:@42295.4]
  assign rport_io_ins_491 = regs_491_io_out; // @[RegFile.scala 97:16:@42296.4]
  assign rport_io_ins_492 = regs_492_io_out; // @[RegFile.scala 97:16:@42297.4]
  assign rport_io_ins_493 = regs_493_io_out; // @[RegFile.scala 97:16:@42298.4]
  assign rport_io_ins_494 = regs_494_io_out; // @[RegFile.scala 97:16:@42299.4]
  assign rport_io_ins_495 = regs_495_io_out; // @[RegFile.scala 97:16:@42300.4]
  assign rport_io_ins_496 = regs_496_io_out; // @[RegFile.scala 97:16:@42301.4]
  assign rport_io_ins_497 = regs_497_io_out; // @[RegFile.scala 97:16:@42302.4]
  assign rport_io_ins_498 = regs_498_io_out; // @[RegFile.scala 97:16:@42303.4]
  assign rport_io_ins_499 = regs_499_io_out; // @[RegFile.scala 97:16:@42304.4]
  assign rport_io_ins_500 = regs_500_io_out; // @[RegFile.scala 97:16:@42305.4]
  assign rport_io_ins_501 = regs_501_io_out; // @[RegFile.scala 97:16:@42306.4]
  assign rport_io_ins_502 = regs_502_io_out; // @[RegFile.scala 97:16:@42307.4]
  assign rport_io_sel = io_raddr[8:0]; // @[RegFile.scala 106:18:@42308.4]
endmodule
module RetimeWrapper_518( // @[:@42330.2]
  input         clock, // @[:@42331.4]
  input         reset, // @[:@42332.4]
  input  [39:0] io_in, // @[:@42333.4]
  output [39:0] io_out // @[:@42333.4]
);
  wire [39:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@42335.4]
  wire [39:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@42335.4]
  wire [39:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@42335.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@42335.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@42335.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@42335.4]
  RetimeShiftRegister #(.WIDTH(40), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@42335.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@42348.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@42347.4]
  assign sr_init = 40'h0; // @[RetimeShiftRegister.scala 19:16:@42346.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@42345.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@42344.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@42342.4]
endmodule
module FringeFF_503( // @[:@42350.2]
  input         clock, // @[:@42351.4]
  input         reset, // @[:@42352.4]
  input  [39:0] io_in, // @[:@42353.4]
  output [39:0] io_out, // @[:@42353.4]
  input         io_enable // @[:@42353.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@42356.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@42356.4]
  wire [39:0] RetimeWrapper_io_in; // @[package.scala 93:22:@42356.4]
  wire [39:0] RetimeWrapper_io_out; // @[package.scala 93:22:@42356.4]
  wire [39:0] _T_18; // @[package.scala 96:25:@42361.4 package.scala 96:25:@42362.4]
  RetimeWrapper_518 RetimeWrapper ( // @[package.scala 93:22:@42356.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@42361.4 package.scala 96:25:@42362.4]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@42373.4]
  assign RetimeWrapper_clock = clock; // @[:@42357.4]
  assign RetimeWrapper_reset = reset; // @[:@42358.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _T_18; // @[package.scala 94:16:@42359.4]
endmodule
module FringeCounter( // @[:@42375.2]
  input   clock, // @[:@42376.4]
  input   reset, // @[:@42377.4]
  input   io_enable, // @[:@42378.4]
  output  io_done // @[:@42378.4]
);
  wire  reg$_clock; // @[FringeCounter.scala 24:19:@42380.4]
  wire  reg$_reset; // @[FringeCounter.scala 24:19:@42380.4]
  wire [39:0] reg$_io_in; // @[FringeCounter.scala 24:19:@42380.4]
  wire [39:0] reg$_io_out; // @[FringeCounter.scala 24:19:@42380.4]
  wire  reg$_io_enable; // @[FringeCounter.scala 24:19:@42380.4]
  wire [40:0] count; // @[Cat.scala 30:58:@42387.4]
  wire [41:0] _T_25; // @[FringeCounter.scala 31:22:@42388.4]
  wire [40:0] newval; // @[FringeCounter.scala 31:22:@42389.4]
  wire  isMax; // @[FringeCounter.scala 32:22:@42390.4]
  wire [40:0] next; // @[FringeCounter.scala 33:17:@42392.4]
  FringeFF_503 reg$ ( // @[FringeCounter.scala 24:19:@42380.4]
    .clock(reg$_clock),
    .reset(reg$_reset),
    .io_in(reg$_io_in),
    .io_out(reg$_io_out),
    .io_enable(reg$_io_enable)
  );
  assign count = {1'h0,reg$_io_out}; // @[Cat.scala 30:58:@42387.4]
  assign _T_25 = count + 41'h1; // @[FringeCounter.scala 31:22:@42388.4]
  assign newval = count + 41'h1; // @[FringeCounter.scala 31:22:@42389.4]
  assign isMax = newval >= 41'h2cb417800; // @[FringeCounter.scala 32:22:@42390.4]
  assign next = isMax ? count : newval; // @[FringeCounter.scala 33:17:@42392.4]
  assign io_done = io_enable & isMax; // @[FringeCounter.scala 43:11:@42403.4]
  assign reg$_clock = clock; // @[:@42381.4]
  assign reg$_reset = reset; // @[:@42382.4]
  assign reg$_io_in = next[39:0]; // @[FringeCounter.scala 35:15:@42394.6 FringeCounter.scala 37:15:@42397.6]
  assign reg$_io_enable = io_enable; // @[FringeCounter.scala 27:17:@42385.4]
endmodule
module FringeFF_504( // @[:@42437.2]
  input   clock, // @[:@42438.4]
  input   reset, // @[:@42439.4]
  input   io_in, // @[:@42440.4]
  input   io_reset, // @[:@42440.4]
  output  io_out, // @[:@42440.4]
  input   io_enable // @[:@42440.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@42443.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@42443.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@42443.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@42443.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@42443.4]
  wire  _T_18; // @[package.scala 96:25:@42448.4 package.scala 96:25:@42449.4]
  wire  _GEN_0; // @[FringeFF.scala 21:27:@42454.6]
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@42443.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@42448.4 package.scala 96:25:@42449.4]
  assign _GEN_0 = io_reset ? 1'h0 : _T_18; // @[FringeFF.scala 21:27:@42454.6]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@42460.4]
  assign RetimeWrapper_clock = clock; // @[:@42444.4]
  assign RetimeWrapper_reset = reset; // @[:@42445.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@42447.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _GEN_0; // @[package.scala 94:16:@42446.4]
endmodule
module Depulser( // @[:@42462.2]
  input   clock, // @[:@42463.4]
  input   reset, // @[:@42464.4]
  input   io_in, // @[:@42465.4]
  input   io_rst, // @[:@42465.4]
  output  io_out // @[:@42465.4]
);
  wire  r_clock; // @[Depulser.scala 14:17:@42467.4]
  wire  r_reset; // @[Depulser.scala 14:17:@42467.4]
  wire  r_io_in; // @[Depulser.scala 14:17:@42467.4]
  wire  r_io_reset; // @[Depulser.scala 14:17:@42467.4]
  wire  r_io_out; // @[Depulser.scala 14:17:@42467.4]
  wire  r_io_enable; // @[Depulser.scala 14:17:@42467.4]
  FringeFF_504 r ( // @[Depulser.scala 14:17:@42467.4]
    .clock(r_clock),
    .reset(r_reset),
    .io_in(r_io_in),
    .io_reset(r_io_reset),
    .io_out(r_io_out),
    .io_enable(r_io_enable)
  );
  assign io_out = r_io_out; // @[Depulser.scala 19:10:@42476.4]
  assign r_clock = clock; // @[:@42468.4]
  assign r_reset = reset; // @[:@42469.4]
  assign r_io_in = io_rst ? 1'h0 : io_in; // @[Depulser.scala 15:11:@42471.4]
  assign r_io_reset = io_rst; // @[Depulser.scala 18:14:@42475.4]
  assign r_io_enable = io_in | io_rst; // @[Depulser.scala 17:15:@42474.4]
endmodule
module Fringe( // @[:@42478.2]
  input         clock, // @[:@42479.4]
  input         reset, // @[:@42480.4]
  input  [31:0] io_raddr, // @[:@42481.4]
  input         io_wen, // @[:@42481.4]
  input  [31:0] io_waddr, // @[:@42481.4]
  input  [63:0] io_wdata, // @[:@42481.4]
  output [63:0] io_rdata, // @[:@42481.4]
  output        io_enable, // @[:@42481.4]
  input         io_done, // @[:@42481.4]
  output        io_reset, // @[:@42481.4]
  output [63:0] io_argIns_0, // @[:@42481.4]
  input         io_argOuts_0_valid, // @[:@42481.4]
  input  [63:0] io_argOuts_0_bits, // @[:@42481.4]
  input         io_heap_0_req_valid, // @[:@42481.4]
  input         io_heap_0_req_bits_allocDealloc, // @[:@42481.4]
  input  [63:0] io_heap_0_req_bits_sizeAddr, // @[:@42481.4]
  output        io_heap_0_resp_valid, // @[:@42481.4]
  output        io_heap_0_resp_bits_allocDealloc, // @[:@42481.4]
  output [63:0] io_heap_0_resp_bits_sizeAddr // @[:@42481.4]
);
  wire  heap_io_accel_0_req_valid; // @[Fringe.scala 107:20:@43510.4]
  wire  heap_io_accel_0_req_bits_allocDealloc; // @[Fringe.scala 107:20:@43510.4]
  wire [63:0] heap_io_accel_0_req_bits_sizeAddr; // @[Fringe.scala 107:20:@43510.4]
  wire  heap_io_accel_0_resp_valid; // @[Fringe.scala 107:20:@43510.4]
  wire  heap_io_accel_0_resp_bits_allocDealloc; // @[Fringe.scala 107:20:@43510.4]
  wire [63:0] heap_io_accel_0_resp_bits_sizeAddr; // @[Fringe.scala 107:20:@43510.4]
  wire  heap_io_host_0_req_valid; // @[Fringe.scala 107:20:@43510.4]
  wire  heap_io_host_0_req_bits_allocDealloc; // @[Fringe.scala 107:20:@43510.4]
  wire [63:0] heap_io_host_0_req_bits_sizeAddr; // @[Fringe.scala 107:20:@43510.4]
  wire  heap_io_host_0_resp_valid; // @[Fringe.scala 107:20:@43510.4]
  wire  heap_io_host_0_resp_bits_allocDealloc; // @[Fringe.scala 107:20:@43510.4]
  wire [63:0] heap_io_host_0_resp_bits_sizeAddr; // @[Fringe.scala 107:20:@43510.4]
  wire  regs_clock; // @[Fringe.scala 116:20:@43519.4]
  wire  regs_reset; // @[Fringe.scala 116:20:@43519.4]
  wire [31:0] regs_io_raddr; // @[Fringe.scala 116:20:@43519.4]
  wire  regs_io_wen; // @[Fringe.scala 116:20:@43519.4]
  wire [31:0] regs_io_waddr; // @[Fringe.scala 116:20:@43519.4]
  wire [63:0] regs_io_wdata; // @[Fringe.scala 116:20:@43519.4]
  wire [63:0] regs_io_rdata; // @[Fringe.scala 116:20:@43519.4]
  wire  regs_io_reset; // @[Fringe.scala 116:20:@43519.4]
  wire [63:0] regs_io_argIns_0; // @[Fringe.scala 116:20:@43519.4]
  wire [63:0] regs_io_argIns_1; // @[Fringe.scala 116:20:@43519.4]
  wire [63:0] regs_io_argIns_2; // @[Fringe.scala 116:20:@43519.4]
  wire  regs_io_argOuts_0_valid; // @[Fringe.scala 116:20:@43519.4]
  wire [63:0] regs_io_argOuts_0_bits; // @[Fringe.scala 116:20:@43519.4]
  wire  regs_io_argOuts_1_valid; // @[Fringe.scala 116:20:@43519.4]
  wire [63:0] regs_io_argOuts_1_bits; // @[Fringe.scala 116:20:@43519.4]
  wire  timeoutCtr_clock; // @[Fringe.scala 143:26:@45568.4]
  wire  timeoutCtr_reset; // @[Fringe.scala 143:26:@45568.4]
  wire  timeoutCtr_io_enable; // @[Fringe.scala 143:26:@45568.4]
  wire  timeoutCtr_io_done; // @[Fringe.scala 143:26:@45568.4]
  wire  depulser_clock; // @[Fringe.scala 153:24:@45586.4]
  wire  depulser_reset; // @[Fringe.scala 153:24:@45586.4]
  wire  depulser_io_in; // @[Fringe.scala 153:24:@45586.4]
  wire  depulser_io_rst; // @[Fringe.scala 153:24:@45586.4]
  wire  depulser_io_out; // @[Fringe.scala 153:24:@45586.4]
  wire [63:0] _T_826; // @[:@45545.4 :@45546.4]
  wire  curStatus_done; // @[Fringe.scala 133:45:@45547.4]
  wire  curStatus_timeout; // @[Fringe.scala 133:45:@45549.4]
  wire [2:0] curStatus_allocDealloc; // @[Fringe.scala 133:45:@45551.4]
  wire [58:0] curStatus_sizeAddr; // @[Fringe.scala 133:45:@45553.4]
  wire  _T_831; // @[Fringe.scala 134:28:@45555.4]
  wire  _T_835; // @[Fringe.scala 134:42:@45557.4]
  wire  _T_836; // @[Fringe.scala 135:27:@45559.4]
  wire [63:0] _T_846; // @[Fringe.scala 156:22:@45594.4]
  reg  _T_853; // @[package.scala 152:20:@45597.4]
  reg [31:0] _RAND_0;
  wire  _T_854; // @[package.scala 153:13:@45599.4]
  wire  _T_855; // @[package.scala 153:8:@45600.4]
  wire  _T_858; // @[Fringe.scala 160:55:@45604.4]
  wire  status_bits_done; // @[Fringe.scala 160:26:@45605.4]
  wire  _T_861; // @[Fringe.scala 161:58:@45608.4]
  wire  status_bits_timeout; // @[Fringe.scala 161:29:@45609.4]
  wire [1:0] _T_865; // @[Fringe.scala 162:57:@45611.4]
  wire [1:0] _T_867; // @[Fringe.scala 162:34:@45612.4]
  wire [63:0] _T_869; // @[Fringe.scala 163:30:@45614.4]
  wire [1:0] _T_870; // @[Fringe.scala 171:37:@45617.4]
  wire [58:0] status_bits_sizeAddr; // @[Fringe.scala 158:20:@45596.4 Fringe.scala 163:24:@45615.4]
  wire [2:0] status_bits_allocDealloc; // @[Fringe.scala 158:20:@45596.4 Fringe.scala 162:28:@45613.4]
  wire [61:0] _T_871; // @[Fringe.scala 171:37:@45618.4]
  wire  alloc; // @[Fringe.scala 202:38:@46903.4]
  wire  dealloc; // @[Fringe.scala 203:40:@46904.4]
  wire  _T_1375; // @[Fringe.scala 204:37:@46905.4]
  reg  _T_1378; // @[package.scala 152:20:@46906.4]
  reg [31:0] _RAND_1;
  wire  _T_1379; // @[package.scala 153:13:@46908.4]
  DRAMHeap heap ( // @[Fringe.scala 107:20:@43510.4]
    .io_accel_0_req_valid(heap_io_accel_0_req_valid),
    .io_accel_0_req_bits_allocDealloc(heap_io_accel_0_req_bits_allocDealloc),
    .io_accel_0_req_bits_sizeAddr(heap_io_accel_0_req_bits_sizeAddr),
    .io_accel_0_resp_valid(heap_io_accel_0_resp_valid),
    .io_accel_0_resp_bits_allocDealloc(heap_io_accel_0_resp_bits_allocDealloc),
    .io_accel_0_resp_bits_sizeAddr(heap_io_accel_0_resp_bits_sizeAddr),
    .io_host_0_req_valid(heap_io_host_0_req_valid),
    .io_host_0_req_bits_allocDealloc(heap_io_host_0_req_bits_allocDealloc),
    .io_host_0_req_bits_sizeAddr(heap_io_host_0_req_bits_sizeAddr),
    .io_host_0_resp_valid(heap_io_host_0_resp_valid),
    .io_host_0_resp_bits_allocDealloc(heap_io_host_0_resp_bits_allocDealloc),
    .io_host_0_resp_bits_sizeAddr(heap_io_host_0_resp_bits_sizeAddr)
  );
  RegFile regs ( // @[Fringe.scala 116:20:@43519.4]
    .clock(regs_clock),
    .reset(regs_reset),
    .io_raddr(regs_io_raddr),
    .io_wen(regs_io_wen),
    .io_waddr(regs_io_waddr),
    .io_wdata(regs_io_wdata),
    .io_rdata(regs_io_rdata),
    .io_reset(regs_io_reset),
    .io_argIns_0(regs_io_argIns_0),
    .io_argIns_1(regs_io_argIns_1),
    .io_argIns_2(regs_io_argIns_2),
    .io_argOuts_0_valid(regs_io_argOuts_0_valid),
    .io_argOuts_0_bits(regs_io_argOuts_0_bits),
    .io_argOuts_1_valid(regs_io_argOuts_1_valid),
    .io_argOuts_1_bits(regs_io_argOuts_1_bits)
  );
  FringeCounter timeoutCtr ( // @[Fringe.scala 143:26:@45568.4]
    .clock(timeoutCtr_clock),
    .reset(timeoutCtr_reset),
    .io_enable(timeoutCtr_io_enable),
    .io_done(timeoutCtr_io_done)
  );
  Depulser depulser ( // @[Fringe.scala 153:24:@45586.4]
    .clock(depulser_clock),
    .reset(depulser_reset),
    .io_in(depulser_io_in),
    .io_rst(depulser_io_rst),
    .io_out(depulser_io_out)
  );
  assign _T_826 = regs_io_argIns_1; // @[:@45545.4 :@45546.4]
  assign curStatus_done = _T_826[0]; // @[Fringe.scala 133:45:@45547.4]
  assign curStatus_timeout = _T_826[1]; // @[Fringe.scala 133:45:@45549.4]
  assign curStatus_allocDealloc = _T_826[4:2]; // @[Fringe.scala 133:45:@45551.4]
  assign curStatus_sizeAddr = _T_826[63:5]; // @[Fringe.scala 133:45:@45553.4]
  assign _T_831 = regs_io_argIns_0[0]; // @[Fringe.scala 134:28:@45555.4]
  assign _T_835 = curStatus_done == 1'h0; // @[Fringe.scala 134:42:@45557.4]
  assign _T_836 = regs_io_argIns_0[1]; // @[Fringe.scala 135:27:@45559.4]
  assign _T_846 = ~ regs_io_argIns_0; // @[Fringe.scala 156:22:@45594.4]
  assign _T_854 = _T_853 ^ heap_io_host_0_req_valid; // @[package.scala 153:13:@45599.4]
  assign _T_855 = heap_io_host_0_req_valid & _T_854; // @[package.scala 153:8:@45600.4]
  assign _T_858 = _T_831 & depulser_io_out; // @[Fringe.scala 160:55:@45604.4]
  assign status_bits_done = depulser_io_out ? _T_858 : curStatus_done; // @[Fringe.scala 160:26:@45605.4]
  assign _T_861 = _T_831 & timeoutCtr_io_done; // @[Fringe.scala 161:58:@45608.4]
  assign status_bits_timeout = depulser_io_out ? _T_861 : curStatus_timeout; // @[Fringe.scala 161:29:@45609.4]
  assign _T_865 = heap_io_host_0_req_bits_allocDealloc ? 2'h1 : 2'h2; // @[Fringe.scala 162:57:@45611.4]
  assign _T_867 = heap_io_host_0_req_valid ? _T_865 : 2'h0; // @[Fringe.scala 162:34:@45612.4]
  assign _T_869 = heap_io_host_0_req_valid ? heap_io_host_0_req_bits_sizeAddr : 64'h0; // @[Fringe.scala 163:30:@45614.4]
  assign _T_870 = {status_bits_timeout,status_bits_done}; // @[Fringe.scala 171:37:@45617.4]
  assign status_bits_sizeAddr = _T_869[58:0]; // @[Fringe.scala 158:20:@45596.4 Fringe.scala 163:24:@45615.4]
  assign status_bits_allocDealloc = {{1'd0}, _T_867}; // @[Fringe.scala 158:20:@45596.4 Fringe.scala 162:28:@45613.4]
  assign _T_871 = {status_bits_sizeAddr,status_bits_allocDealloc}; // @[Fringe.scala 171:37:@45618.4]
  assign alloc = curStatus_allocDealloc == 3'h3; // @[Fringe.scala 202:38:@46903.4]
  assign dealloc = curStatus_allocDealloc == 3'h4; // @[Fringe.scala 203:40:@46904.4]
  assign _T_1375 = alloc | dealloc; // @[Fringe.scala 204:37:@46905.4]
  assign _T_1379 = _T_1378 ^ _T_1375; // @[package.scala 153:13:@46908.4]
  assign io_rdata = regs_io_rdata; // @[Fringe.scala 125:14:@45543.4]
  assign io_enable = _T_831 & _T_835; // @[Fringe.scala 136:13:@45563.4]
  assign io_reset = _T_836 | reset; // @[Fringe.scala 137:12:@45564.4]
  assign io_argIns_0 = regs_io_argIns_2; // @[Fringe.scala 151:51:@45585.4]
  assign io_heap_0_resp_valid = heap_io_accel_0_resp_valid; // @[Fringe.scala 108:17:@43515.4]
  assign io_heap_0_resp_bits_allocDealloc = heap_io_accel_0_resp_bits_allocDealloc; // @[Fringe.scala 108:17:@43514.4]
  assign io_heap_0_resp_bits_sizeAddr = heap_io_accel_0_resp_bits_sizeAddr; // @[Fringe.scala 108:17:@43513.4]
  assign heap_io_accel_0_req_valid = io_heap_0_req_valid; // @[Fringe.scala 108:17:@43518.4]
  assign heap_io_accel_0_req_bits_allocDealloc = io_heap_0_req_bits_allocDealloc; // @[Fringe.scala 108:17:@43517.4]
  assign heap_io_accel_0_req_bits_sizeAddr = io_heap_0_req_bits_sizeAddr; // @[Fringe.scala 108:17:@43516.4]
  assign heap_io_host_0_resp_valid = _T_1375 & _T_1379; // @[Fringe.scala 204:22:@46910.4]
  assign heap_io_host_0_resp_bits_allocDealloc = curStatus_allocDealloc == 3'h3; // @[Fringe.scala 205:34:@46911.4]
  assign heap_io_host_0_resp_bits_sizeAddr = {{5'd0}, curStatus_sizeAddr}; // @[Fringe.scala 206:30:@46912.4]
  assign regs_clock = clock; // @[:@43520.4]
  assign regs_reset = reset; // @[:@43521.4 Fringe.scala 139:14:@45567.4]
  assign regs_io_raddr = io_raddr; // @[Fringe.scala 118:17:@45539.4]
  assign regs_io_wen = io_wen; // @[Fringe.scala 120:15:@45541.4]
  assign regs_io_waddr = io_waddr; // @[Fringe.scala 119:17:@45540.4]
  assign regs_io_wdata = io_wdata; // @[Fringe.scala 121:17:@45542.4]
  assign regs_io_reset = _T_836 | reset; // @[Fringe.scala 138:17:@45565.4]
  assign regs_io_argOuts_0_valid = depulser_io_out | _T_855; // @[Fringe.scala 170:23:@45616.4]
  assign regs_io_argOuts_0_bits = {_T_871,_T_870}; // @[Fringe.scala 171:22:@45620.4]
  assign regs_io_argOuts_1_valid = io_argOuts_0_valid; // @[Fringe.scala 176:23:@45623.4]
  assign regs_io_argOuts_1_bits = io_argOuts_0_bits; // @[Fringe.scala 175:22:@45622.4]
  assign timeoutCtr_clock = clock; // @[:@45569.4]
  assign timeoutCtr_reset = reset; // @[:@45570.4]
  assign timeoutCtr_io_enable = _T_831 & _T_835; // @[Fringe.scala 149:24:@45584.4]
  assign depulser_clock = clock; // @[:@45587.4]
  assign depulser_reset = reset; // @[:@45588.4]
  assign depulser_io_in = io_done | timeoutCtr_io_done; // @[Fringe.scala 155:18:@45593.4]
  assign depulser_io_rst = _T_846[0]; // @[Fringe.scala 156:19:@45595.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_853 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1378 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_853 <= 1'h0;
    end else begin
      _T_853 <= heap_io_host_0_req_valid;
    end
    if (reset) begin
      _T_1378 <= 1'h0;
    end else begin
      _T_1378 <= _T_1375;
    end
  end
endmodule
module AXI4LiteToRFBridgeKCU1500( // @[:@46927.2]
  input         clock, // @[:@46928.4]
  input         reset, // @[:@46929.4]
  input  [31:0] io_S_AXI_AWADDR, // @[:@46930.4]
  input  [2:0]  io_S_AXI_AWPROT, // @[:@46930.4]
  input         io_S_AXI_AWVALID, // @[:@46930.4]
  output        io_S_AXI_AWREADY, // @[:@46930.4]
  input  [31:0] io_S_AXI_ARADDR, // @[:@46930.4]
  input  [2:0]  io_S_AXI_ARPROT, // @[:@46930.4]
  input         io_S_AXI_ARVALID, // @[:@46930.4]
  output        io_S_AXI_ARREADY, // @[:@46930.4]
  input  [31:0] io_S_AXI_WDATA, // @[:@46930.4]
  input  [3:0]  io_S_AXI_WSTRB, // @[:@46930.4]
  input         io_S_AXI_WVALID, // @[:@46930.4]
  output        io_S_AXI_WREADY, // @[:@46930.4]
  output [31:0] io_S_AXI_RDATA, // @[:@46930.4]
  output [1:0]  io_S_AXI_RRESP, // @[:@46930.4]
  output        io_S_AXI_RVALID, // @[:@46930.4]
  input         io_S_AXI_RREADY, // @[:@46930.4]
  output [1:0]  io_S_AXI_BRESP, // @[:@46930.4]
  output        io_S_AXI_BVALID, // @[:@46930.4]
  input         io_S_AXI_BREADY, // @[:@46930.4]
  output [31:0] io_raddr, // @[:@46930.4]
  output        io_wen, // @[:@46930.4]
  output [31:0] io_waddr, // @[:@46930.4]
  output [31:0] io_wdata, // @[:@46930.4]
  input  [31:0] io_rdata // @[:@46930.4]
);
  wire [31:0] d_rf_rdata; // @[AXI4LiteToRFBridge.scala 109:17:@46932.4]
  wire [31:0] d_rf_wdata; // @[AXI4LiteToRFBridge.scala 109:17:@46932.4]
  wire [31:0] d_rf_waddr; // @[AXI4LiteToRFBridge.scala 109:17:@46932.4]
  wire  d_rf_wen; // @[AXI4LiteToRFBridge.scala 109:17:@46932.4]
  wire [31:0] d_rf_raddr; // @[AXI4LiteToRFBridge.scala 109:17:@46932.4]
  wire  d_S_AXI_ARESETN; // @[AXI4LiteToRFBridge.scala 109:17:@46932.4]
  wire  d_S_AXI_ACLK; // @[AXI4LiteToRFBridge.scala 109:17:@46932.4]
  wire [31:0] d_S_AXI_AWADDR; // @[AXI4LiteToRFBridge.scala 109:17:@46932.4]
  wire [2:0] d_S_AXI_AWPROT; // @[AXI4LiteToRFBridge.scala 109:17:@46932.4]
  wire  d_S_AXI_AWVALID; // @[AXI4LiteToRFBridge.scala 109:17:@46932.4]
  wire  d_S_AXI_AWREADY; // @[AXI4LiteToRFBridge.scala 109:17:@46932.4]
  wire [31:0] d_S_AXI_ARADDR; // @[AXI4LiteToRFBridge.scala 109:17:@46932.4]
  wire [2:0] d_S_AXI_ARPROT; // @[AXI4LiteToRFBridge.scala 109:17:@46932.4]
  wire  d_S_AXI_ARVALID; // @[AXI4LiteToRFBridge.scala 109:17:@46932.4]
  wire  d_S_AXI_ARREADY; // @[AXI4LiteToRFBridge.scala 109:17:@46932.4]
  wire [31:0] d_S_AXI_WDATA; // @[AXI4LiteToRFBridge.scala 109:17:@46932.4]
  wire [3:0] d_S_AXI_WSTRB; // @[AXI4LiteToRFBridge.scala 109:17:@46932.4]
  wire  d_S_AXI_WVALID; // @[AXI4LiteToRFBridge.scala 109:17:@46932.4]
  wire  d_S_AXI_WREADY; // @[AXI4LiteToRFBridge.scala 109:17:@46932.4]
  wire [31:0] d_S_AXI_RDATA; // @[AXI4LiteToRFBridge.scala 109:17:@46932.4]
  wire [1:0] d_S_AXI_RRESP; // @[AXI4LiteToRFBridge.scala 109:17:@46932.4]
  wire  d_S_AXI_RVALID; // @[AXI4LiteToRFBridge.scala 109:17:@46932.4]
  wire  d_S_AXI_RREADY; // @[AXI4LiteToRFBridge.scala 109:17:@46932.4]
  wire [1:0] d_S_AXI_BRESP; // @[AXI4LiteToRFBridge.scala 109:17:@46932.4]
  wire  d_S_AXI_BVALID; // @[AXI4LiteToRFBridge.scala 109:17:@46932.4]
  wire  d_S_AXI_BREADY; // @[AXI4LiteToRFBridge.scala 109:17:@46932.4]
  AXI4LiteToRFBridgeVerilog d ( // @[AXI4LiteToRFBridge.scala 109:17:@46932.4]
    .rf_rdata(d_rf_rdata),
    .rf_wdata(d_rf_wdata),
    .rf_waddr(d_rf_waddr),
    .rf_wen(d_rf_wen),
    .rf_raddr(d_rf_raddr),
    .S_AXI_ARESETN(d_S_AXI_ARESETN),
    .S_AXI_ACLK(d_S_AXI_ACLK),
    .S_AXI_AWADDR(d_S_AXI_AWADDR),
    .S_AXI_AWPROT(d_S_AXI_AWPROT),
    .S_AXI_AWVALID(d_S_AXI_AWVALID),
    .S_AXI_AWREADY(d_S_AXI_AWREADY),
    .S_AXI_ARADDR(d_S_AXI_ARADDR),
    .S_AXI_ARPROT(d_S_AXI_ARPROT),
    .S_AXI_ARVALID(d_S_AXI_ARVALID),
    .S_AXI_ARREADY(d_S_AXI_ARREADY),
    .S_AXI_WDATA(d_S_AXI_WDATA),
    .S_AXI_WSTRB(d_S_AXI_WSTRB),
    .S_AXI_WVALID(d_S_AXI_WVALID),
    .S_AXI_WREADY(d_S_AXI_WREADY),
    .S_AXI_RDATA(d_S_AXI_RDATA),
    .S_AXI_RRESP(d_S_AXI_RRESP),
    .S_AXI_RVALID(d_S_AXI_RVALID),
    .S_AXI_RREADY(d_S_AXI_RREADY),
    .S_AXI_BRESP(d_S_AXI_BRESP),
    .S_AXI_BVALID(d_S_AXI_BVALID),
    .S_AXI_BREADY(d_S_AXI_BREADY)
  );
  assign io_S_AXI_AWREADY = d_S_AXI_AWREADY; // @[AXI4LiteToRFBridge.scala 111:14:@46956.4]
  assign io_S_AXI_ARREADY = d_S_AXI_ARREADY; // @[AXI4LiteToRFBridge.scala 111:14:@46952.4]
  assign io_S_AXI_WREADY = d_S_AXI_WREADY; // @[AXI4LiteToRFBridge.scala 111:14:@46948.4]
  assign io_S_AXI_RDATA = d_S_AXI_RDATA; // @[AXI4LiteToRFBridge.scala 111:14:@46947.4]
  assign io_S_AXI_RRESP = d_S_AXI_RRESP; // @[AXI4LiteToRFBridge.scala 111:14:@46946.4]
  assign io_S_AXI_RVALID = d_S_AXI_RVALID; // @[AXI4LiteToRFBridge.scala 111:14:@46945.4]
  assign io_S_AXI_BRESP = d_S_AXI_BRESP; // @[AXI4LiteToRFBridge.scala 111:14:@46943.4]
  assign io_S_AXI_BVALID = d_S_AXI_BVALID; // @[AXI4LiteToRFBridge.scala 111:14:@46942.4]
  assign io_raddr = d_rf_raddr; // @[AXI4LiteToRFBridge.scala 115:12:@46964.4]
  assign io_wen = d_rf_wen; // @[AXI4LiteToRFBridge.scala 118:12:@46967.4]
  assign io_waddr = d_rf_waddr; // @[AXI4LiteToRFBridge.scala 116:12:@46965.4]
  assign io_wdata = d_rf_wdata; // @[AXI4LiteToRFBridge.scala 117:12:@46966.4]
  assign d_rf_rdata = io_rdata; // @[AXI4LiteToRFBridge.scala 119:17:@46968.4]
  assign d_S_AXI_ARESETN = ~ reset; // @[AXI4LiteToRFBridge.scala 113:22:@46963.4]
  assign d_S_AXI_ACLK = clock; // @[AXI4LiteToRFBridge.scala 112:19:@46960.4]
  assign d_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[AXI4LiteToRFBridge.scala 111:14:@46959.4]
  assign d_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[AXI4LiteToRFBridge.scala 111:14:@46958.4]
  assign d_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[AXI4LiteToRFBridge.scala 111:14:@46957.4]
  assign d_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[AXI4LiteToRFBridge.scala 111:14:@46955.4]
  assign d_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[AXI4LiteToRFBridge.scala 111:14:@46954.4]
  assign d_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[AXI4LiteToRFBridge.scala 111:14:@46953.4]
  assign d_S_AXI_WDATA = io_S_AXI_WDATA; // @[AXI4LiteToRFBridge.scala 111:14:@46951.4]
  assign d_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[AXI4LiteToRFBridge.scala 111:14:@46950.4]
  assign d_S_AXI_WVALID = io_S_AXI_WVALID; // @[AXI4LiteToRFBridge.scala 111:14:@46949.4]
  assign d_S_AXI_RREADY = io_S_AXI_RREADY; // @[AXI4LiteToRFBridge.scala 111:14:@46944.4]
  assign d_S_AXI_BREADY = io_S_AXI_BREADY; // @[AXI4LiteToRFBridge.scala 111:14:@46941.4]
endmodule
module MAGToAXI4Bridge( // @[:@46970.2]
  output [7:0] io_M_AXI_AWLEN, // @[:@46973.4]
  output [7:0] io_M_AXI_ARLEN // @[:@46973.4]
);
  wire [32:0] _T_218; // @[MAGToAXI4Bridge.scala 27:29:@47130.4]
  wire [32:0] _T_219; // @[MAGToAXI4Bridge.scala 27:29:@47131.4]
  wire [31:0] _T_220; // @[MAGToAXI4Bridge.scala 27:29:@47132.4]
  assign _T_218 = 32'h0 - 32'h1; // @[MAGToAXI4Bridge.scala 27:29:@47130.4]
  assign _T_219 = $unsigned(_T_218); // @[MAGToAXI4Bridge.scala 27:29:@47131.4]
  assign _T_220 = _T_219[31:0]; // @[MAGToAXI4Bridge.scala 27:29:@47132.4]
  assign io_M_AXI_AWLEN = _T_220[7:0]; // @[MAGToAXI4Bridge.scala 41:21:@47150.4]
  assign io_M_AXI_ARLEN = _T_220[7:0]; // @[MAGToAXI4Bridge.scala 27:21:@47133.4]
endmodule
module FringeZynq( // @[:@47298.2]
  input         clock, // @[:@47299.4]
  input         reset, // @[:@47300.4]
  input  [31:0] io_S_AXI_AWADDR, // @[:@47301.4]
  input  [2:0]  io_S_AXI_AWPROT, // @[:@47301.4]
  input         io_S_AXI_AWVALID, // @[:@47301.4]
  output        io_S_AXI_AWREADY, // @[:@47301.4]
  input  [31:0] io_S_AXI_ARADDR, // @[:@47301.4]
  input  [2:0]  io_S_AXI_ARPROT, // @[:@47301.4]
  input         io_S_AXI_ARVALID, // @[:@47301.4]
  output        io_S_AXI_ARREADY, // @[:@47301.4]
  input  [31:0] io_S_AXI_WDATA, // @[:@47301.4]
  input  [3:0]  io_S_AXI_WSTRB, // @[:@47301.4]
  input         io_S_AXI_WVALID, // @[:@47301.4]
  output        io_S_AXI_WREADY, // @[:@47301.4]
  output [31:0] io_S_AXI_RDATA, // @[:@47301.4]
  output [1:0]  io_S_AXI_RRESP, // @[:@47301.4]
  output        io_S_AXI_RVALID, // @[:@47301.4]
  input         io_S_AXI_RREADY, // @[:@47301.4]
  output [1:0]  io_S_AXI_BRESP, // @[:@47301.4]
  output        io_S_AXI_BVALID, // @[:@47301.4]
  input         io_S_AXI_BREADY, // @[:@47301.4]
  output [7:0]  io_M_AXI_0_AWLEN, // @[:@47301.4]
  output [7:0]  io_M_AXI_0_ARLEN, // @[:@47301.4]
  output        io_enable, // @[:@47301.4]
  input         io_done, // @[:@47301.4]
  output        io_reset, // @[:@47301.4]
  output [63:0] io_argIns_0, // @[:@47301.4]
  input         io_argOuts_0_valid, // @[:@47301.4]
  input  [63:0] io_argOuts_0_bits, // @[:@47301.4]
  input         io_heap_0_req_valid, // @[:@47301.4]
  input         io_heap_0_req_bits_allocDealloc, // @[:@47301.4]
  input  [63:0] io_heap_0_req_bits_sizeAddr, // @[:@47301.4]
  output        io_heap_0_resp_valid, // @[:@47301.4]
  output        io_heap_0_resp_bits_allocDealloc, // @[:@47301.4]
  output [63:0] io_heap_0_resp_bits_sizeAddr // @[:@47301.4]
);
  wire  fringeCommon_clock; // @[FringeZynq.scala 68:28:@47663.4]
  wire  fringeCommon_reset; // @[FringeZynq.scala 68:28:@47663.4]
  wire [31:0] fringeCommon_io_raddr; // @[FringeZynq.scala 68:28:@47663.4]
  wire  fringeCommon_io_wen; // @[FringeZynq.scala 68:28:@47663.4]
  wire [31:0] fringeCommon_io_waddr; // @[FringeZynq.scala 68:28:@47663.4]
  wire [63:0] fringeCommon_io_wdata; // @[FringeZynq.scala 68:28:@47663.4]
  wire [63:0] fringeCommon_io_rdata; // @[FringeZynq.scala 68:28:@47663.4]
  wire  fringeCommon_io_enable; // @[FringeZynq.scala 68:28:@47663.4]
  wire  fringeCommon_io_done; // @[FringeZynq.scala 68:28:@47663.4]
  wire  fringeCommon_io_reset; // @[FringeZynq.scala 68:28:@47663.4]
  wire [63:0] fringeCommon_io_argIns_0; // @[FringeZynq.scala 68:28:@47663.4]
  wire  fringeCommon_io_argOuts_0_valid; // @[FringeZynq.scala 68:28:@47663.4]
  wire [63:0] fringeCommon_io_argOuts_0_bits; // @[FringeZynq.scala 68:28:@47663.4]
  wire  fringeCommon_io_heap_0_req_valid; // @[FringeZynq.scala 68:28:@47663.4]
  wire  fringeCommon_io_heap_0_req_bits_allocDealloc; // @[FringeZynq.scala 68:28:@47663.4]
  wire [63:0] fringeCommon_io_heap_0_req_bits_sizeAddr; // @[FringeZynq.scala 68:28:@47663.4]
  wire  fringeCommon_io_heap_0_resp_valid; // @[FringeZynq.scala 68:28:@47663.4]
  wire  fringeCommon_io_heap_0_resp_bits_allocDealloc; // @[FringeZynq.scala 68:28:@47663.4]
  wire [63:0] fringeCommon_io_heap_0_resp_bits_sizeAddr; // @[FringeZynq.scala 68:28:@47663.4]
  wire  AXI4LiteToRFBridgeKCU1500_clock; // @[FringeZynq.scala 78:31:@48247.4]
  wire  AXI4LiteToRFBridgeKCU1500_reset; // @[FringeZynq.scala 78:31:@48247.4]
  wire [31:0] AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWADDR; // @[FringeZynq.scala 78:31:@48247.4]
  wire [2:0] AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWPROT; // @[FringeZynq.scala 78:31:@48247.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWVALID; // @[FringeZynq.scala 78:31:@48247.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWREADY; // @[FringeZynq.scala 78:31:@48247.4]
  wire [31:0] AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARADDR; // @[FringeZynq.scala 78:31:@48247.4]
  wire [2:0] AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARPROT; // @[FringeZynq.scala 78:31:@48247.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARVALID; // @[FringeZynq.scala 78:31:@48247.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARREADY; // @[FringeZynq.scala 78:31:@48247.4]
  wire [31:0] AXI4LiteToRFBridgeKCU1500_io_S_AXI_WDATA; // @[FringeZynq.scala 78:31:@48247.4]
  wire [3:0] AXI4LiteToRFBridgeKCU1500_io_S_AXI_WSTRB; // @[FringeZynq.scala 78:31:@48247.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_WVALID; // @[FringeZynq.scala 78:31:@48247.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_WREADY; // @[FringeZynq.scala 78:31:@48247.4]
  wire [31:0] AXI4LiteToRFBridgeKCU1500_io_S_AXI_RDATA; // @[FringeZynq.scala 78:31:@48247.4]
  wire [1:0] AXI4LiteToRFBridgeKCU1500_io_S_AXI_RRESP; // @[FringeZynq.scala 78:31:@48247.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_RVALID; // @[FringeZynq.scala 78:31:@48247.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_RREADY; // @[FringeZynq.scala 78:31:@48247.4]
  wire [1:0] AXI4LiteToRFBridgeKCU1500_io_S_AXI_BRESP; // @[FringeZynq.scala 78:31:@48247.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_BVALID; // @[FringeZynq.scala 78:31:@48247.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_BREADY; // @[FringeZynq.scala 78:31:@48247.4]
  wire [31:0] AXI4LiteToRFBridgeKCU1500_io_raddr; // @[FringeZynq.scala 78:31:@48247.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_wen; // @[FringeZynq.scala 78:31:@48247.4]
  wire [31:0] AXI4LiteToRFBridgeKCU1500_io_waddr; // @[FringeZynq.scala 78:31:@48247.4]
  wire [31:0] AXI4LiteToRFBridgeKCU1500_io_wdata; // @[FringeZynq.scala 78:31:@48247.4]
  wire [31:0] AXI4LiteToRFBridgeKCU1500_io_rdata; // @[FringeZynq.scala 78:31:@48247.4]
  wire [7:0] MAGToAXI4Bridge_io_M_AXI_AWLEN; // @[FringeZynq.scala 130:27:@48413.4]
  wire [7:0] MAGToAXI4Bridge_io_M_AXI_ARLEN; // @[FringeZynq.scala 130:27:@48413.4]
  Fringe fringeCommon ( // @[FringeZynq.scala 68:28:@47663.4]
    .clock(fringeCommon_clock),
    .reset(fringeCommon_reset),
    .io_raddr(fringeCommon_io_raddr),
    .io_wen(fringeCommon_io_wen),
    .io_waddr(fringeCommon_io_waddr),
    .io_wdata(fringeCommon_io_wdata),
    .io_rdata(fringeCommon_io_rdata),
    .io_enable(fringeCommon_io_enable),
    .io_done(fringeCommon_io_done),
    .io_reset(fringeCommon_io_reset),
    .io_argIns_0(fringeCommon_io_argIns_0),
    .io_argOuts_0_valid(fringeCommon_io_argOuts_0_valid),
    .io_argOuts_0_bits(fringeCommon_io_argOuts_0_bits),
    .io_heap_0_req_valid(fringeCommon_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(fringeCommon_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(fringeCommon_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(fringeCommon_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(fringeCommon_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(fringeCommon_io_heap_0_resp_bits_sizeAddr)
  );
  AXI4LiteToRFBridgeKCU1500 AXI4LiteToRFBridgeKCU1500 ( // @[FringeZynq.scala 78:31:@48247.4]
    .clock(AXI4LiteToRFBridgeKCU1500_clock),
    .reset(AXI4LiteToRFBridgeKCU1500_reset),
    .io_S_AXI_AWADDR(AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWADDR),
    .io_S_AXI_AWPROT(AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWPROT),
    .io_S_AXI_AWVALID(AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWVALID),
    .io_S_AXI_AWREADY(AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWREADY),
    .io_S_AXI_ARADDR(AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARADDR),
    .io_S_AXI_ARPROT(AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARPROT),
    .io_S_AXI_ARVALID(AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARVALID),
    .io_S_AXI_ARREADY(AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARREADY),
    .io_S_AXI_WDATA(AXI4LiteToRFBridgeKCU1500_io_S_AXI_WDATA),
    .io_S_AXI_WSTRB(AXI4LiteToRFBridgeKCU1500_io_S_AXI_WSTRB),
    .io_S_AXI_WVALID(AXI4LiteToRFBridgeKCU1500_io_S_AXI_WVALID),
    .io_S_AXI_WREADY(AXI4LiteToRFBridgeKCU1500_io_S_AXI_WREADY),
    .io_S_AXI_RDATA(AXI4LiteToRFBridgeKCU1500_io_S_AXI_RDATA),
    .io_S_AXI_RRESP(AXI4LiteToRFBridgeKCU1500_io_S_AXI_RRESP),
    .io_S_AXI_RVALID(AXI4LiteToRFBridgeKCU1500_io_S_AXI_RVALID),
    .io_S_AXI_RREADY(AXI4LiteToRFBridgeKCU1500_io_S_AXI_RREADY),
    .io_S_AXI_BRESP(AXI4LiteToRFBridgeKCU1500_io_S_AXI_BRESP),
    .io_S_AXI_BVALID(AXI4LiteToRFBridgeKCU1500_io_S_AXI_BVALID),
    .io_S_AXI_BREADY(AXI4LiteToRFBridgeKCU1500_io_S_AXI_BREADY),
    .io_raddr(AXI4LiteToRFBridgeKCU1500_io_raddr),
    .io_wen(AXI4LiteToRFBridgeKCU1500_io_wen),
    .io_waddr(AXI4LiteToRFBridgeKCU1500_io_waddr),
    .io_wdata(AXI4LiteToRFBridgeKCU1500_io_wdata),
    .io_rdata(AXI4LiteToRFBridgeKCU1500_io_rdata)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge ( // @[FringeZynq.scala 130:27:@48413.4]
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_io_M_AXI_AWLEN),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_io_M_AXI_ARLEN)
  );
  assign io_S_AXI_AWREADY = AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWREADY; // @[FringeZynq.scala 79:28:@48265.4]
  assign io_S_AXI_ARREADY = AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARREADY; // @[FringeZynq.scala 79:28:@48261.4]
  assign io_S_AXI_WREADY = AXI4LiteToRFBridgeKCU1500_io_S_AXI_WREADY; // @[FringeZynq.scala 79:28:@48257.4]
  assign io_S_AXI_RDATA = AXI4LiteToRFBridgeKCU1500_io_S_AXI_RDATA; // @[FringeZynq.scala 79:28:@48256.4]
  assign io_S_AXI_RRESP = AXI4LiteToRFBridgeKCU1500_io_S_AXI_RRESP; // @[FringeZynq.scala 79:28:@48255.4]
  assign io_S_AXI_RVALID = AXI4LiteToRFBridgeKCU1500_io_S_AXI_RVALID; // @[FringeZynq.scala 79:28:@48254.4]
  assign io_S_AXI_BRESP = AXI4LiteToRFBridgeKCU1500_io_S_AXI_BRESP; // @[FringeZynq.scala 79:28:@48252.4]
  assign io_S_AXI_BVALID = AXI4LiteToRFBridgeKCU1500_io_S_AXI_BVALID; // @[FringeZynq.scala 79:28:@48251.4]
  assign io_M_AXI_0_AWLEN = MAGToAXI4Bridge_io_M_AXI_AWLEN; // @[FringeZynq.scala 132:10:@48565.4]
  assign io_M_AXI_0_ARLEN = MAGToAXI4Bridge_io_M_AXI_ARLEN; // @[FringeZynq.scala 132:10:@48553.4]
  assign io_enable = fringeCommon_io_enable; // @[FringeZynq.scala 114:13:@48277.4]
  assign io_reset = fringeCommon_io_reset; // @[FringeZynq.scala 118:12:@48281.4]
  assign io_argIns_0 = fringeCommon_io_argIns_0; // @[FringeZynq.scala 120:13:@48282.4]
  assign io_heap_0_resp_valid = fringeCommon_io_heap_0_resp_valid; // @[FringeZynq.scala 126:11:@48409.4]
  assign io_heap_0_resp_bits_allocDealloc = fringeCommon_io_heap_0_resp_bits_allocDealloc; // @[FringeZynq.scala 126:11:@48408.4]
  assign io_heap_0_resp_bits_sizeAddr = fringeCommon_io_heap_0_resp_bits_sizeAddr; // @[FringeZynq.scala 126:11:@48407.4]
  assign fringeCommon_clock = clock; // @[:@47664.4]
  assign fringeCommon_reset = reset; // @[:@47665.4 FringeZynq.scala 81:24:@48270.4 FringeZynq.scala 116:22:@48280.4]
  assign fringeCommon_io_raddr = AXI4LiteToRFBridgeKCU1500_io_raddr; // @[FringeZynq.scala 82:27:@48271.4]
  assign fringeCommon_io_wen = AXI4LiteToRFBridgeKCU1500_io_wen; // @[FringeZynq.scala 83:27:@48272.4]
  assign fringeCommon_io_waddr = AXI4LiteToRFBridgeKCU1500_io_waddr; // @[FringeZynq.scala 84:27:@48273.4]
  assign fringeCommon_io_wdata = {{32'd0}, AXI4LiteToRFBridgeKCU1500_io_wdata}; // @[FringeZynq.scala 85:27:@48274.4]
  assign fringeCommon_io_done = io_done; // @[FringeZynq.scala 115:24:@48278.4]
  assign fringeCommon_io_argOuts_0_valid = io_argOuts_0_valid; // @[FringeZynq.scala 121:27:@48284.4]
  assign fringeCommon_io_argOuts_0_bits = io_argOuts_0_bits; // @[FringeZynq.scala 121:27:@48283.4]
  assign fringeCommon_io_heap_0_req_valid = io_heap_0_req_valid; // @[FringeZynq.scala 126:11:@48412.4]
  assign fringeCommon_io_heap_0_req_bits_allocDealloc = io_heap_0_req_bits_allocDealloc; // @[FringeZynq.scala 126:11:@48411.4]
  assign fringeCommon_io_heap_0_req_bits_sizeAddr = io_heap_0_req_bits_sizeAddr; // @[FringeZynq.scala 126:11:@48410.4]
  assign AXI4LiteToRFBridgeKCU1500_clock = clock; // @[:@48248.4]
  assign AXI4LiteToRFBridgeKCU1500_reset = reset; // @[:@48249.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[FringeZynq.scala 79:28:@48268.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[FringeZynq.scala 79:28:@48267.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[FringeZynq.scala 79:28:@48266.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[FringeZynq.scala 79:28:@48264.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[FringeZynq.scala 79:28:@48263.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[FringeZynq.scala 79:28:@48262.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_WDATA = io_S_AXI_WDATA; // @[FringeZynq.scala 79:28:@48260.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[FringeZynq.scala 79:28:@48259.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_WVALID = io_S_AXI_WVALID; // @[FringeZynq.scala 79:28:@48258.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_RREADY = io_S_AXI_RREADY; // @[FringeZynq.scala 79:28:@48253.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_BREADY = io_S_AXI_BREADY; // @[FringeZynq.scala 79:28:@48250.4]
  assign AXI4LiteToRFBridgeKCU1500_io_rdata = fringeCommon_io_rdata[31:0]; // @[FringeZynq.scala 86:28:@48275.4]
endmodule
module Top( // @[:@48570.2]
  input          clock, // @[:@48571.4]
  input          reset, // @[:@48572.4]
  input          io_raddr, // @[:@48573.4]
  input          io_wen, // @[:@48573.4]
  input          io_waddr, // @[:@48573.4]
  input          io_wdata, // @[:@48573.4]
  output         io_rdata, // @[:@48573.4]
  input  [31:0]  io_S_AXI_AWADDR, // @[:@48573.4]
  input  [2:0]   io_S_AXI_AWPROT, // @[:@48573.4]
  input          io_S_AXI_AWVALID, // @[:@48573.4]
  output         io_S_AXI_AWREADY, // @[:@48573.4]
  input  [31:0]  io_S_AXI_ARADDR, // @[:@48573.4]
  input  [2:0]   io_S_AXI_ARPROT, // @[:@48573.4]
  input          io_S_AXI_ARVALID, // @[:@48573.4]
  output         io_S_AXI_ARREADY, // @[:@48573.4]
  input  [31:0]  io_S_AXI_WDATA, // @[:@48573.4]
  input  [3:0]   io_S_AXI_WSTRB, // @[:@48573.4]
  input          io_S_AXI_WVALID, // @[:@48573.4]
  output         io_S_AXI_WREADY, // @[:@48573.4]
  output [31:0]  io_S_AXI_RDATA, // @[:@48573.4]
  output [1:0]   io_S_AXI_RRESP, // @[:@48573.4]
  output         io_S_AXI_RVALID, // @[:@48573.4]
  input          io_S_AXI_RREADY, // @[:@48573.4]
  output [1:0]   io_S_AXI_BRESP, // @[:@48573.4]
  output         io_S_AXI_BVALID, // @[:@48573.4]
  input          io_S_AXI_BREADY, // @[:@48573.4]
  output [3:0]   io_M_AXI_0_AWID, // @[:@48573.4]
  output [3:0]   io_M_AXI_0_AWUSER, // @[:@48573.4]
  output [31:0]  io_M_AXI_0_AWADDR, // @[:@48573.4]
  output [7:0]   io_M_AXI_0_AWLEN, // @[:@48573.4]
  output [2:0]   io_M_AXI_0_AWSIZE, // @[:@48573.4]
  output [1:0]   io_M_AXI_0_AWBURST, // @[:@48573.4]
  output         io_M_AXI_0_AWLOCK, // @[:@48573.4]
  output [3:0]   io_M_AXI_0_AWCACHE, // @[:@48573.4]
  output [2:0]   io_M_AXI_0_AWPROT, // @[:@48573.4]
  output [3:0]   io_M_AXI_0_AWQOS, // @[:@48573.4]
  output         io_M_AXI_0_AWVALID, // @[:@48573.4]
  input          io_M_AXI_0_AWREADY, // @[:@48573.4]
  output [3:0]   io_M_AXI_0_ARID, // @[:@48573.4]
  output [3:0]   io_M_AXI_0_ARUSER, // @[:@48573.4]
  output [31:0]  io_M_AXI_0_ARADDR, // @[:@48573.4]
  output [7:0]   io_M_AXI_0_ARLEN, // @[:@48573.4]
  output [2:0]   io_M_AXI_0_ARSIZE, // @[:@48573.4]
  output [1:0]   io_M_AXI_0_ARBURST, // @[:@48573.4]
  output         io_M_AXI_0_ARLOCK, // @[:@48573.4]
  output [3:0]   io_M_AXI_0_ARCACHE, // @[:@48573.4]
  output [2:0]   io_M_AXI_0_ARPROT, // @[:@48573.4]
  output [3:0]   io_M_AXI_0_ARQOS, // @[:@48573.4]
  output         io_M_AXI_0_ARVALID, // @[:@48573.4]
  input          io_M_AXI_0_ARREADY, // @[:@48573.4]
  output [511:0] io_M_AXI_0_WDATA, // @[:@48573.4]
  output [63:0]  io_M_AXI_0_WSTRB, // @[:@48573.4]
  output         io_M_AXI_0_WLAST, // @[:@48573.4]
  output         io_M_AXI_0_WVALID, // @[:@48573.4]
  input          io_M_AXI_0_WREADY, // @[:@48573.4]
  input  [3:0]   io_M_AXI_0_RID, // @[:@48573.4]
  input  [31:0]  io_M_AXI_0_RUSER, // @[:@48573.4]
  input  [511:0] io_M_AXI_0_RDATA, // @[:@48573.4]
  input  [1:0]   io_M_AXI_0_RRESP, // @[:@48573.4]
  input          io_M_AXI_0_RLAST, // @[:@48573.4]
  input          io_M_AXI_0_RVALID, // @[:@48573.4]
  output         io_M_AXI_0_RREADY, // @[:@48573.4]
  input  [3:0]   io_M_AXI_0_BID, // @[:@48573.4]
  input  [3:0]   io_M_AXI_0_BUSER, // @[:@48573.4]
  input  [1:0]   io_M_AXI_0_BRESP, // @[:@48573.4]
  input          io_M_AXI_0_BVALID, // @[:@48573.4]
  output         io_M_AXI_0_BREADY // @[:@48573.4]
);
  wire  accel_clock; // @[Instantiator.scala 54:38:@48575.4]
  wire  accel_reset; // @[Instantiator.scala 54:38:@48575.4]
  wire  accel_io_enable; // @[Instantiator.scala 54:38:@48575.4]
  wire  accel_io_done; // @[Instantiator.scala 54:38:@48575.4]
  wire  accel_io_reset; // @[Instantiator.scala 54:38:@48575.4]
  wire  accel_io_memStreams_loads_0_cmd_ready; // @[Instantiator.scala 54:38:@48575.4]
  wire  accel_io_memStreams_loads_0_cmd_valid; // @[Instantiator.scala 54:38:@48575.4]
  wire [63:0] accel_io_memStreams_loads_0_cmd_bits_addr; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_loads_0_cmd_bits_size; // @[Instantiator.scala 54:38:@48575.4]
  wire  accel_io_memStreams_loads_0_data_ready; // @[Instantiator.scala 54:38:@48575.4]
  wire  accel_io_memStreams_loads_0_data_valid; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_0; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_1; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_2; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_3; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_4; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_5; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_6; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_7; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_8; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_9; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_10; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_11; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_12; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_13; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_14; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_15; // @[Instantiator.scala 54:38:@48575.4]
  wire  accel_io_memStreams_stores_0_cmd_ready; // @[Instantiator.scala 54:38:@48575.4]
  wire  accel_io_memStreams_stores_0_cmd_valid; // @[Instantiator.scala 54:38:@48575.4]
  wire [63:0] accel_io_memStreams_stores_0_cmd_bits_addr; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_stores_0_cmd_bits_size; // @[Instantiator.scala 54:38:@48575.4]
  wire  accel_io_memStreams_stores_0_data_ready; // @[Instantiator.scala 54:38:@48575.4]
  wire  accel_io_memStreams_stores_0_data_valid; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_0; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_1; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_2; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_3; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_4; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_5; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_6; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_7; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_8; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_9; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_10; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_11; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_12; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_13; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_14; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_15; // @[Instantiator.scala 54:38:@48575.4]
  wire [15:0] accel_io_memStreams_stores_0_data_bits_wstrb; // @[Instantiator.scala 54:38:@48575.4]
  wire  accel_io_memStreams_stores_0_wresp_ready; // @[Instantiator.scala 54:38:@48575.4]
  wire  accel_io_memStreams_stores_0_wresp_valid; // @[Instantiator.scala 54:38:@48575.4]
  wire  accel_io_memStreams_stores_0_wresp_bits; // @[Instantiator.scala 54:38:@48575.4]
  wire  accel_io_memStreams_gathers_0_cmd_ready; // @[Instantiator.scala 54:38:@48575.4]
  wire  accel_io_memStreams_gathers_0_cmd_valid; // @[Instantiator.scala 54:38:@48575.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_0; // @[Instantiator.scala 54:38:@48575.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_1; // @[Instantiator.scala 54:38:@48575.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_2; // @[Instantiator.scala 54:38:@48575.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_3; // @[Instantiator.scala 54:38:@48575.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_4; // @[Instantiator.scala 54:38:@48575.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_5; // @[Instantiator.scala 54:38:@48575.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_6; // @[Instantiator.scala 54:38:@48575.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_7; // @[Instantiator.scala 54:38:@48575.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_8; // @[Instantiator.scala 54:38:@48575.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_9; // @[Instantiator.scala 54:38:@48575.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_10; // @[Instantiator.scala 54:38:@48575.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_11; // @[Instantiator.scala 54:38:@48575.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_12; // @[Instantiator.scala 54:38:@48575.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_13; // @[Instantiator.scala 54:38:@48575.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_14; // @[Instantiator.scala 54:38:@48575.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_15; // @[Instantiator.scala 54:38:@48575.4]
  wire  accel_io_memStreams_gathers_0_data_ready; // @[Instantiator.scala 54:38:@48575.4]
  wire  accel_io_memStreams_gathers_0_data_valid; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_0; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_1; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_2; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_3; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_4; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_5; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_6; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_7; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_8; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_9; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_10; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_11; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_12; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_13; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_14; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_15; // @[Instantiator.scala 54:38:@48575.4]
  wire  accel_io_memStreams_scatters_0_cmd_ready; // @[Instantiator.scala 54:38:@48575.4]
  wire  accel_io_memStreams_scatters_0_cmd_valid; // @[Instantiator.scala 54:38:@48575.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0; // @[Instantiator.scala 54:38:@48575.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1; // @[Instantiator.scala 54:38:@48575.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2; // @[Instantiator.scala 54:38:@48575.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3; // @[Instantiator.scala 54:38:@48575.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4; // @[Instantiator.scala 54:38:@48575.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5; // @[Instantiator.scala 54:38:@48575.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6; // @[Instantiator.scala 54:38:@48575.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7; // @[Instantiator.scala 54:38:@48575.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8; // @[Instantiator.scala 54:38:@48575.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9; // @[Instantiator.scala 54:38:@48575.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10; // @[Instantiator.scala 54:38:@48575.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11; // @[Instantiator.scala 54:38:@48575.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12; // @[Instantiator.scala 54:38:@48575.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13; // @[Instantiator.scala 54:38:@48575.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14; // @[Instantiator.scala 54:38:@48575.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_0; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_1; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_2; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_3; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_4; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_5; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_6; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_7; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_8; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_9; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_10; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_11; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_12; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_13; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_14; // @[Instantiator.scala 54:38:@48575.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_15; // @[Instantiator.scala 54:38:@48575.4]
  wire  accel_io_memStreams_scatters_0_wresp_ready; // @[Instantiator.scala 54:38:@48575.4]
  wire  accel_io_memStreams_scatters_0_wresp_valid; // @[Instantiator.scala 54:38:@48575.4]
  wire  accel_io_memStreams_scatters_0_wresp_bits; // @[Instantiator.scala 54:38:@48575.4]
  wire  accel_io_heap_0_req_valid; // @[Instantiator.scala 54:38:@48575.4]
  wire  accel_io_heap_0_req_bits_allocDealloc; // @[Instantiator.scala 54:38:@48575.4]
  wire [63:0] accel_io_heap_0_req_bits_sizeAddr; // @[Instantiator.scala 54:38:@48575.4]
  wire  accel_io_heap_0_resp_valid; // @[Instantiator.scala 54:38:@48575.4]
  wire  accel_io_heap_0_resp_bits_allocDealloc; // @[Instantiator.scala 54:38:@48575.4]
  wire [63:0] accel_io_heap_0_resp_bits_sizeAddr; // @[Instantiator.scala 54:38:@48575.4]
  wire [63:0] accel_io_argIns_0; // @[Instantiator.scala 54:38:@48575.4]
  wire  accel_io_argOuts_0_port_ready; // @[Instantiator.scala 54:38:@48575.4]
  wire  accel_io_argOuts_0_port_valid; // @[Instantiator.scala 54:38:@48575.4]
  wire [63:0] accel_io_argOuts_0_port_bits; // @[Instantiator.scala 54:38:@48575.4]
  wire [63:0] accel_io_argOuts_0_echo; // @[Instantiator.scala 54:38:@48575.4]
  wire  FringeZynq_clock; // @[KCU1500.scala 21:24:@48713.4]
  wire  FringeZynq_reset; // @[KCU1500.scala 21:24:@48713.4]
  wire [31:0] FringeZynq_io_S_AXI_AWADDR; // @[KCU1500.scala 21:24:@48713.4]
  wire [2:0] FringeZynq_io_S_AXI_AWPROT; // @[KCU1500.scala 21:24:@48713.4]
  wire  FringeZynq_io_S_AXI_AWVALID; // @[KCU1500.scala 21:24:@48713.4]
  wire  FringeZynq_io_S_AXI_AWREADY; // @[KCU1500.scala 21:24:@48713.4]
  wire [31:0] FringeZynq_io_S_AXI_ARADDR; // @[KCU1500.scala 21:24:@48713.4]
  wire [2:0] FringeZynq_io_S_AXI_ARPROT; // @[KCU1500.scala 21:24:@48713.4]
  wire  FringeZynq_io_S_AXI_ARVALID; // @[KCU1500.scala 21:24:@48713.4]
  wire  FringeZynq_io_S_AXI_ARREADY; // @[KCU1500.scala 21:24:@48713.4]
  wire [31:0] FringeZynq_io_S_AXI_WDATA; // @[KCU1500.scala 21:24:@48713.4]
  wire [3:0] FringeZynq_io_S_AXI_WSTRB; // @[KCU1500.scala 21:24:@48713.4]
  wire  FringeZynq_io_S_AXI_WVALID; // @[KCU1500.scala 21:24:@48713.4]
  wire  FringeZynq_io_S_AXI_WREADY; // @[KCU1500.scala 21:24:@48713.4]
  wire [31:0] FringeZynq_io_S_AXI_RDATA; // @[KCU1500.scala 21:24:@48713.4]
  wire [1:0] FringeZynq_io_S_AXI_RRESP; // @[KCU1500.scala 21:24:@48713.4]
  wire  FringeZynq_io_S_AXI_RVALID; // @[KCU1500.scala 21:24:@48713.4]
  wire  FringeZynq_io_S_AXI_RREADY; // @[KCU1500.scala 21:24:@48713.4]
  wire [1:0] FringeZynq_io_S_AXI_BRESP; // @[KCU1500.scala 21:24:@48713.4]
  wire  FringeZynq_io_S_AXI_BVALID; // @[KCU1500.scala 21:24:@48713.4]
  wire  FringeZynq_io_S_AXI_BREADY; // @[KCU1500.scala 21:24:@48713.4]
  wire [7:0] FringeZynq_io_M_AXI_0_AWLEN; // @[KCU1500.scala 21:24:@48713.4]
  wire [7:0] FringeZynq_io_M_AXI_0_ARLEN; // @[KCU1500.scala 21:24:@48713.4]
  wire  FringeZynq_io_enable; // @[KCU1500.scala 21:24:@48713.4]
  wire  FringeZynq_io_done; // @[KCU1500.scala 21:24:@48713.4]
  wire  FringeZynq_io_reset; // @[KCU1500.scala 21:24:@48713.4]
  wire [63:0] FringeZynq_io_argIns_0; // @[KCU1500.scala 21:24:@48713.4]
  wire  FringeZynq_io_argOuts_0_valid; // @[KCU1500.scala 21:24:@48713.4]
  wire [63:0] FringeZynq_io_argOuts_0_bits; // @[KCU1500.scala 21:24:@48713.4]
  wire  FringeZynq_io_heap_0_req_valid; // @[KCU1500.scala 21:24:@48713.4]
  wire  FringeZynq_io_heap_0_req_bits_allocDealloc; // @[KCU1500.scala 21:24:@48713.4]
  wire [63:0] FringeZynq_io_heap_0_req_bits_sizeAddr; // @[KCU1500.scala 21:24:@48713.4]
  wire  FringeZynq_io_heap_0_resp_valid; // @[KCU1500.scala 21:24:@48713.4]
  wire  FringeZynq_io_heap_0_resp_bits_allocDealloc; // @[KCU1500.scala 21:24:@48713.4]
  wire [63:0] FringeZynq_io_heap_0_resp_bits_sizeAddr; // @[KCU1500.scala 21:24:@48713.4]
  AccelTop accel ( // @[Instantiator.scala 54:38:@48575.4]
    .clock(accel_clock),
    .reset(accel_reset),
    .io_enable(accel_io_enable),
    .io_done(accel_io_done),
    .io_reset(accel_io_reset),
    .io_memStreams_loads_0_cmd_ready(accel_io_memStreams_loads_0_cmd_ready),
    .io_memStreams_loads_0_cmd_valid(accel_io_memStreams_loads_0_cmd_valid),
    .io_memStreams_loads_0_cmd_bits_addr(accel_io_memStreams_loads_0_cmd_bits_addr),
    .io_memStreams_loads_0_cmd_bits_size(accel_io_memStreams_loads_0_cmd_bits_size),
    .io_memStreams_loads_0_data_ready(accel_io_memStreams_loads_0_data_ready),
    .io_memStreams_loads_0_data_valid(accel_io_memStreams_loads_0_data_valid),
    .io_memStreams_loads_0_data_bits_rdata_0(accel_io_memStreams_loads_0_data_bits_rdata_0),
    .io_memStreams_loads_0_data_bits_rdata_1(accel_io_memStreams_loads_0_data_bits_rdata_1),
    .io_memStreams_loads_0_data_bits_rdata_2(accel_io_memStreams_loads_0_data_bits_rdata_2),
    .io_memStreams_loads_0_data_bits_rdata_3(accel_io_memStreams_loads_0_data_bits_rdata_3),
    .io_memStreams_loads_0_data_bits_rdata_4(accel_io_memStreams_loads_0_data_bits_rdata_4),
    .io_memStreams_loads_0_data_bits_rdata_5(accel_io_memStreams_loads_0_data_bits_rdata_5),
    .io_memStreams_loads_0_data_bits_rdata_6(accel_io_memStreams_loads_0_data_bits_rdata_6),
    .io_memStreams_loads_0_data_bits_rdata_7(accel_io_memStreams_loads_0_data_bits_rdata_7),
    .io_memStreams_loads_0_data_bits_rdata_8(accel_io_memStreams_loads_0_data_bits_rdata_8),
    .io_memStreams_loads_0_data_bits_rdata_9(accel_io_memStreams_loads_0_data_bits_rdata_9),
    .io_memStreams_loads_0_data_bits_rdata_10(accel_io_memStreams_loads_0_data_bits_rdata_10),
    .io_memStreams_loads_0_data_bits_rdata_11(accel_io_memStreams_loads_0_data_bits_rdata_11),
    .io_memStreams_loads_0_data_bits_rdata_12(accel_io_memStreams_loads_0_data_bits_rdata_12),
    .io_memStreams_loads_0_data_bits_rdata_13(accel_io_memStreams_loads_0_data_bits_rdata_13),
    .io_memStreams_loads_0_data_bits_rdata_14(accel_io_memStreams_loads_0_data_bits_rdata_14),
    .io_memStreams_loads_0_data_bits_rdata_15(accel_io_memStreams_loads_0_data_bits_rdata_15),
    .io_memStreams_stores_0_cmd_ready(accel_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(accel_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(accel_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(accel_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(accel_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(accel_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(accel_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wdata_1(accel_io_memStreams_stores_0_data_bits_wdata_1),
    .io_memStreams_stores_0_data_bits_wdata_2(accel_io_memStreams_stores_0_data_bits_wdata_2),
    .io_memStreams_stores_0_data_bits_wdata_3(accel_io_memStreams_stores_0_data_bits_wdata_3),
    .io_memStreams_stores_0_data_bits_wdata_4(accel_io_memStreams_stores_0_data_bits_wdata_4),
    .io_memStreams_stores_0_data_bits_wdata_5(accel_io_memStreams_stores_0_data_bits_wdata_5),
    .io_memStreams_stores_0_data_bits_wdata_6(accel_io_memStreams_stores_0_data_bits_wdata_6),
    .io_memStreams_stores_0_data_bits_wdata_7(accel_io_memStreams_stores_0_data_bits_wdata_7),
    .io_memStreams_stores_0_data_bits_wdata_8(accel_io_memStreams_stores_0_data_bits_wdata_8),
    .io_memStreams_stores_0_data_bits_wdata_9(accel_io_memStreams_stores_0_data_bits_wdata_9),
    .io_memStreams_stores_0_data_bits_wdata_10(accel_io_memStreams_stores_0_data_bits_wdata_10),
    .io_memStreams_stores_0_data_bits_wdata_11(accel_io_memStreams_stores_0_data_bits_wdata_11),
    .io_memStreams_stores_0_data_bits_wdata_12(accel_io_memStreams_stores_0_data_bits_wdata_12),
    .io_memStreams_stores_0_data_bits_wdata_13(accel_io_memStreams_stores_0_data_bits_wdata_13),
    .io_memStreams_stores_0_data_bits_wdata_14(accel_io_memStreams_stores_0_data_bits_wdata_14),
    .io_memStreams_stores_0_data_bits_wdata_15(accel_io_memStreams_stores_0_data_bits_wdata_15),
    .io_memStreams_stores_0_data_bits_wstrb(accel_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(accel_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(accel_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(accel_io_memStreams_stores_0_wresp_bits),
    .io_memStreams_gathers_0_cmd_ready(accel_io_memStreams_gathers_0_cmd_ready),
    .io_memStreams_gathers_0_cmd_valid(accel_io_memStreams_gathers_0_cmd_valid),
    .io_memStreams_gathers_0_cmd_bits_addr_0(accel_io_memStreams_gathers_0_cmd_bits_addr_0),
    .io_memStreams_gathers_0_cmd_bits_addr_1(accel_io_memStreams_gathers_0_cmd_bits_addr_1),
    .io_memStreams_gathers_0_cmd_bits_addr_2(accel_io_memStreams_gathers_0_cmd_bits_addr_2),
    .io_memStreams_gathers_0_cmd_bits_addr_3(accel_io_memStreams_gathers_0_cmd_bits_addr_3),
    .io_memStreams_gathers_0_cmd_bits_addr_4(accel_io_memStreams_gathers_0_cmd_bits_addr_4),
    .io_memStreams_gathers_0_cmd_bits_addr_5(accel_io_memStreams_gathers_0_cmd_bits_addr_5),
    .io_memStreams_gathers_0_cmd_bits_addr_6(accel_io_memStreams_gathers_0_cmd_bits_addr_6),
    .io_memStreams_gathers_0_cmd_bits_addr_7(accel_io_memStreams_gathers_0_cmd_bits_addr_7),
    .io_memStreams_gathers_0_cmd_bits_addr_8(accel_io_memStreams_gathers_0_cmd_bits_addr_8),
    .io_memStreams_gathers_0_cmd_bits_addr_9(accel_io_memStreams_gathers_0_cmd_bits_addr_9),
    .io_memStreams_gathers_0_cmd_bits_addr_10(accel_io_memStreams_gathers_0_cmd_bits_addr_10),
    .io_memStreams_gathers_0_cmd_bits_addr_11(accel_io_memStreams_gathers_0_cmd_bits_addr_11),
    .io_memStreams_gathers_0_cmd_bits_addr_12(accel_io_memStreams_gathers_0_cmd_bits_addr_12),
    .io_memStreams_gathers_0_cmd_bits_addr_13(accel_io_memStreams_gathers_0_cmd_bits_addr_13),
    .io_memStreams_gathers_0_cmd_bits_addr_14(accel_io_memStreams_gathers_0_cmd_bits_addr_14),
    .io_memStreams_gathers_0_cmd_bits_addr_15(accel_io_memStreams_gathers_0_cmd_bits_addr_15),
    .io_memStreams_gathers_0_data_ready(accel_io_memStreams_gathers_0_data_ready),
    .io_memStreams_gathers_0_data_valid(accel_io_memStreams_gathers_0_data_valid),
    .io_memStreams_gathers_0_data_bits_0(accel_io_memStreams_gathers_0_data_bits_0),
    .io_memStreams_gathers_0_data_bits_1(accel_io_memStreams_gathers_0_data_bits_1),
    .io_memStreams_gathers_0_data_bits_2(accel_io_memStreams_gathers_0_data_bits_2),
    .io_memStreams_gathers_0_data_bits_3(accel_io_memStreams_gathers_0_data_bits_3),
    .io_memStreams_gathers_0_data_bits_4(accel_io_memStreams_gathers_0_data_bits_4),
    .io_memStreams_gathers_0_data_bits_5(accel_io_memStreams_gathers_0_data_bits_5),
    .io_memStreams_gathers_0_data_bits_6(accel_io_memStreams_gathers_0_data_bits_6),
    .io_memStreams_gathers_0_data_bits_7(accel_io_memStreams_gathers_0_data_bits_7),
    .io_memStreams_gathers_0_data_bits_8(accel_io_memStreams_gathers_0_data_bits_8),
    .io_memStreams_gathers_0_data_bits_9(accel_io_memStreams_gathers_0_data_bits_9),
    .io_memStreams_gathers_0_data_bits_10(accel_io_memStreams_gathers_0_data_bits_10),
    .io_memStreams_gathers_0_data_bits_11(accel_io_memStreams_gathers_0_data_bits_11),
    .io_memStreams_gathers_0_data_bits_12(accel_io_memStreams_gathers_0_data_bits_12),
    .io_memStreams_gathers_0_data_bits_13(accel_io_memStreams_gathers_0_data_bits_13),
    .io_memStreams_gathers_0_data_bits_14(accel_io_memStreams_gathers_0_data_bits_14),
    .io_memStreams_gathers_0_data_bits_15(accel_io_memStreams_gathers_0_data_bits_15),
    .io_memStreams_scatters_0_cmd_ready(accel_io_memStreams_scatters_0_cmd_ready),
    .io_memStreams_scatters_0_cmd_valid(accel_io_memStreams_scatters_0_cmd_valid),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_0(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_1(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_2(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_3(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_4(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_5(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_6(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_7(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_8(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_9(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_10(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_11(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_12(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_13(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_14(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_15(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15),
    .io_memStreams_scatters_0_cmd_bits_wdata_0(accel_io_memStreams_scatters_0_cmd_bits_wdata_0),
    .io_memStreams_scatters_0_cmd_bits_wdata_1(accel_io_memStreams_scatters_0_cmd_bits_wdata_1),
    .io_memStreams_scatters_0_cmd_bits_wdata_2(accel_io_memStreams_scatters_0_cmd_bits_wdata_2),
    .io_memStreams_scatters_0_cmd_bits_wdata_3(accel_io_memStreams_scatters_0_cmd_bits_wdata_3),
    .io_memStreams_scatters_0_cmd_bits_wdata_4(accel_io_memStreams_scatters_0_cmd_bits_wdata_4),
    .io_memStreams_scatters_0_cmd_bits_wdata_5(accel_io_memStreams_scatters_0_cmd_bits_wdata_5),
    .io_memStreams_scatters_0_cmd_bits_wdata_6(accel_io_memStreams_scatters_0_cmd_bits_wdata_6),
    .io_memStreams_scatters_0_cmd_bits_wdata_7(accel_io_memStreams_scatters_0_cmd_bits_wdata_7),
    .io_memStreams_scatters_0_cmd_bits_wdata_8(accel_io_memStreams_scatters_0_cmd_bits_wdata_8),
    .io_memStreams_scatters_0_cmd_bits_wdata_9(accel_io_memStreams_scatters_0_cmd_bits_wdata_9),
    .io_memStreams_scatters_0_cmd_bits_wdata_10(accel_io_memStreams_scatters_0_cmd_bits_wdata_10),
    .io_memStreams_scatters_0_cmd_bits_wdata_11(accel_io_memStreams_scatters_0_cmd_bits_wdata_11),
    .io_memStreams_scatters_0_cmd_bits_wdata_12(accel_io_memStreams_scatters_0_cmd_bits_wdata_12),
    .io_memStreams_scatters_0_cmd_bits_wdata_13(accel_io_memStreams_scatters_0_cmd_bits_wdata_13),
    .io_memStreams_scatters_0_cmd_bits_wdata_14(accel_io_memStreams_scatters_0_cmd_bits_wdata_14),
    .io_memStreams_scatters_0_cmd_bits_wdata_15(accel_io_memStreams_scatters_0_cmd_bits_wdata_15),
    .io_memStreams_scatters_0_wresp_ready(accel_io_memStreams_scatters_0_wresp_ready),
    .io_memStreams_scatters_0_wresp_valid(accel_io_memStreams_scatters_0_wresp_valid),
    .io_memStreams_scatters_0_wresp_bits(accel_io_memStreams_scatters_0_wresp_bits),
    .io_heap_0_req_valid(accel_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(accel_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(accel_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(accel_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(accel_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(accel_io_heap_0_resp_bits_sizeAddr),
    .io_argIns_0(accel_io_argIns_0),
    .io_argOuts_0_port_ready(accel_io_argOuts_0_port_ready),
    .io_argOuts_0_port_valid(accel_io_argOuts_0_port_valid),
    .io_argOuts_0_port_bits(accel_io_argOuts_0_port_bits),
    .io_argOuts_0_echo(accel_io_argOuts_0_echo)
  );
  FringeZynq FringeZynq ( // @[KCU1500.scala 21:24:@48713.4]
    .clock(FringeZynq_clock),
    .reset(FringeZynq_reset),
    .io_S_AXI_AWADDR(FringeZynq_io_S_AXI_AWADDR),
    .io_S_AXI_AWPROT(FringeZynq_io_S_AXI_AWPROT),
    .io_S_AXI_AWVALID(FringeZynq_io_S_AXI_AWVALID),
    .io_S_AXI_AWREADY(FringeZynq_io_S_AXI_AWREADY),
    .io_S_AXI_ARADDR(FringeZynq_io_S_AXI_ARADDR),
    .io_S_AXI_ARPROT(FringeZynq_io_S_AXI_ARPROT),
    .io_S_AXI_ARVALID(FringeZynq_io_S_AXI_ARVALID),
    .io_S_AXI_ARREADY(FringeZynq_io_S_AXI_ARREADY),
    .io_S_AXI_WDATA(FringeZynq_io_S_AXI_WDATA),
    .io_S_AXI_WSTRB(FringeZynq_io_S_AXI_WSTRB),
    .io_S_AXI_WVALID(FringeZynq_io_S_AXI_WVALID),
    .io_S_AXI_WREADY(FringeZynq_io_S_AXI_WREADY),
    .io_S_AXI_RDATA(FringeZynq_io_S_AXI_RDATA),
    .io_S_AXI_RRESP(FringeZynq_io_S_AXI_RRESP),
    .io_S_AXI_RVALID(FringeZynq_io_S_AXI_RVALID),
    .io_S_AXI_RREADY(FringeZynq_io_S_AXI_RREADY),
    .io_S_AXI_BRESP(FringeZynq_io_S_AXI_BRESP),
    .io_S_AXI_BVALID(FringeZynq_io_S_AXI_BVALID),
    .io_S_AXI_BREADY(FringeZynq_io_S_AXI_BREADY),
    .io_M_AXI_0_AWLEN(FringeZynq_io_M_AXI_0_AWLEN),
    .io_M_AXI_0_ARLEN(FringeZynq_io_M_AXI_0_ARLEN),
    .io_enable(FringeZynq_io_enable),
    .io_done(FringeZynq_io_done),
    .io_reset(FringeZynq_io_reset),
    .io_argIns_0(FringeZynq_io_argIns_0),
    .io_argOuts_0_valid(FringeZynq_io_argOuts_0_valid),
    .io_argOuts_0_bits(FringeZynq_io_argOuts_0_bits),
    .io_heap_0_req_valid(FringeZynq_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(FringeZynq_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(FringeZynq_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(FringeZynq_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(FringeZynq_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(FringeZynq_io_heap_0_resp_bits_sizeAddr)
  );
  assign io_rdata = 1'h0;
  assign io_S_AXI_AWREADY = FringeZynq_io_S_AXI_AWREADY; // @[KCU1500.scala 24:21:@48731.4]
  assign io_S_AXI_ARREADY = FringeZynq_io_S_AXI_ARREADY; // @[KCU1500.scala 24:21:@48727.4]
  assign io_S_AXI_WREADY = FringeZynq_io_S_AXI_WREADY; // @[KCU1500.scala 24:21:@48723.4]
  assign io_S_AXI_RDATA = FringeZynq_io_S_AXI_RDATA; // @[KCU1500.scala 24:21:@48722.4]
  assign io_S_AXI_RRESP = FringeZynq_io_S_AXI_RRESP; // @[KCU1500.scala 24:21:@48721.4]
  assign io_S_AXI_RVALID = FringeZynq_io_S_AXI_RVALID; // @[KCU1500.scala 24:21:@48720.4]
  assign io_S_AXI_BRESP = FringeZynq_io_S_AXI_BRESP; // @[KCU1500.scala 24:21:@48718.4]
  assign io_S_AXI_BVALID = FringeZynq_io_S_AXI_BVALID; // @[KCU1500.scala 24:21:@48717.4]
  assign io_M_AXI_0_AWID = 4'h0; // @[KCU1500.scala 27:14:@48775.4]
  assign io_M_AXI_0_AWUSER = 4'h0; // @[KCU1500.scala 27:14:@48774.4]
  assign io_M_AXI_0_AWADDR = 32'h0; // @[KCU1500.scala 27:14:@48773.4]
  assign io_M_AXI_0_AWLEN = FringeZynq_io_M_AXI_0_AWLEN; // @[KCU1500.scala 27:14:@48772.4]
  assign io_M_AXI_0_AWSIZE = 3'h6; // @[KCU1500.scala 27:14:@48771.4]
  assign io_M_AXI_0_AWBURST = 2'h1; // @[KCU1500.scala 27:14:@48770.4]
  assign io_M_AXI_0_AWLOCK = 1'h0; // @[KCU1500.scala 27:14:@48769.4]
  assign io_M_AXI_0_AWCACHE = 4'h3; // @[KCU1500.scala 27:14:@48768.4]
  assign io_M_AXI_0_AWPROT = 3'h0; // @[KCU1500.scala 27:14:@48767.4]
  assign io_M_AXI_0_AWQOS = 4'h0; // @[KCU1500.scala 27:14:@48766.4]
  assign io_M_AXI_0_AWVALID = 1'h0; // @[KCU1500.scala 27:14:@48765.4]
  assign io_M_AXI_0_ARID = 4'h0; // @[KCU1500.scala 27:14:@48763.4]
  assign io_M_AXI_0_ARUSER = 4'h0; // @[KCU1500.scala 27:14:@48762.4]
  assign io_M_AXI_0_ARADDR = 32'h0; // @[KCU1500.scala 27:14:@48761.4]
  assign io_M_AXI_0_ARLEN = FringeZynq_io_M_AXI_0_ARLEN; // @[KCU1500.scala 27:14:@48760.4]
  assign io_M_AXI_0_ARSIZE = 3'h6; // @[KCU1500.scala 27:14:@48759.4]
  assign io_M_AXI_0_ARBURST = 2'h1; // @[KCU1500.scala 27:14:@48758.4]
  assign io_M_AXI_0_ARLOCK = 1'h0; // @[KCU1500.scala 27:14:@48757.4]
  assign io_M_AXI_0_ARCACHE = 4'h3; // @[KCU1500.scala 27:14:@48756.4]
  assign io_M_AXI_0_ARPROT = 3'h0; // @[KCU1500.scala 27:14:@48755.4]
  assign io_M_AXI_0_ARQOS = 4'h0; // @[KCU1500.scala 27:14:@48754.4]
  assign io_M_AXI_0_ARVALID = 1'h0; // @[KCU1500.scala 27:14:@48753.4]
  assign io_M_AXI_0_WDATA = 512'h0; // @[KCU1500.scala 27:14:@48751.4]
  assign io_M_AXI_0_WSTRB = 64'h0; // @[KCU1500.scala 27:14:@48750.4]
  assign io_M_AXI_0_WLAST = 1'h0; // @[KCU1500.scala 27:14:@48749.4]
  assign io_M_AXI_0_WVALID = 1'h0; // @[KCU1500.scala 27:14:@48748.4]
  assign io_M_AXI_0_RREADY = 1'h0; // @[KCU1500.scala 27:14:@48740.4]
  assign io_M_AXI_0_BREADY = 1'h0; // @[KCU1500.scala 27:14:@48735.4]
  assign accel_clock = clock; // @[:@48576.4]
  assign accel_reset = FringeZynq_io_reset; // @[:@48577.4 KCU1500.scala 57:17:@49077.4]
  assign accel_io_enable = FringeZynq_io_enable; // @[KCU1500.scala 54:21:@49073.4]
  assign accel_io_reset = 1'h0;
  assign accel_io_memStreams_loads_0_cmd_ready = 1'h0; // @[KCU1500.scala 52:26:@49066.4]
  assign accel_io_memStreams_loads_0_data_valid = 1'h0; // @[KCU1500.scala 52:26:@49061.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_0 = 32'h0; // @[KCU1500.scala 52:26:@49045.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_1 = 32'h0; // @[KCU1500.scala 52:26:@49046.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_2 = 32'h0; // @[KCU1500.scala 52:26:@49047.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_3 = 32'h0; // @[KCU1500.scala 52:26:@49048.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_4 = 32'h0; // @[KCU1500.scala 52:26:@49049.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_5 = 32'h0; // @[KCU1500.scala 52:26:@49050.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_6 = 32'h0; // @[KCU1500.scala 52:26:@49051.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_7 = 32'h0; // @[KCU1500.scala 52:26:@49052.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_8 = 32'h0; // @[KCU1500.scala 52:26:@49053.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_9 = 32'h0; // @[KCU1500.scala 52:26:@49054.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_10 = 32'h0; // @[KCU1500.scala 52:26:@49055.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_11 = 32'h0; // @[KCU1500.scala 52:26:@49056.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_12 = 32'h0; // @[KCU1500.scala 52:26:@49057.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_13 = 32'h0; // @[KCU1500.scala 52:26:@49058.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_14 = 32'h0; // @[KCU1500.scala 52:26:@49059.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_15 = 32'h0; // @[KCU1500.scala 52:26:@49060.4]
  assign accel_io_memStreams_stores_0_cmd_ready = 1'h0; // @[KCU1500.scala 52:26:@49044.4]
  assign accel_io_memStreams_stores_0_data_ready = 1'h0; // @[KCU1500.scala 52:26:@49040.4]
  assign accel_io_memStreams_stores_0_wresp_valid = 1'h0; // @[KCU1500.scala 52:26:@49020.4]
  assign accel_io_memStreams_stores_0_wresp_bits = 1'h0; // @[KCU1500.scala 52:26:@49019.4]
  assign accel_io_memStreams_gathers_0_cmd_ready = 1'h0; // @[KCU1500.scala 52:26:@49018.4]
  assign accel_io_memStreams_gathers_0_data_valid = 1'h0; // @[KCU1500.scala 52:26:@48999.4]
  assign accel_io_memStreams_gathers_0_data_bits_0 = 32'h0; // @[KCU1500.scala 52:26:@48983.4]
  assign accel_io_memStreams_gathers_0_data_bits_1 = 32'h0; // @[KCU1500.scala 52:26:@48984.4]
  assign accel_io_memStreams_gathers_0_data_bits_2 = 32'h0; // @[KCU1500.scala 52:26:@48985.4]
  assign accel_io_memStreams_gathers_0_data_bits_3 = 32'h0; // @[KCU1500.scala 52:26:@48986.4]
  assign accel_io_memStreams_gathers_0_data_bits_4 = 32'h0; // @[KCU1500.scala 52:26:@48987.4]
  assign accel_io_memStreams_gathers_0_data_bits_5 = 32'h0; // @[KCU1500.scala 52:26:@48988.4]
  assign accel_io_memStreams_gathers_0_data_bits_6 = 32'h0; // @[KCU1500.scala 52:26:@48989.4]
  assign accel_io_memStreams_gathers_0_data_bits_7 = 32'h0; // @[KCU1500.scala 52:26:@48990.4]
  assign accel_io_memStreams_gathers_0_data_bits_8 = 32'h0; // @[KCU1500.scala 52:26:@48991.4]
  assign accel_io_memStreams_gathers_0_data_bits_9 = 32'h0; // @[KCU1500.scala 52:26:@48992.4]
  assign accel_io_memStreams_gathers_0_data_bits_10 = 32'h0; // @[KCU1500.scala 52:26:@48993.4]
  assign accel_io_memStreams_gathers_0_data_bits_11 = 32'h0; // @[KCU1500.scala 52:26:@48994.4]
  assign accel_io_memStreams_gathers_0_data_bits_12 = 32'h0; // @[KCU1500.scala 52:26:@48995.4]
  assign accel_io_memStreams_gathers_0_data_bits_13 = 32'h0; // @[KCU1500.scala 52:26:@48996.4]
  assign accel_io_memStreams_gathers_0_data_bits_14 = 32'h0; // @[KCU1500.scala 52:26:@48997.4]
  assign accel_io_memStreams_gathers_0_data_bits_15 = 32'h0; // @[KCU1500.scala 52:26:@48998.4]
  assign accel_io_memStreams_scatters_0_cmd_ready = 1'h0; // @[KCU1500.scala 52:26:@48982.4]
  assign accel_io_memStreams_scatters_0_wresp_valid = 1'h0; // @[KCU1500.scala 52:26:@48947.4]
  assign accel_io_memStreams_scatters_0_wresp_bits = 1'h0; // @[KCU1500.scala 52:26:@48946.4]
  assign accel_io_heap_0_resp_valid = FringeZynq_io_heap_0_resp_valid; // @[KCU1500.scala 53:20:@49069.4]
  assign accel_io_heap_0_resp_bits_allocDealloc = FringeZynq_io_heap_0_resp_bits_allocDealloc; // @[KCU1500.scala 53:20:@49068.4]
  assign accel_io_heap_0_resp_bits_sizeAddr = FringeZynq_io_heap_0_resp_bits_sizeAddr; // @[KCU1500.scala 53:20:@49067.4]
  assign accel_io_argIns_0 = FringeZynq_io_argIns_0; // @[KCU1500.scala 37:21:@48941.4]
  assign accel_io_argOuts_0_port_ready = 1'h0;
  assign accel_io_argOuts_0_echo = 64'h0; // @[KCU1500.scala 43:24:@48944.4]
  assign FringeZynq_clock = clock; // @[:@48714.4]
  assign FringeZynq_reset = reset; // @[:@48715.4 KCU1500.scala 56:18:@49076.4]
  assign FringeZynq_io_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[KCU1500.scala 24:21:@48734.4]
  assign FringeZynq_io_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[KCU1500.scala 24:21:@48733.4]
  assign FringeZynq_io_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[KCU1500.scala 24:21:@48732.4]
  assign FringeZynq_io_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[KCU1500.scala 24:21:@48730.4]
  assign FringeZynq_io_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[KCU1500.scala 24:21:@48729.4]
  assign FringeZynq_io_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[KCU1500.scala 24:21:@48728.4]
  assign FringeZynq_io_S_AXI_WDATA = io_S_AXI_WDATA; // @[KCU1500.scala 24:21:@48726.4]
  assign FringeZynq_io_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[KCU1500.scala 24:21:@48725.4]
  assign FringeZynq_io_S_AXI_WVALID = io_S_AXI_WVALID; // @[KCU1500.scala 24:21:@48724.4]
  assign FringeZynq_io_S_AXI_RREADY = io_S_AXI_RREADY; // @[KCU1500.scala 24:21:@48719.4]
  assign FringeZynq_io_S_AXI_BREADY = io_S_AXI_BREADY; // @[KCU1500.scala 24:21:@48716.4]
  assign FringeZynq_io_done = accel_io_done; // @[KCU1500.scala 55:20:@49074.4]
  assign FringeZynq_io_argOuts_0_valid = accel_io_argOuts_0_port_valid; // @[KCU1500.scala 40:26:@48943.4]
  assign FringeZynq_io_argOuts_0_bits = accel_io_argOuts_0_port_bits; // @[KCU1500.scala 39:25:@48942.4]
  assign FringeZynq_io_heap_0_req_valid = accel_io_heap_0_req_valid; // @[KCU1500.scala 53:20:@49072.4]
  assign FringeZynq_io_heap_0_req_bits_allocDealloc = accel_io_heap_0_req_bits_allocDealloc; // @[KCU1500.scala 53:20:@49071.4]
  assign FringeZynq_io_heap_0_req_bits_sizeAddr = accel_io_heap_0_req_bits_sizeAddr; // @[KCU1500.scala 53:20:@49070.4]
endmodule
module SRAMVerilogAWS
#(
    parameter WORDS = 1024,
    parameter AWIDTH = 10,
    parameter DWIDTH = 32)
(
    input clk,
    input [AWIDTH-1:0] raddr,
    input [AWIDTH-1:0] waddr,
    input raddrEn,
    input waddrEn,
    input wen,
    input [DWIDTH-1:0] wdata,
    input backpressure,
    output reg [DWIDTH-1:0] rdata
);

    reg [DWIDTH-1:0] mem [0:WORDS-1];

    always @(posedge clk) begin
      if (wen) mem[waddr] <= wdata;
      if (backpressure) rdata <= mem[raddr];
    end

endmodule
