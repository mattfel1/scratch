module FF( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  output [31:0] io_rPort_0_output_0, // @[:@6.4]
  input  [31:0] io_wPort_0_data_0, // @[:@6.4]
  input         io_wPort_0_reset, // @[:@6.4]
  input         io_wPort_0_en_0 // @[:@6.4]
);
  reg [31:0] ff; // @[MemPrimitives.scala 173:19:@21.4]
  reg [31:0] _RAND_0;
  wire [31:0] _T_68; // @[MemPrimitives.scala 177:32:@23.4]
  wire [31:0] _T_69; // @[MemPrimitives.scala 177:12:@24.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 177:32:@23.4]
  assign _T_69 = io_wPort_0_reset ? 32'h0 : _T_68; // @[MemPrimitives.scala 177:12:@24.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 178:34:@26.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 32'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 32'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SRFF( // @[:@28.2]
  input   clock, // @[:@29.4]
  input   reset, // @[:@30.4]
  input   io_input_set, // @[:@31.4]
  input   io_input_reset, // @[:@31.4]
  input   io_input_asyn_reset, // @[:@31.4]
  output  io_output // @[:@31.4]
);
  reg  _T_15; // @[SRFF.scala 20:21:@33.4]
  reg [31:0] _RAND_0;
  wire  _T_19; // @[SRFF.scala 21:74:@34.4]
  wire  _T_20; // @[SRFF.scala 21:48:@35.4]
  wire  _T_21; // @[SRFF.scala 21:14:@36.4]
  assign _T_19 = io_input_reset ? 1'h0 : _T_15; // @[SRFF.scala 21:74:@34.4]
  assign _T_20 = io_input_set ? 1'h1 : _T_19; // @[SRFF.scala 21:48:@35.4]
  assign _T_21 = io_input_asyn_reset ? 1'h0 : _T_20; // @[SRFF.scala 21:14:@36.4]
  assign io_output = io_input_asyn_reset ? 1'h0 : _T_15; // @[SRFF.scala 22:15:@39.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_15 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_15 <= 1'h0;
    end else begin
      if (io_input_asyn_reset) begin
        _T_15 <= 1'h0;
      end else begin
        if (io_input_set) begin
          _T_15 <= 1'h1;
        end else begin
          if (io_input_reset) begin
            _T_15 <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module SingleCounter( // @[:@41.2]
  input   clock, // @[:@42.4]
  input   reset, // @[:@43.4]
  input   io_input_reset, // @[:@44.4]
  output  io_output_done // @[:@44.4]
);
  wire  bases_0_clock; // @[Counter.scala 253:53:@57.4]
  wire  bases_0_reset; // @[Counter.scala 253:53:@57.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 253:53:@57.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 253:53:@57.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 253:53:@57.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 253:53:@57.4]
  wire  SRFF_clock; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_reset; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_input_set; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_output; // @[Counter.scala 255:22:@73.4]
  wire [31:0] _T_48; // @[Counter.scala 279:52:@101.4]
  wire [32:0] _T_50; // @[Counter.scala 283:33:@102.4]
  wire [31:0] _T_51; // @[Counter.scala 283:33:@103.4]
  wire [31:0] _T_52; // @[Counter.scala 283:33:@104.4]
  wire  _T_57; // @[Counter.scala 285:18:@106.4]
  wire [31:0] _T_68; // @[Counter.scala 291:115:@114.4]
  wire [31:0] _T_71; // @[Counter.scala 291:152:@117.4]
  wire [31:0] _T_72; // @[Counter.scala 291:74:@118.4]
  FF bases_0 ( // @[Counter.scala 253:53:@57.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 255:22:@73.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 279:52:@101.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@102.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@103.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 283:33:@104.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh1); // @[Counter.scala 285:18:@106.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 291:115:@114.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 291:152:@117.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 291:74:@118.4]
  assign io_output_done = $signed(_T_52) >= $signed(32'sh1); // @[Counter.scala 325:20:@127.4]
  assign bases_0_clock = clock; // @[:@58.4]
  assign bases_0_reset = reset; // @[:@59.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 291:31:@120.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 273:27:@99.4]
  assign bases_0_io_wPort_0_en_0 = 1'h1; // @[Counter.scala 276:29:@100.4]
  assign SRFF_clock = clock; // @[:@74.4]
  assign SRFF_reset = reset; // @[:@75.4]
  assign SRFF_io_input_set = io_input_reset == 1'h0; // @[Counter.scala 256:23:@78.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 257:25:@80.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 258:30:@81.4]
endmodule
module RetimeWrapper( // @[:@144.2]
  input   clock, // @[:@145.4]
  input   reset, // @[:@146.4]
  input   io_flow, // @[:@147.4]
  input   io_in, // @[:@147.4]
  output  io_out // @[:@147.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@149.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@149.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@162.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@161.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@160.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@159.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@158.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@156.4]
endmodule
module RootController_sm( // @[:@351.2]
  input   clock, // @[:@352.4]
  input   reset, // @[:@353.4]
  input   io_enable, // @[:@354.4]
  output  io_done, // @[:@354.4]
  input   io_rst, // @[:@354.4]
  input   io_ctrDone, // @[:@354.4]
  output  io_ctrInc, // @[:@354.4]
  input   io_doneIn_0, // @[:@354.4]
  input   io_doneIn_1, // @[:@354.4]
  output  io_enableOut_0, // @[:@354.4]
  output  io_enableOut_1, // @[:@354.4]
  output  io_childAck_0, // @[:@354.4]
  output  io_childAck_1 // @[:@354.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@357.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@357.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@357.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@357.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@357.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@357.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@360.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@360.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@360.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@360.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@360.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@360.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@363.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@363.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@363.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@363.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@363.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@363.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@366.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@366.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@366.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@366.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@366.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@366.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@395.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@395.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@395.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@395.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@395.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@395.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@398.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@398.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@398.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@398.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@398.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@398.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@427.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@427.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@427.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@427.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@427.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@523.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@523.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@523.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@523.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@523.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@540.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@540.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@540.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@540.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@540.4]
  wire  allDone; // @[Controllers.scala 80:47:@369.4]
  wire  _T_77; // @[Controllers.scala 81:26:@370.4]
  wire  finished; // @[Controllers.scala 81:37:@371.4]
  wire  synchronize; // @[package.scala 96:25:@432.4 package.scala 96:25:@433.4]
  wire  _T_144; // @[Controllers.scala 128:33:@441.4]
  wire  _T_146; // @[Controllers.scala 128:54:@442.4]
  wire  _T_147; // @[Controllers.scala 128:52:@443.4]
  wire  _T_148; // @[Controllers.scala 128:66:@444.4]
  wire  _T_150; // @[Controllers.scala 128:98:@446.4]
  wire  _T_151; // @[Controllers.scala 128:96:@447.4]
  wire  _T_153; // @[Controllers.scala 128:123:@448.4]
  wire  _T_155; // @[Controllers.scala 129:48:@451.4]
  wire  _T_160; // @[Controllers.scala 130:52:@456.4]
  wire  _T_161; // @[Controllers.scala 130:50:@457.4]
  wire  _T_169; // @[Controllers.scala 130:129:@463.4]
  wire  _T_172; // @[Controllers.scala 131:45:@466.4]
  wire  _T_175; // @[Controllers.scala 135:80:@470.4]
  wire  _T_176; // @[Controllers.scala 135:78:@471.4]
  wire  _T_178; // @[Controllers.scala 135:105:@472.4]
  wire  _T_179; // @[Controllers.scala 135:103:@473.4]
  wire  _T_180; // @[Controllers.scala 135:119:@474.4]
  wire  _T_182; // @[Controllers.scala 135:51:@476.4]
  wire  _T_205; // @[Controllers.scala 213:68:@501.4]
  wire  _T_207; // @[Controllers.scala 213:90:@503.4]
  wire  _T_209; // @[Controllers.scala 213:132:@505.4]
  wire  _T_210; // @[Controllers.scala 213:130:@506.4]
  wire  _T_211; // @[Controllers.scala 213:156:@507.4]
  wire  _T_213; // @[Controllers.scala 213:68:@510.4]
  wire  _T_215; // @[Controllers.scala 213:90:@512.4]
  wire  _T_222; // @[package.scala 100:49:@518.4]
  reg  _T_225; // @[package.scala 48:56:@519.4]
  reg [31:0] _RAND_0;
  reg  _T_239; // @[package.scala 48:56:@537.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@357.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@360.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@363.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@366.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@395.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@398.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@427.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@523.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@540.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  assign allDone = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@369.4]
  assign _T_77 = allDone | io_done; // @[Controllers.scala 81:26:@370.4]
  assign finished = _T_77 | done_1_io_input_set; // @[Controllers.scala 81:37:@371.4]
  assign synchronize = RetimeWrapper_io_out; // @[package.scala 96:25:@432.4 package.scala 96:25:@433.4]
  assign _T_144 = done_0_io_output == 1'h0; // @[Controllers.scala 128:33:@441.4]
  assign _T_146 = io_ctrDone == 1'h0; // @[Controllers.scala 128:54:@442.4]
  assign _T_147 = _T_144 & _T_146; // @[Controllers.scala 128:52:@443.4]
  assign _T_148 = _T_147 & io_enable; // @[Controllers.scala 128:66:@444.4]
  assign _T_150 = ~ iterDone_0_io_output; // @[Controllers.scala 128:98:@446.4]
  assign _T_151 = _T_148 & _T_150; // @[Controllers.scala 128:96:@447.4]
  assign _T_153 = io_doneIn_0 == 1'h0; // @[Controllers.scala 128:123:@448.4]
  assign _T_155 = io_doneIn_0 | io_rst; // @[Controllers.scala 129:48:@451.4]
  assign _T_160 = synchronize == 1'h0; // @[Controllers.scala 130:52:@456.4]
  assign _T_161 = io_doneIn_0 & _T_160; // @[Controllers.scala 130:50:@457.4]
  assign _T_169 = finished == 1'h0; // @[Controllers.scala 130:129:@463.4]
  assign _T_172 = io_rst == 1'h0; // @[Controllers.scala 131:45:@466.4]
  assign _T_175 = ~ iterDone_1_io_output; // @[Controllers.scala 135:80:@470.4]
  assign _T_176 = iterDone_0_io_output & _T_175; // @[Controllers.scala 135:78:@471.4]
  assign _T_178 = io_doneIn_1 == 1'h0; // @[Controllers.scala 135:105:@472.4]
  assign _T_179 = _T_176 & _T_178; // @[Controllers.scala 135:103:@473.4]
  assign _T_180 = _T_179 & io_enable; // @[Controllers.scala 135:119:@474.4]
  assign _T_182 = io_doneIn_0 | _T_180; // @[Controllers.scala 135:51:@476.4]
  assign _T_205 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@501.4]
  assign _T_207 = _T_205 & _T_150; // @[Controllers.scala 213:90:@503.4]
  assign _T_209 = ~ allDone; // @[Controllers.scala 213:132:@505.4]
  assign _T_210 = _T_207 & _T_209; // @[Controllers.scala 213:130:@506.4]
  assign _T_211 = ~ io_ctrDone; // @[Controllers.scala 213:156:@507.4]
  assign _T_213 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@510.4]
  assign _T_215 = _T_213 & _T_175; // @[Controllers.scala 213:90:@512.4]
  assign _T_222 = allDone == 1'h0; // @[package.scala 100:49:@518.4]
  assign io_done = RetimeWrapper_2_io_out; // @[Controllers.scala 245:13:@547.4]
  assign io_ctrInc = io_doneIn_1; // @[Controllers.scala 122:17:@426.4]
  assign io_enableOut_0 = _T_210 & _T_211; // @[Controllers.scala 213:55:@509.4]
  assign io_enableOut_1 = _T_215 & _T_209; // @[Controllers.scala 213:55:@517.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@498.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@500.4]
  assign active_0_clock = clock; // @[:@358.4]
  assign active_0_reset = reset; // @[:@359.4]
  assign active_0_io_input_set = _T_151 & _T_153; // @[Controllers.scala 128:30:@450.4]
  assign active_0_io_input_reset = _T_155 | allDone; // @[Controllers.scala 129:32:@455.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@372.4]
  assign active_1_clock = clock; // @[:@361.4]
  assign active_1_reset = reset; // @[:@362.4]
  assign active_1_io_input_set = _T_182 & _T_160; // @[Controllers.scala 135:32:@479.4]
  assign active_1_io_input_reset = io_doneIn_1 | io_rst; // @[Controllers.scala 136:34:@483.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@373.4]
  assign done_0_clock = clock; // @[:@364.4]
  assign done_0_reset = reset; // @[:@365.4]
  assign done_0_io_input_set = io_ctrDone & _T_172; // @[Controllers.scala 131:28:@469.4]
  assign done_0_io_input_reset = io_rst | allDone; // @[Controllers.scala 86:33:@384.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@374.4]
  assign done_1_clock = clock; // @[:@367.4]
  assign done_1_reset = reset; // @[:@368.4]
  assign done_1_io_input_set = io_ctrDone & _T_172; // @[Controllers.scala 138:30:@496.4]
  assign done_1_io_input_reset = io_rst | allDone; // @[Controllers.scala 86:33:@393.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@375.4]
  assign iterDone_0_clock = clock; // @[:@396.4]
  assign iterDone_0_reset = reset; // @[:@397.4]
  assign iterDone_0_io_input_set = _T_161 & _T_169; // @[Controllers.scala 130:32:@465.4]
  assign iterDone_0_io_input_reset = synchronize | io_rst; // @[Controllers.scala 92:37:@411.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@401.4]
  assign iterDone_1_clock = clock; // @[:@399.4]
  assign iterDone_1_reset = reset; // @[:@400.4]
  assign iterDone_1_io_input_set = io_doneIn_1 & _T_160; // @[Controllers.scala 137:34:@492.4]
  assign iterDone_1_io_input_reset = synchronize | io_rst; // @[Controllers.scala 92:37:@420.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@402.4]
  assign RetimeWrapper_clock = clock; // @[:@428.4]
  assign RetimeWrapper_reset = reset; // @[:@429.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@431.4]
  assign RetimeWrapper_io_in = io_doneIn_1; // @[package.scala 94:16:@430.4]
  assign RetimeWrapper_1_clock = clock; // @[:@524.4]
  assign RetimeWrapper_1_reset = reset; // @[:@525.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@527.4]
  assign RetimeWrapper_1_io_in = allDone & _T_225; // @[package.scala 94:16:@526.4]
  assign RetimeWrapper_2_clock = clock; // @[:@541.4]
  assign RetimeWrapper_2_reset = reset; // @[:@542.4]
  assign RetimeWrapper_2_io_flow = io_enable; // @[package.scala 95:18:@544.4]
  assign RetimeWrapper_2_io_in = allDone & _T_239; // @[package.scala 94:16:@543.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_225 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_239 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_225 <= 1'h0;
    end else begin
      _T_225 <= _T_222;
    end
    if (reset) begin
      _T_239 <= 1'h0;
    end else begin
      _T_239 <= _T_222;
    end
  end
endmodule
module SRAM( // @[:@613.2]
  input         clock, // @[:@614.4]
  input         reset, // @[:@615.4]
  input  [1:0]  io_raddr, // @[:@616.4]
  input         io_wen, // @[:@616.4]
  input  [1:0]  io_waddr, // @[:@616.4]
  input  [63:0] io_wdata, // @[:@616.4]
  output [63:0] io_rdata, // @[:@616.4]
  input         io_backpressure // @[:@616.4]
);
  wire [63:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 124:30:@618.4]
  wire [63:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 124:30:@618.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 124:30:@618.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 124:30:@618.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 124:30:@618.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 124:30:@618.4]
  wire [1:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 124:30:@618.4]
  wire [1:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 124:30:@618.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 124:30:@618.4]
  wire  _T_19; // @[SRAM.scala 137:49:@636.4]
  wire  _T_20; // @[SRAM.scala 137:37:@637.4]
  reg  _T_23; // @[SRAM.scala 137:29:@638.4]
  reg [31:0] _RAND_0;
  reg [63:0] _T_26; // @[SRAM.scala 138:29:@640.4]
  reg [63:0] _RAND_1;
  SRAMVerilogAWS #(.DWIDTH(64), .WORDS(4), .AWIDTH(2)) SRAMVerilogAWS ( // @[SRAM.scala 124:30:@618.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_19 = io_raddr == io_waddr; // @[SRAM.scala 137:49:@636.4]
  assign _T_20 = io_wen & _T_19; // @[SRAM.scala 137:37:@637.4]
  assign io_rdata = _T_23 ? _T_26 : SRAMVerilogAWS_rdata; // @[SRAM.scala 139:16:@645.4]
  assign SRAMVerilogAWS_wdata = io_wdata; // @[SRAM.scala 130:20:@632.4]
  assign SRAMVerilogAWS_backpressure = io_backpressure; // @[SRAM.scala 131:27:@633.4]
  assign SRAMVerilogAWS_wen = io_wen; // @[SRAM.scala 128:18:@630.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 133:22:@635.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 132:22:@634.4]
  assign SRAMVerilogAWS_waddr = io_waddr; // @[SRAM.scala 129:20:@631.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 127:20:@629.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 126:18:@628.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_23 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {2{`RANDOM}};
  _T_26 = _RAND_1[63:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_23 <= 1'h0;
    end else begin
      _T_23 <= _T_20;
    end
    if (reset) begin
      _T_26 <= 64'h0;
    end else begin
      _T_26 <= io_wdata;
    end
  end
endmodule
module RetimeWrapper_5( // @[:@659.2]
  input        clock, // @[:@660.4]
  input        reset, // @[:@661.4]
  input        io_flow, // @[:@662.4]
  input  [2:0] io_in, // @[:@662.4]
  output [2:0] io_out // @[:@662.4]
);
  wire [2:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@664.4]
  wire [2:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@664.4]
  wire [2:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@664.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@664.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@664.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@664.4]
  RetimeShiftRegister #(.WIDTH(3), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@664.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@677.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@676.4]
  assign sr_init = 3'h0; // @[RetimeShiftRegister.scala 19:16:@675.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@674.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@673.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@671.4]
endmodule
module Mem1D( // @[:@679.2]
  input         clock, // @[:@680.4]
  input         reset, // @[:@681.4]
  input  [2:0]  io_r_ofs_0, // @[:@682.4]
  input         io_r_backpressure, // @[:@682.4]
  input  [2:0]  io_w_ofs_0, // @[:@682.4]
  input  [63:0] io_w_data_0, // @[:@682.4]
  input         io_w_en_0, // @[:@682.4]
  output [63:0] io_output // @[:@682.4]
);
  wire  SRAM_clock; // @[MemPrimitives.scala 567:21:@686.4]
  wire  SRAM_reset; // @[MemPrimitives.scala 567:21:@686.4]
  wire [1:0] SRAM_io_raddr; // @[MemPrimitives.scala 567:21:@686.4]
  wire  SRAM_io_wen; // @[MemPrimitives.scala 567:21:@686.4]
  wire [1:0] SRAM_io_waddr; // @[MemPrimitives.scala 567:21:@686.4]
  wire [63:0] SRAM_io_wdata; // @[MemPrimitives.scala 567:21:@686.4]
  wire [63:0] SRAM_io_rdata; // @[MemPrimitives.scala 567:21:@686.4]
  wire  SRAM_io_backpressure; // @[MemPrimitives.scala 567:21:@686.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@689.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@689.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@689.4]
  wire [2:0] RetimeWrapper_io_in; // @[package.scala 93:22:@689.4]
  wire [2:0] RetimeWrapper_io_out; // @[package.scala 93:22:@689.4]
  wire  wInBound; // @[MemPrimitives.scala 554:32:@684.4]
  wire [2:0] _T_126; // @[package.scala 96:25:@694.4 package.scala 96:25:@695.4]
  SRAM SRAM ( // @[MemPrimitives.scala 567:21:@686.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata(SRAM_io_wdata),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  RetimeWrapper_5 RetimeWrapper ( // @[package.scala 93:22:@689.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign wInBound = io_w_ofs_0 <= 3'h4; // @[MemPrimitives.scala 554:32:@684.4]
  assign _T_126 = RetimeWrapper_io_out; // @[package.scala 96:25:@694.4 package.scala 96:25:@695.4]
  assign io_output = SRAM_io_rdata; // @[MemPrimitives.scala 574:17:@702.4]
  assign SRAM_clock = clock; // @[:@687.4]
  assign SRAM_reset = reset; // @[:@688.4]
  assign SRAM_io_raddr = _T_126[1:0]; // @[MemPrimitives.scala 568:37:@696.4]
  assign SRAM_io_wen = io_w_en_0 & wInBound; // @[MemPrimitives.scala 571:22:@699.4]
  assign SRAM_io_waddr = io_w_ofs_0[1:0]; // @[MemPrimitives.scala 570:22:@697.4]
  assign SRAM_io_wdata = io_w_data_0; // @[MemPrimitives.scala 572:22:@700.4]
  assign SRAM_io_backpressure = io_r_backpressure; // @[MemPrimitives.scala 573:30:@701.4]
  assign RetimeWrapper_clock = clock; // @[:@690.4]
  assign RetimeWrapper_reset = reset; // @[:@691.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@693.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@692.4]
endmodule
module StickySelects( // @[:@1453.2]
  input   io_ins_0, // @[:@1456.4]
  output  io_outs_0 // @[:@1456.4]
);
  assign io_outs_0 = io_ins_0; // @[StickySelects.scala 12:26:@1458.4]
endmodule
module RetimeWrapper_13( // @[:@1521.2]
  input   clock, // @[:@1522.4]
  input   reset, // @[:@1523.4]
  input   io_in, // @[:@1524.4]
  output  io_out // @[:@1524.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@1526.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@1526.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@1526.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@1526.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@1526.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@1526.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@1526.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@1539.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@1538.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@1537.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@1536.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@1535.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@1533.4]
endmodule
module x452_a_0( // @[:@1765.2]
  input         clock, // @[:@1766.4]
  input         reset, // @[:@1767.4]
  input         io_rPort_7_en_0, // @[:@1768.4]
  output [63:0] io_rPort_7_output_0, // @[:@1768.4]
  input         io_rPort_6_en_0, // @[:@1768.4]
  output [63:0] io_rPort_6_output_0, // @[:@1768.4]
  input         io_rPort_5_en_0, // @[:@1768.4]
  output [63:0] io_rPort_5_output_0, // @[:@1768.4]
  input         io_rPort_4_en_0, // @[:@1768.4]
  output [63:0] io_rPort_4_output_0, // @[:@1768.4]
  input         io_rPort_3_en_0, // @[:@1768.4]
  output [63:0] io_rPort_3_output_0, // @[:@1768.4]
  input         io_rPort_2_en_0, // @[:@1768.4]
  output [63:0] io_rPort_2_output_0, // @[:@1768.4]
  input         io_rPort_1_en_0, // @[:@1768.4]
  output [63:0] io_rPort_1_output_0, // @[:@1768.4]
  input         io_rPort_0_en_0, // @[:@1768.4]
  output [63:0] io_rPort_0_output_0, // @[:@1768.4]
  input  [3:0]  io_wPort_0_banks_0, // @[:@1768.4]
  input  [2:0]  io_wPort_0_ofs_0, // @[:@1768.4]
  input  [63:0] io_wPort_0_data_0, // @[:@1768.4]
  input         io_wPort_0_en_0 // @[:@1768.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@1818.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@1818.4]
  wire [2:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@1818.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@1818.4]
  wire [2:0] Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@1818.4]
  wire [63:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@1818.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@1818.4]
  wire [63:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@1818.4]
  wire  Mem1D_1_clock; // @[MemPrimitives.scala 64:21:@1834.4]
  wire  Mem1D_1_reset; // @[MemPrimitives.scala 64:21:@1834.4]
  wire [2:0] Mem1D_1_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@1834.4]
  wire  Mem1D_1_io_r_backpressure; // @[MemPrimitives.scala 64:21:@1834.4]
  wire [2:0] Mem1D_1_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@1834.4]
  wire [63:0] Mem1D_1_io_w_data_0; // @[MemPrimitives.scala 64:21:@1834.4]
  wire  Mem1D_1_io_w_en_0; // @[MemPrimitives.scala 64:21:@1834.4]
  wire [63:0] Mem1D_1_io_output; // @[MemPrimitives.scala 64:21:@1834.4]
  wire  Mem1D_2_clock; // @[MemPrimitives.scala 64:21:@1850.4]
  wire  Mem1D_2_reset; // @[MemPrimitives.scala 64:21:@1850.4]
  wire [2:0] Mem1D_2_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@1850.4]
  wire  Mem1D_2_io_r_backpressure; // @[MemPrimitives.scala 64:21:@1850.4]
  wire [2:0] Mem1D_2_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@1850.4]
  wire [63:0] Mem1D_2_io_w_data_0; // @[MemPrimitives.scala 64:21:@1850.4]
  wire  Mem1D_2_io_w_en_0; // @[MemPrimitives.scala 64:21:@1850.4]
  wire [63:0] Mem1D_2_io_output; // @[MemPrimitives.scala 64:21:@1850.4]
  wire  Mem1D_3_clock; // @[MemPrimitives.scala 64:21:@1866.4]
  wire  Mem1D_3_reset; // @[MemPrimitives.scala 64:21:@1866.4]
  wire [2:0] Mem1D_3_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@1866.4]
  wire  Mem1D_3_io_r_backpressure; // @[MemPrimitives.scala 64:21:@1866.4]
  wire [2:0] Mem1D_3_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@1866.4]
  wire [63:0] Mem1D_3_io_w_data_0; // @[MemPrimitives.scala 64:21:@1866.4]
  wire  Mem1D_3_io_w_en_0; // @[MemPrimitives.scala 64:21:@1866.4]
  wire [63:0] Mem1D_3_io_output; // @[MemPrimitives.scala 64:21:@1866.4]
  wire  Mem1D_4_clock; // @[MemPrimitives.scala 64:21:@1882.4]
  wire  Mem1D_4_reset; // @[MemPrimitives.scala 64:21:@1882.4]
  wire [2:0] Mem1D_4_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@1882.4]
  wire  Mem1D_4_io_r_backpressure; // @[MemPrimitives.scala 64:21:@1882.4]
  wire [2:0] Mem1D_4_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@1882.4]
  wire [63:0] Mem1D_4_io_w_data_0; // @[MemPrimitives.scala 64:21:@1882.4]
  wire  Mem1D_4_io_w_en_0; // @[MemPrimitives.scala 64:21:@1882.4]
  wire [63:0] Mem1D_4_io_output; // @[MemPrimitives.scala 64:21:@1882.4]
  wire  Mem1D_5_clock; // @[MemPrimitives.scala 64:21:@1898.4]
  wire  Mem1D_5_reset; // @[MemPrimitives.scala 64:21:@1898.4]
  wire [2:0] Mem1D_5_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@1898.4]
  wire  Mem1D_5_io_r_backpressure; // @[MemPrimitives.scala 64:21:@1898.4]
  wire [2:0] Mem1D_5_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@1898.4]
  wire [63:0] Mem1D_5_io_w_data_0; // @[MemPrimitives.scala 64:21:@1898.4]
  wire  Mem1D_5_io_w_en_0; // @[MemPrimitives.scala 64:21:@1898.4]
  wire [63:0] Mem1D_5_io_output; // @[MemPrimitives.scala 64:21:@1898.4]
  wire  Mem1D_6_clock; // @[MemPrimitives.scala 64:21:@1914.4]
  wire  Mem1D_6_reset; // @[MemPrimitives.scala 64:21:@1914.4]
  wire [2:0] Mem1D_6_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@1914.4]
  wire  Mem1D_6_io_r_backpressure; // @[MemPrimitives.scala 64:21:@1914.4]
  wire [2:0] Mem1D_6_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@1914.4]
  wire [63:0] Mem1D_6_io_w_data_0; // @[MemPrimitives.scala 64:21:@1914.4]
  wire  Mem1D_6_io_w_en_0; // @[MemPrimitives.scala 64:21:@1914.4]
  wire [63:0] Mem1D_6_io_output; // @[MemPrimitives.scala 64:21:@1914.4]
  wire  Mem1D_7_clock; // @[MemPrimitives.scala 64:21:@1930.4]
  wire  Mem1D_7_reset; // @[MemPrimitives.scala 64:21:@1930.4]
  wire [2:0] Mem1D_7_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@1930.4]
  wire  Mem1D_7_io_r_backpressure; // @[MemPrimitives.scala 64:21:@1930.4]
  wire [2:0] Mem1D_7_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@1930.4]
  wire [63:0] Mem1D_7_io_w_data_0; // @[MemPrimitives.scala 64:21:@1930.4]
  wire  Mem1D_7_io_w_en_0; // @[MemPrimitives.scala 64:21:@1930.4]
  wire [63:0] Mem1D_7_io_output; // @[MemPrimitives.scala 64:21:@1930.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 121:29:@2027.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 121:29:@2027.4]
  wire  StickySelects_1_io_ins_0; // @[MemPrimitives.scala 121:29:@2041.4]
  wire  StickySelects_1_io_outs_0; // @[MemPrimitives.scala 121:29:@2041.4]
  wire  StickySelects_2_io_ins_0; // @[MemPrimitives.scala 121:29:@2055.4]
  wire  StickySelects_2_io_outs_0; // @[MemPrimitives.scala 121:29:@2055.4]
  wire  StickySelects_3_io_ins_0; // @[MemPrimitives.scala 121:29:@2069.4]
  wire  StickySelects_3_io_outs_0; // @[MemPrimitives.scala 121:29:@2069.4]
  wire  StickySelects_4_io_ins_0; // @[MemPrimitives.scala 121:29:@2083.4]
  wire  StickySelects_4_io_outs_0; // @[MemPrimitives.scala 121:29:@2083.4]
  wire  StickySelects_5_io_ins_0; // @[MemPrimitives.scala 121:29:@2097.4]
  wire  StickySelects_5_io_outs_0; // @[MemPrimitives.scala 121:29:@2097.4]
  wire  StickySelects_6_io_ins_0; // @[MemPrimitives.scala 121:29:@2111.4]
  wire  StickySelects_6_io_outs_0; // @[MemPrimitives.scala 121:29:@2111.4]
  wire  StickySelects_7_io_ins_0; // @[MemPrimitives.scala 121:29:@2125.4]
  wire  StickySelects_7_io_outs_0; // @[MemPrimitives.scala 121:29:@2125.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@2139.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@2139.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@2139.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@2139.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@2148.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@2148.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@2148.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@2148.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@2157.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@2157.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@2157.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@2157.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@2166.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@2166.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@2166.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@2166.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@2175.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@2175.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@2175.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@2175.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@2184.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@2184.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@2184.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@2184.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@2193.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@2193.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@2193.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@2193.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@2202.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@2202.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@2202.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@2202.4]
  wire  _T_250; // @[MemPrimitives.scala 82:210:@1946.4]
  wire  _T_251; // @[MemPrimitives.scala 83:102:@1947.4]
  wire [67:0] _T_253; // @[Cat.scala 30:58:@1949.4]
  wire  _T_258; // @[MemPrimitives.scala 82:210:@1956.4]
  wire  _T_259; // @[MemPrimitives.scala 83:102:@1957.4]
  wire [67:0] _T_261; // @[Cat.scala 30:58:@1959.4]
  wire  _T_266; // @[MemPrimitives.scala 82:210:@1966.4]
  wire  _T_267; // @[MemPrimitives.scala 83:102:@1967.4]
  wire [67:0] _T_269; // @[Cat.scala 30:58:@1969.4]
  wire  _T_274; // @[MemPrimitives.scala 82:210:@1976.4]
  wire  _T_275; // @[MemPrimitives.scala 83:102:@1977.4]
  wire [67:0] _T_277; // @[Cat.scala 30:58:@1979.4]
  wire  _T_282; // @[MemPrimitives.scala 82:210:@1986.4]
  wire  _T_283; // @[MemPrimitives.scala 83:102:@1987.4]
  wire [67:0] _T_285; // @[Cat.scala 30:58:@1989.4]
  wire  _T_290; // @[MemPrimitives.scala 82:210:@1996.4]
  wire  _T_291; // @[MemPrimitives.scala 83:102:@1997.4]
  wire [67:0] _T_293; // @[Cat.scala 30:58:@1999.4]
  wire  _T_298; // @[MemPrimitives.scala 82:210:@2006.4]
  wire  _T_299; // @[MemPrimitives.scala 83:102:@2007.4]
  wire [67:0] _T_301; // @[Cat.scala 30:58:@2009.4]
  wire  _T_306; // @[MemPrimitives.scala 82:210:@2016.4]
  wire  _T_307; // @[MemPrimitives.scala 83:102:@2017.4]
  wire [67:0] _T_309; // @[Cat.scala 30:58:@2019.4]
  wire  _T_315; // @[MemPrimitives.scala 123:41:@2031.4]
  wire [4:0] _T_317; // @[Cat.scala 30:58:@2033.4]
  wire  _T_323; // @[MemPrimitives.scala 123:41:@2045.4]
  wire [4:0] _T_325; // @[Cat.scala 30:58:@2047.4]
  wire  _T_331; // @[MemPrimitives.scala 123:41:@2059.4]
  wire [4:0] _T_333; // @[Cat.scala 30:58:@2061.4]
  wire  _T_339; // @[MemPrimitives.scala 123:41:@2073.4]
  wire [4:0] _T_341; // @[Cat.scala 30:58:@2075.4]
  wire  _T_347; // @[MemPrimitives.scala 123:41:@2087.4]
  wire [4:0] _T_349; // @[Cat.scala 30:58:@2089.4]
  wire  _T_355; // @[MemPrimitives.scala 123:41:@2101.4]
  wire [4:0] _T_357; // @[Cat.scala 30:58:@2103.4]
  wire  _T_363; // @[MemPrimitives.scala 123:41:@2115.4]
  wire [4:0] _T_365; // @[Cat.scala 30:58:@2117.4]
  wire  _T_371; // @[MemPrimitives.scala 123:41:@2129.4]
  wire [4:0] _T_373; // @[Cat.scala 30:58:@2131.4]
  Mem1D Mem1D ( // @[MemPrimitives.scala 64:21:@1818.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  Mem1D Mem1D_1 ( // @[MemPrimitives.scala 64:21:@1834.4]
    .clock(Mem1D_1_clock),
    .reset(Mem1D_1_reset),
    .io_r_ofs_0(Mem1D_1_io_r_ofs_0),
    .io_r_backpressure(Mem1D_1_io_r_backpressure),
    .io_w_ofs_0(Mem1D_1_io_w_ofs_0),
    .io_w_data_0(Mem1D_1_io_w_data_0),
    .io_w_en_0(Mem1D_1_io_w_en_0),
    .io_output(Mem1D_1_io_output)
  );
  Mem1D Mem1D_2 ( // @[MemPrimitives.scala 64:21:@1850.4]
    .clock(Mem1D_2_clock),
    .reset(Mem1D_2_reset),
    .io_r_ofs_0(Mem1D_2_io_r_ofs_0),
    .io_r_backpressure(Mem1D_2_io_r_backpressure),
    .io_w_ofs_0(Mem1D_2_io_w_ofs_0),
    .io_w_data_0(Mem1D_2_io_w_data_0),
    .io_w_en_0(Mem1D_2_io_w_en_0),
    .io_output(Mem1D_2_io_output)
  );
  Mem1D Mem1D_3 ( // @[MemPrimitives.scala 64:21:@1866.4]
    .clock(Mem1D_3_clock),
    .reset(Mem1D_3_reset),
    .io_r_ofs_0(Mem1D_3_io_r_ofs_0),
    .io_r_backpressure(Mem1D_3_io_r_backpressure),
    .io_w_ofs_0(Mem1D_3_io_w_ofs_0),
    .io_w_data_0(Mem1D_3_io_w_data_0),
    .io_w_en_0(Mem1D_3_io_w_en_0),
    .io_output(Mem1D_3_io_output)
  );
  Mem1D Mem1D_4 ( // @[MemPrimitives.scala 64:21:@1882.4]
    .clock(Mem1D_4_clock),
    .reset(Mem1D_4_reset),
    .io_r_ofs_0(Mem1D_4_io_r_ofs_0),
    .io_r_backpressure(Mem1D_4_io_r_backpressure),
    .io_w_ofs_0(Mem1D_4_io_w_ofs_0),
    .io_w_data_0(Mem1D_4_io_w_data_0),
    .io_w_en_0(Mem1D_4_io_w_en_0),
    .io_output(Mem1D_4_io_output)
  );
  Mem1D Mem1D_5 ( // @[MemPrimitives.scala 64:21:@1898.4]
    .clock(Mem1D_5_clock),
    .reset(Mem1D_5_reset),
    .io_r_ofs_0(Mem1D_5_io_r_ofs_0),
    .io_r_backpressure(Mem1D_5_io_r_backpressure),
    .io_w_ofs_0(Mem1D_5_io_w_ofs_0),
    .io_w_data_0(Mem1D_5_io_w_data_0),
    .io_w_en_0(Mem1D_5_io_w_en_0),
    .io_output(Mem1D_5_io_output)
  );
  Mem1D Mem1D_6 ( // @[MemPrimitives.scala 64:21:@1914.4]
    .clock(Mem1D_6_clock),
    .reset(Mem1D_6_reset),
    .io_r_ofs_0(Mem1D_6_io_r_ofs_0),
    .io_r_backpressure(Mem1D_6_io_r_backpressure),
    .io_w_ofs_0(Mem1D_6_io_w_ofs_0),
    .io_w_data_0(Mem1D_6_io_w_data_0),
    .io_w_en_0(Mem1D_6_io_w_en_0),
    .io_output(Mem1D_6_io_output)
  );
  Mem1D Mem1D_7 ( // @[MemPrimitives.scala 64:21:@1930.4]
    .clock(Mem1D_7_clock),
    .reset(Mem1D_7_reset),
    .io_r_ofs_0(Mem1D_7_io_r_ofs_0),
    .io_r_backpressure(Mem1D_7_io_r_backpressure),
    .io_w_ofs_0(Mem1D_7_io_w_ofs_0),
    .io_w_data_0(Mem1D_7_io_w_data_0),
    .io_w_en_0(Mem1D_7_io_w_en_0),
    .io_output(Mem1D_7_io_output)
  );
  StickySelects StickySelects ( // @[MemPrimitives.scala 121:29:@2027.4]
    .io_ins_0(StickySelects_io_ins_0),
    .io_outs_0(StickySelects_io_outs_0)
  );
  StickySelects StickySelects_1 ( // @[MemPrimitives.scala 121:29:@2041.4]
    .io_ins_0(StickySelects_1_io_ins_0),
    .io_outs_0(StickySelects_1_io_outs_0)
  );
  StickySelects StickySelects_2 ( // @[MemPrimitives.scala 121:29:@2055.4]
    .io_ins_0(StickySelects_2_io_ins_0),
    .io_outs_0(StickySelects_2_io_outs_0)
  );
  StickySelects StickySelects_3 ( // @[MemPrimitives.scala 121:29:@2069.4]
    .io_ins_0(StickySelects_3_io_ins_0),
    .io_outs_0(StickySelects_3_io_outs_0)
  );
  StickySelects StickySelects_4 ( // @[MemPrimitives.scala 121:29:@2083.4]
    .io_ins_0(StickySelects_4_io_ins_0),
    .io_outs_0(StickySelects_4_io_outs_0)
  );
  StickySelects StickySelects_5 ( // @[MemPrimitives.scala 121:29:@2097.4]
    .io_ins_0(StickySelects_5_io_ins_0),
    .io_outs_0(StickySelects_5_io_outs_0)
  );
  StickySelects StickySelects_6 ( // @[MemPrimitives.scala 121:29:@2111.4]
    .io_ins_0(StickySelects_6_io_ins_0),
    .io_outs_0(StickySelects_6_io_outs_0)
  );
  StickySelects StickySelects_7 ( // @[MemPrimitives.scala 121:29:@2125.4]
    .io_ins_0(StickySelects_7_io_ins_0),
    .io_outs_0(StickySelects_7_io_outs_0)
  );
  RetimeWrapper_13 RetimeWrapper ( // @[package.scala 93:22:@2139.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_13 RetimeWrapper_1 ( // @[package.scala 93:22:@2148.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_13 RetimeWrapper_2 ( // @[package.scala 93:22:@2157.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_13 RetimeWrapper_3 ( // @[package.scala 93:22:@2166.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_13 RetimeWrapper_4 ( // @[package.scala 93:22:@2175.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_13 RetimeWrapper_5 ( // @[package.scala 93:22:@2184.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_13 RetimeWrapper_6 ( // @[package.scala 93:22:@2193.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_13 RetimeWrapper_7 ( // @[package.scala 93:22:@2202.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  assign _T_250 = io_wPort_0_banks_0 == 4'h0; // @[MemPrimitives.scala 82:210:@1946.4]
  assign _T_251 = io_wPort_0_en_0 & _T_250; // @[MemPrimitives.scala 83:102:@1947.4]
  assign _T_253 = {_T_251,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@1949.4]
  assign _T_258 = io_wPort_0_banks_0 == 4'h1; // @[MemPrimitives.scala 82:210:@1956.4]
  assign _T_259 = io_wPort_0_en_0 & _T_258; // @[MemPrimitives.scala 83:102:@1957.4]
  assign _T_261 = {_T_259,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@1959.4]
  assign _T_266 = io_wPort_0_banks_0 == 4'h2; // @[MemPrimitives.scala 82:210:@1966.4]
  assign _T_267 = io_wPort_0_en_0 & _T_266; // @[MemPrimitives.scala 83:102:@1967.4]
  assign _T_269 = {_T_267,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@1969.4]
  assign _T_274 = io_wPort_0_banks_0 == 4'h3; // @[MemPrimitives.scala 82:210:@1976.4]
  assign _T_275 = io_wPort_0_en_0 & _T_274; // @[MemPrimitives.scala 83:102:@1977.4]
  assign _T_277 = {_T_275,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@1979.4]
  assign _T_282 = io_wPort_0_banks_0 == 4'h4; // @[MemPrimitives.scala 82:210:@1986.4]
  assign _T_283 = io_wPort_0_en_0 & _T_282; // @[MemPrimitives.scala 83:102:@1987.4]
  assign _T_285 = {_T_283,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@1989.4]
  assign _T_290 = io_wPort_0_banks_0 == 4'h5; // @[MemPrimitives.scala 82:210:@1996.4]
  assign _T_291 = io_wPort_0_en_0 & _T_290; // @[MemPrimitives.scala 83:102:@1997.4]
  assign _T_293 = {_T_291,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@1999.4]
  assign _T_298 = io_wPort_0_banks_0 == 4'h6; // @[MemPrimitives.scala 82:210:@2006.4]
  assign _T_299 = io_wPort_0_en_0 & _T_298; // @[MemPrimitives.scala 83:102:@2007.4]
  assign _T_301 = {_T_299,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@2009.4]
  assign _T_306 = io_wPort_0_banks_0 == 4'h7; // @[MemPrimitives.scala 82:210:@2016.4]
  assign _T_307 = io_wPort_0_en_0 & _T_306; // @[MemPrimitives.scala 83:102:@2017.4]
  assign _T_309 = {_T_307,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@2019.4]
  assign _T_315 = StickySelects_io_outs_0; // @[MemPrimitives.scala 123:41:@2031.4]
  assign _T_317 = {_T_315,1'h1,3'h0}; // @[Cat.scala 30:58:@2033.4]
  assign _T_323 = StickySelects_1_io_outs_0; // @[MemPrimitives.scala 123:41:@2045.4]
  assign _T_325 = {_T_323,1'h1,3'h0}; // @[Cat.scala 30:58:@2047.4]
  assign _T_331 = StickySelects_2_io_outs_0; // @[MemPrimitives.scala 123:41:@2059.4]
  assign _T_333 = {_T_331,1'h1,3'h0}; // @[Cat.scala 30:58:@2061.4]
  assign _T_339 = StickySelects_3_io_outs_0; // @[MemPrimitives.scala 123:41:@2073.4]
  assign _T_341 = {_T_339,1'h1,3'h0}; // @[Cat.scala 30:58:@2075.4]
  assign _T_347 = StickySelects_4_io_outs_0; // @[MemPrimitives.scala 123:41:@2087.4]
  assign _T_349 = {_T_347,1'h1,3'h0}; // @[Cat.scala 30:58:@2089.4]
  assign _T_355 = StickySelects_5_io_outs_0; // @[MemPrimitives.scala 123:41:@2101.4]
  assign _T_357 = {_T_355,1'h1,3'h0}; // @[Cat.scala 30:58:@2103.4]
  assign _T_363 = StickySelects_6_io_outs_0; // @[MemPrimitives.scala 123:41:@2115.4]
  assign _T_365 = {_T_363,1'h1,3'h0}; // @[Cat.scala 30:58:@2117.4]
  assign _T_371 = StickySelects_7_io_outs_0; // @[MemPrimitives.scala 123:41:@2129.4]
  assign _T_373 = {_T_371,1'h1,3'h0}; // @[Cat.scala 30:58:@2131.4]
  assign io_rPort_7_output_0 = Mem1D_1_io_output; // @[MemPrimitives.scala 148:13:@2209.4]
  assign io_rPort_6_output_0 = Mem1D_7_io_output; // @[MemPrimitives.scala 148:13:@2200.4]
  assign io_rPort_5_output_0 = Mem1D_2_io_output; // @[MemPrimitives.scala 148:13:@2191.4]
  assign io_rPort_4_output_0 = Mem1D_5_io_output; // @[MemPrimitives.scala 148:13:@2182.4]
  assign io_rPort_3_output_0 = Mem1D_io_output; // @[MemPrimitives.scala 148:13:@2173.4]
  assign io_rPort_2_output_0 = Mem1D_3_io_output; // @[MemPrimitives.scala 148:13:@2164.4]
  assign io_rPort_1_output_0 = Mem1D_6_io_output; // @[MemPrimitives.scala 148:13:@2155.4]
  assign io_rPort_0_output_0 = Mem1D_4_io_output; // @[MemPrimitives.scala 148:13:@2146.4]
  assign Mem1D_clock = clock; // @[:@1819.4]
  assign Mem1D_reset = reset; // @[:@1820.4]
  assign Mem1D_io_r_ofs_0 = _T_317[2:0]; // @[MemPrimitives.scala 127:28:@2037.4]
  assign Mem1D_io_r_backpressure = _T_317[3]; // @[MemPrimitives.scala 128:32:@2038.4]
  assign Mem1D_io_w_ofs_0 = _T_253[2:0]; // @[MemPrimitives.scala 94:28:@1953.4]
  assign Mem1D_io_w_data_0 = _T_253[66:3]; // @[MemPrimitives.scala 95:29:@1954.4]
  assign Mem1D_io_w_en_0 = _T_253[67]; // @[MemPrimitives.scala 96:27:@1955.4]
  assign Mem1D_1_clock = clock; // @[:@1835.4]
  assign Mem1D_1_reset = reset; // @[:@1836.4]
  assign Mem1D_1_io_r_ofs_0 = _T_325[2:0]; // @[MemPrimitives.scala 127:28:@2051.4]
  assign Mem1D_1_io_r_backpressure = _T_325[3]; // @[MemPrimitives.scala 128:32:@2052.4]
  assign Mem1D_1_io_w_ofs_0 = _T_261[2:0]; // @[MemPrimitives.scala 94:28:@1963.4]
  assign Mem1D_1_io_w_data_0 = _T_261[66:3]; // @[MemPrimitives.scala 95:29:@1964.4]
  assign Mem1D_1_io_w_en_0 = _T_261[67]; // @[MemPrimitives.scala 96:27:@1965.4]
  assign Mem1D_2_clock = clock; // @[:@1851.4]
  assign Mem1D_2_reset = reset; // @[:@1852.4]
  assign Mem1D_2_io_r_ofs_0 = _T_333[2:0]; // @[MemPrimitives.scala 127:28:@2065.4]
  assign Mem1D_2_io_r_backpressure = _T_333[3]; // @[MemPrimitives.scala 128:32:@2066.4]
  assign Mem1D_2_io_w_ofs_0 = _T_269[2:0]; // @[MemPrimitives.scala 94:28:@1973.4]
  assign Mem1D_2_io_w_data_0 = _T_269[66:3]; // @[MemPrimitives.scala 95:29:@1974.4]
  assign Mem1D_2_io_w_en_0 = _T_269[67]; // @[MemPrimitives.scala 96:27:@1975.4]
  assign Mem1D_3_clock = clock; // @[:@1867.4]
  assign Mem1D_3_reset = reset; // @[:@1868.4]
  assign Mem1D_3_io_r_ofs_0 = _T_341[2:0]; // @[MemPrimitives.scala 127:28:@2079.4]
  assign Mem1D_3_io_r_backpressure = _T_341[3]; // @[MemPrimitives.scala 128:32:@2080.4]
  assign Mem1D_3_io_w_ofs_0 = _T_277[2:0]; // @[MemPrimitives.scala 94:28:@1983.4]
  assign Mem1D_3_io_w_data_0 = _T_277[66:3]; // @[MemPrimitives.scala 95:29:@1984.4]
  assign Mem1D_3_io_w_en_0 = _T_277[67]; // @[MemPrimitives.scala 96:27:@1985.4]
  assign Mem1D_4_clock = clock; // @[:@1883.4]
  assign Mem1D_4_reset = reset; // @[:@1884.4]
  assign Mem1D_4_io_r_ofs_0 = _T_349[2:0]; // @[MemPrimitives.scala 127:28:@2093.4]
  assign Mem1D_4_io_r_backpressure = _T_349[3]; // @[MemPrimitives.scala 128:32:@2094.4]
  assign Mem1D_4_io_w_ofs_0 = _T_285[2:0]; // @[MemPrimitives.scala 94:28:@1993.4]
  assign Mem1D_4_io_w_data_0 = _T_285[66:3]; // @[MemPrimitives.scala 95:29:@1994.4]
  assign Mem1D_4_io_w_en_0 = _T_285[67]; // @[MemPrimitives.scala 96:27:@1995.4]
  assign Mem1D_5_clock = clock; // @[:@1899.4]
  assign Mem1D_5_reset = reset; // @[:@1900.4]
  assign Mem1D_5_io_r_ofs_0 = _T_357[2:0]; // @[MemPrimitives.scala 127:28:@2107.4]
  assign Mem1D_5_io_r_backpressure = _T_357[3]; // @[MemPrimitives.scala 128:32:@2108.4]
  assign Mem1D_5_io_w_ofs_0 = _T_293[2:0]; // @[MemPrimitives.scala 94:28:@2003.4]
  assign Mem1D_5_io_w_data_0 = _T_293[66:3]; // @[MemPrimitives.scala 95:29:@2004.4]
  assign Mem1D_5_io_w_en_0 = _T_293[67]; // @[MemPrimitives.scala 96:27:@2005.4]
  assign Mem1D_6_clock = clock; // @[:@1915.4]
  assign Mem1D_6_reset = reset; // @[:@1916.4]
  assign Mem1D_6_io_r_ofs_0 = _T_365[2:0]; // @[MemPrimitives.scala 127:28:@2121.4]
  assign Mem1D_6_io_r_backpressure = _T_365[3]; // @[MemPrimitives.scala 128:32:@2122.4]
  assign Mem1D_6_io_w_ofs_0 = _T_301[2:0]; // @[MemPrimitives.scala 94:28:@2013.4]
  assign Mem1D_6_io_w_data_0 = _T_301[66:3]; // @[MemPrimitives.scala 95:29:@2014.4]
  assign Mem1D_6_io_w_en_0 = _T_301[67]; // @[MemPrimitives.scala 96:27:@2015.4]
  assign Mem1D_7_clock = clock; // @[:@1931.4]
  assign Mem1D_7_reset = reset; // @[:@1932.4]
  assign Mem1D_7_io_r_ofs_0 = _T_373[2:0]; // @[MemPrimitives.scala 127:28:@2135.4]
  assign Mem1D_7_io_r_backpressure = _T_373[3]; // @[MemPrimitives.scala 128:32:@2136.4]
  assign Mem1D_7_io_w_ofs_0 = _T_309[2:0]; // @[MemPrimitives.scala 94:28:@2023.4]
  assign Mem1D_7_io_w_data_0 = _T_309[66:3]; // @[MemPrimitives.scala 95:29:@2024.4]
  assign Mem1D_7_io_w_en_0 = _T_309[67]; // @[MemPrimitives.scala 96:27:@2025.4]
  assign StickySelects_io_ins_0 = io_rPort_3_en_0; // @[MemPrimitives.scala 122:60:@2030.4]
  assign StickySelects_1_io_ins_0 = io_rPort_7_en_0; // @[MemPrimitives.scala 122:60:@2044.4]
  assign StickySelects_2_io_ins_0 = io_rPort_5_en_0; // @[MemPrimitives.scala 122:60:@2058.4]
  assign StickySelects_3_io_ins_0 = io_rPort_2_en_0; // @[MemPrimitives.scala 122:60:@2072.4]
  assign StickySelects_4_io_ins_0 = io_rPort_0_en_0; // @[MemPrimitives.scala 122:60:@2086.4]
  assign StickySelects_5_io_ins_0 = io_rPort_4_en_0; // @[MemPrimitives.scala 122:60:@2100.4]
  assign StickySelects_6_io_ins_0 = io_rPort_1_en_0; // @[MemPrimitives.scala 122:60:@2114.4]
  assign StickySelects_7_io_ins_0 = io_rPort_6_en_0; // @[MemPrimitives.scala 122:60:@2128.4]
  assign RetimeWrapper_clock = clock; // @[:@2140.4]
  assign RetimeWrapper_reset = reset; // @[:@2141.4]
  assign RetimeWrapper_io_in = io_rPort_0_en_0; // @[package.scala 94:16:@2142.4]
  assign RetimeWrapper_1_clock = clock; // @[:@2149.4]
  assign RetimeWrapper_1_reset = reset; // @[:@2150.4]
  assign RetimeWrapper_1_io_in = io_rPort_1_en_0; // @[package.scala 94:16:@2151.4]
  assign RetimeWrapper_2_clock = clock; // @[:@2158.4]
  assign RetimeWrapper_2_reset = reset; // @[:@2159.4]
  assign RetimeWrapper_2_io_in = io_rPort_2_en_0; // @[package.scala 94:16:@2160.4]
  assign RetimeWrapper_3_clock = clock; // @[:@2167.4]
  assign RetimeWrapper_3_reset = reset; // @[:@2168.4]
  assign RetimeWrapper_3_io_in = io_rPort_3_en_0; // @[package.scala 94:16:@2169.4]
  assign RetimeWrapper_4_clock = clock; // @[:@2176.4]
  assign RetimeWrapper_4_reset = reset; // @[:@2177.4]
  assign RetimeWrapper_4_io_in = io_rPort_4_en_0; // @[package.scala 94:16:@2178.4]
  assign RetimeWrapper_5_clock = clock; // @[:@2185.4]
  assign RetimeWrapper_5_reset = reset; // @[:@2186.4]
  assign RetimeWrapper_5_io_in = io_rPort_5_en_0; // @[package.scala 94:16:@2187.4]
  assign RetimeWrapper_6_clock = clock; // @[:@2194.4]
  assign RetimeWrapper_6_reset = reset; // @[:@2195.4]
  assign RetimeWrapper_6_io_in = io_rPort_6_en_0; // @[package.scala 94:16:@2196.4]
  assign RetimeWrapper_7_clock = clock; // @[:@2203.4]
  assign RetimeWrapper_7_reset = reset; // @[:@2204.4]
  assign RetimeWrapper_7_io_in = io_rPort_7_en_0; // @[package.scala 94:16:@2205.4]
endmodule
module x466_outr_UnitPipe_sm( // @[:@2410.2]
  input   clock, // @[:@2411.4]
  input   reset, // @[:@2412.4]
  input   io_enable, // @[:@2413.4]
  output  io_done, // @[:@2413.4]
  input   io_parentAck, // @[:@2413.4]
  input   io_doneIn_0, // @[:@2413.4]
  output  io_enableOut_0, // @[:@2413.4]
  output  io_childAck_0, // @[:@2413.4]
  input   io_ctrCopyDone_0 // @[:@2413.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@2416.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@2416.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@2416.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@2416.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@2416.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@2416.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@2419.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@2419.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@2419.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@2419.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@2419.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@2419.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@2436.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@2436.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@2436.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@2436.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@2436.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@2436.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@2467.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@2467.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@2467.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@2467.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@2467.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@2481.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@2481.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@2481.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@2481.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@2481.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@2499.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@2499.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@2499.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@2499.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@2499.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@2536.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@2536.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@2536.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@2536.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@2536.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@2553.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@2553.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@2553.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@2553.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@2553.4]
  wire  _T_105; // @[Controllers.scala 165:35:@2451.4]
  wire  _T_107; // @[Controllers.scala 165:60:@2452.4]
  wire  _T_108; // @[Controllers.scala 165:58:@2453.4]
  wire  _T_110; // @[Controllers.scala 165:76:@2454.4]
  wire  _T_111; // @[Controllers.scala 165:74:@2455.4]
  wire  _T_115; // @[Controllers.scala 165:109:@2458.4]
  wire  _T_118; // @[Controllers.scala 165:141:@2460.4]
  wire  _T_126; // @[package.scala 96:25:@2472.4 package.scala 96:25:@2473.4]
  wire  _T_130; // @[Controllers.scala 167:54:@2475.4]
  wire  _T_131; // @[Controllers.scala 167:52:@2476.4]
  wire  _T_138; // @[package.scala 96:25:@2486.4 package.scala 96:25:@2487.4]
  wire  _T_156; // @[package.scala 96:25:@2504.4 package.scala 96:25:@2505.4]
  wire  _T_160; // @[Controllers.scala 169:67:@2507.4]
  wire  _T_161; // @[Controllers.scala 169:86:@2508.4]
  wire  _T_174; // @[Controllers.scala 213:68:@2522.4]
  wire  _T_176; // @[Controllers.scala 213:90:@2524.4]
  wire  _T_178; // @[Controllers.scala 213:132:@2526.4]
  reg  _T_186; // @[package.scala 48:56:@2532.4]
  reg [31:0] _RAND_0;
  wire  _T_187; // @[package.scala 100:41:@2534.4]
  reg  _T_200; // @[package.scala 48:56:@2550.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@2416.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@2419.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@2436.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@2467.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@2481.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@2499.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@2536.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@2553.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_105 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@2451.4]
  assign _T_107 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@2452.4]
  assign _T_108 = _T_105 & _T_107; // @[Controllers.scala 165:58:@2453.4]
  assign _T_110 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@2454.4]
  assign _T_111 = _T_108 & _T_110; // @[Controllers.scala 165:74:@2455.4]
  assign _T_115 = _T_111 & io_enable; // @[Controllers.scala 165:109:@2458.4]
  assign _T_118 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@2460.4]
  assign _T_126 = RetimeWrapper_io_out; // @[package.scala 96:25:@2472.4 package.scala 96:25:@2473.4]
  assign _T_130 = _T_126 == 1'h0; // @[Controllers.scala 167:54:@2475.4]
  assign _T_131 = io_doneIn_0 | _T_130; // @[Controllers.scala 167:52:@2476.4]
  assign _T_138 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@2486.4 package.scala 96:25:@2487.4]
  assign _T_156 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@2504.4 package.scala 96:25:@2505.4]
  assign _T_160 = _T_156 == 1'h0; // @[Controllers.scala 169:67:@2507.4]
  assign _T_161 = _T_160 & io_enable; // @[Controllers.scala 169:86:@2508.4]
  assign _T_174 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@2522.4]
  assign _T_176 = _T_174 & _T_105; // @[Controllers.scala 213:90:@2524.4]
  assign _T_178 = ~ done_0_io_output; // @[Controllers.scala 213:132:@2526.4]
  assign _T_187 = done_0_io_output & _T_186; // @[package.scala 100:41:@2534.4]
  assign io_done = RetimeWrapper_4_io_out; // @[Controllers.scala 245:13:@2560.4]
  assign io_enableOut_0 = _T_176 & _T_178; // @[Controllers.scala 213:55:@2530.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@2521.4]
  assign active_0_clock = clock; // @[:@2417.4]
  assign active_0_reset = reset; // @[:@2418.4]
  assign active_0_io_input_set = _T_115 & _T_118; // @[Controllers.scala 165:32:@2462.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@2466.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@2424.4]
  assign done_0_clock = clock; // @[:@2420.4]
  assign done_0_reset = reset; // @[:@2421.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_161; // @[Controllers.scala 169:30:@2512.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@2434.4 Controllers.scala 170:32:@2519.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@2425.4]
  assign iterDone_0_clock = clock; // @[:@2437.4]
  assign iterDone_0_reset = reset; // @[:@2438.4]
  assign iterDone_0_io_input_set = _T_131 & io_enable; // @[Controllers.scala 167:34:@2480.4]
  assign iterDone_0_io_input_reset = _T_138 | io_parentAck; // @[Controllers.scala 92:37:@2448.4 Controllers.scala 168:36:@2496.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@2439.4]
  assign RetimeWrapper_clock = clock; // @[:@2468.4]
  assign RetimeWrapper_reset = reset; // @[:@2469.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@2471.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@2470.4]
  assign RetimeWrapper_1_clock = clock; // @[:@2482.4]
  assign RetimeWrapper_1_reset = reset; // @[:@2483.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@2485.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@2484.4]
  assign RetimeWrapper_2_clock = clock; // @[:@2500.4]
  assign RetimeWrapper_2_reset = reset; // @[:@2501.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@2503.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@2502.4]
  assign RetimeWrapper_3_clock = clock; // @[:@2537.4]
  assign RetimeWrapper_3_reset = reset; // @[:@2538.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@2540.4]
  assign RetimeWrapper_3_io_in = _T_187 | io_parentAck; // @[package.scala 94:16:@2539.4]
  assign RetimeWrapper_4_clock = clock; // @[:@2554.4]
  assign RetimeWrapper_4_reset = reset; // @[:@2555.4]
  assign RetimeWrapper_4_io_flow = io_enable; // @[package.scala 95:18:@2557.4]
  assign RetimeWrapper_4_io_in = done_0_io_output & _T_200; // @[package.scala 94:16:@2556.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_186 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_200 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_186 <= 1'h0;
    end else begin
      _T_186 <= _T_110;
    end
    if (reset) begin
      _T_200 <= 1'h0;
    end else begin
      _T_200 <= _T_110;
    end
  end
endmodule
module SingleCounter_1( // @[:@2680.2]
  input         clock, // @[:@2681.4]
  input         reset, // @[:@2682.4]
  input         io_input_reset, // @[:@2683.4]
  input         io_input_enable, // @[:@2683.4]
  output [31:0] io_output_count_0, // @[:@2683.4]
  output        io_output_oobs_0, // @[:@2683.4]
  output        io_output_done // @[:@2683.4]
);
  wire  bases_0_clock; // @[Counter.scala 253:53:@2696.4]
  wire  bases_0_reset; // @[Counter.scala 253:53:@2696.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 253:53:@2696.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 253:53:@2696.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 253:53:@2696.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 253:53:@2696.4]
  wire  SRFF_clock; // @[Counter.scala 255:22:@2712.4]
  wire  SRFF_reset; // @[Counter.scala 255:22:@2712.4]
  wire  SRFF_io_input_set; // @[Counter.scala 255:22:@2712.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 255:22:@2712.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 255:22:@2712.4]
  wire  SRFF_io_output; // @[Counter.scala 255:22:@2712.4]
  wire  _T_36; // @[Counter.scala 256:45:@2715.4]
  wire [31:0] _T_48; // @[Counter.scala 279:52:@2740.4]
  wire [32:0] _T_50; // @[Counter.scala 283:33:@2741.4]
  wire [31:0] _T_51; // @[Counter.scala 283:33:@2742.4]
  wire [31:0] _T_52; // @[Counter.scala 283:33:@2743.4]
  wire  _T_57; // @[Counter.scala 285:18:@2745.4]
  wire [31:0] _T_68; // @[Counter.scala 291:115:@2753.4]
  wire [31:0] _T_71; // @[Counter.scala 291:152:@2756.4]
  wire [31:0] _T_72; // @[Counter.scala 291:74:@2757.4]
  wire  _T_75; // @[Counter.scala 314:102:@2761.4]
  wire  _T_77; // @[Counter.scala 314:130:@2762.4]
  FF bases_0 ( // @[Counter.scala 253:53:@2696.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 255:22:@2712.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 256:45:@2715.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 279:52:@2740.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@2741.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@2742.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 283:33:@2743.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh8); // @[Counter.scala 285:18:@2745.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 291:115:@2753.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 291:152:@2756.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 291:74:@2757.4]
  assign _T_75 = $signed(_T_48) < $signed(32'sh0); // @[Counter.scala 314:102:@2761.4]
  assign _T_77 = $signed(_T_48) >= $signed(32'sh8); // @[Counter.scala 314:130:@2762.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 296:28:@2760.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 314:60:@2764.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 325:20:@2766.4]
  assign bases_0_clock = clock; // @[:@2697.4]
  assign bases_0_reset = reset; // @[:@2698.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 291:31:@2759.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 273:27:@2738.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 276:29:@2739.4]
  assign SRFF_clock = clock; // @[:@2713.4]
  assign SRFF_reset = reset; // @[:@2714.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 256:23:@2717.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 257:25:@2719.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 258:30:@2720.4]
endmodule
module x454_ctrchain( // @[:@2771.2]
  input         clock, // @[:@2772.4]
  input         reset, // @[:@2773.4]
  input         io_input_reset, // @[:@2774.4]
  input         io_input_enable, // @[:@2774.4]
  output [31:0] io_output_counts_0, // @[:@2774.4]
  output        io_output_oobs_0, // @[:@2774.4]
  output        io_output_done // @[:@2774.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 505:46:@2776.4]
  wire  ctrs_0_reset; // @[Counter.scala 505:46:@2776.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 505:46:@2776.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 505:46:@2776.4]
  wire [31:0] ctrs_0_io_output_count_0; // @[Counter.scala 505:46:@2776.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 505:46:@2776.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 505:46:@2776.4]
  reg  wasDone; // @[Counter.scala 534:24:@2785.4]
  reg [31:0] _RAND_0;
  wire  _T_45; // @[Counter.scala 538:69:@2791.4]
  wire  _T_47; // @[Counter.scala 538:80:@2792.4]
  reg  doneLatch; // @[Counter.scala 542:26:@2797.4]
  reg [31:0] _RAND_1;
  wire  _T_54; // @[Counter.scala 543:48:@2798.4]
  wire  _T_55; // @[Counter.scala 543:19:@2799.4]
  SingleCounter_1 ctrs_0 ( // @[Counter.scala 505:46:@2776.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done)
  );
  assign _T_45 = io_input_enable & ctrs_0_io_output_done; // @[Counter.scala 538:69:@2791.4]
  assign _T_47 = wasDone == 1'h0; // @[Counter.scala 538:80:@2792.4]
  assign _T_54 = ctrs_0_io_output_done ? 1'h1 : doneLatch; // @[Counter.scala 543:48:@2798.4]
  assign _T_55 = io_input_reset ? 1'h0 : _T_54; // @[Counter.scala 543:19:@2799.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 549:32:@2801.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 550:30:@2803.4]
  assign io_output_done = _T_45 & _T_47; // @[Counter.scala 538:18:@2794.4]
  assign ctrs_0_clock = clock; // @[:@2777.4]
  assign ctrs_0_reset = reset; // @[:@2778.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 512:24:@2782.4]
  assign ctrs_0_io_input_enable = io_input_enable; // @[Counter.scala 516:33:@2783.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= ctrs_0_io_output_done;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (ctrs_0_io_output_done) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module x465_inr_Foreach_sm( // @[:@2991.2]
  input   clock, // @[:@2992.4]
  input   reset, // @[:@2993.4]
  input   io_enable, // @[:@2994.4]
  output  io_done, // @[:@2994.4]
  output  io_doneLatch, // @[:@2994.4]
  input   io_ctrDone, // @[:@2994.4]
  output  io_datapathEn, // @[:@2994.4]
  output  io_ctrInc, // @[:@2994.4]
  output  io_ctrRst, // @[:@2994.4]
  input   io_parentAck, // @[:@2994.4]
  input   io_break // @[:@2994.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@2996.4]
  wire  active_reset; // @[Controllers.scala 261:22:@2996.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@2996.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@2996.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@2996.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@2996.4]
  wire  done_clock; // @[Controllers.scala 262:20:@2999.4]
  wire  done_reset; // @[Controllers.scala 262:20:@2999.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@2999.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@2999.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@2999.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@2999.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3033.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3033.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@3033.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@3033.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@3055.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@3055.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@3055.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@3055.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@3067.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@3067.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@3067.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@3067.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@3067.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@3075.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@3075.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@3075.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@3075.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@3075.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@3091.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@3091.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@3091.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@3091.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@3091.4]
  wire  _T_80; // @[Controllers.scala 264:48:@3004.4]
  wire  _T_81; // @[Controllers.scala 264:46:@3005.4]
  wire  _T_82; // @[Controllers.scala 264:62:@3006.4]
  wire  _T_100; // @[package.scala 100:49:@3024.4]
  reg  _T_103; // @[package.scala 48:56:@3025.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@3038.4 package.scala 96:25:@3039.4]
  wire  _T_110; // @[package.scala 100:49:@3040.4]
  reg  _T_113; // @[package.scala 48:56:@3041.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@3043.4]
  wire  _T_118; // @[Controllers.scala 283:41:@3048.4]
  wire  _T_124; // @[package.scala 96:25:@3060.4 package.scala 96:25:@3061.4]
  wire  _T_126; // @[package.scala 100:49:@3062.4]
  reg  _T_129; // @[package.scala 48:56:@3063.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@3085.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@3087.4]
  reg  _T_153; // @[package.scala 48:56:@3088.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@3096.4 package.scala 96:25:@3097.4]
  wire  _T_158; // @[Controllers.scala 292:61:@3098.4]
  wire  _T_159; // @[Controllers.scala 292:24:@3099.4]
  SRFF active ( // @[Controllers.scala 261:22:@2996.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@2999.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_13 RetimeWrapper ( // @[package.scala 93:22:@3033.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_13 RetimeWrapper_1 ( // @[package.scala 93:22:@3055.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@3067.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@3075.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@3091.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@3004.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@3005.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@3006.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@3024.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@3038.4 package.scala 96:25:@3039.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@3040.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@3043.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@3048.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@3060.4 package.scala 96:25:@3061.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@3062.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@3087.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@3096.4 package.scala 96:25:@3097.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@3098.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@3099.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@3066.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@3101.4]
  assign io_datapathEn = _T_118 & io_enable; // @[Controllers.scala 283:21:@3051.4]
  assign io_ctrInc = active_io_output & io_enable; // @[Controllers.scala 284:17:@3054.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@3046.4]
  assign active_clock = clock; // @[:@2997.4]
  assign active_reset = reset; // @[:@2998.4]
  assign active_io_input_set = _T_81 & _T_82; // @[Controllers.scala 264:23:@3009.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@3013.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@3014.4]
  assign done_clock = clock; // @[:@3000.4]
  assign done_reset = reset; // @[:@3001.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@3029.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@3022.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@3023.4]
  assign RetimeWrapper_clock = clock; // @[:@3034.4]
  assign RetimeWrapper_reset = reset; // @[:@3035.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@3036.4]
  assign RetimeWrapper_1_clock = clock; // @[:@3056.4]
  assign RetimeWrapper_1_reset = reset; // @[:@3057.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@3058.4]
  assign RetimeWrapper_2_clock = clock; // @[:@3068.4]
  assign RetimeWrapper_2_reset = reset; // @[:@3069.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@3071.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@3070.4]
  assign RetimeWrapper_3_clock = clock; // @[:@3076.4]
  assign RetimeWrapper_3_reset = reset; // @[:@3077.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@3079.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@3078.4]
  assign RetimeWrapper_4_clock = clock; // @[:@3092.4]
  assign RetimeWrapper_4_reset = reset; // @[:@3093.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@3095.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@3094.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module fix2fixBox( // @[:@3207.2]
  input  [31:0] io_a, // @[:@3210.4]
  output [31:0] io_b // @[:@3210.4]
);
  assign io_b = io_a; // @[Converter.scala 95:38:@3220.4]
endmodule
module _( // @[:@3222.2]
  input  [31:0] io_b, // @[:@3225.4]
  output [31:0] io_result // @[:@3225.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@3230.4]
  wire [31:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@3230.4]
  fix2fixBox fix2fixBox ( // @[BigIPZynq.scala 219:30:@3230.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 706:17:@3238.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@3233.4]
endmodule
module RetimeWrapper_36( // @[:@3252.2]
  input          clock, // @[:@3253.4]
  input          reset, // @[:@3254.4]
  input  [368:0] io_in, // @[:@3255.4]
  output [368:0] io_out // @[:@3255.4]
);
  wire [368:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@3257.4]
  wire [368:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@3257.4]
  wire [368:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@3257.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3257.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3257.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3257.4]
  RetimeShiftRegister #(.WIDTH(369), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@3257.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3270.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3269.4]
  assign sr_init = 369'h0; // @[RetimeShiftRegister.scala 19:16:@3268.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@3267.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3266.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3264.4]
endmodule
module RetimeWrapper_37( // @[:@3284.2]
  input         clock, // @[:@3285.4]
  input         reset, // @[:@3286.4]
  input  [31:0] io_in, // @[:@3287.4]
  output [31:0] io_out // @[:@3287.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@3289.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@3289.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@3289.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3289.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3289.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3289.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@3289.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3302.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3301.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@3300.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@3299.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3298.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3296.4]
endmodule
module x465_inr_Foreach_kernelx465_inr_Foreach_concrete1( // @[:@3400.2]
  input          clock, // @[:@3401.4]
  input          reset, // @[:@3402.4]
  output         io_in_x416_TREADY, // @[:@3403.4]
  input  [255:0] io_in_x416_TDATA, // @[:@3403.4]
  output [3:0]   io_in_x452_a_0_wPort_0_banks_0, // @[:@3403.4]
  output [2:0]   io_in_x452_a_0_wPort_0_ofs_0, // @[:@3403.4]
  output [63:0]  io_in_x452_a_0_wPort_0_data_0, // @[:@3403.4]
  output         io_in_x452_a_0_wPort_0_en_0, // @[:@3403.4]
  input          io_sigsIn_datapathEn, // @[:@3403.4]
  input          io_sigsIn_break, // @[:@3403.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_0, // @[:@3403.4]
  input          io_sigsIn_cchainOutputs_0_oobs_0, // @[:@3403.4]
  input          io_rr // @[:@3403.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@3465.4]
  wire [31:0] __io_result; // @[Math.scala 709:24:@3465.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3479.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3479.4]
  wire [368:0] RetimeWrapper_io_in; // @[package.scala 93:22:@3479.4]
  wire [368:0] RetimeWrapper_io_out; // @[package.scala 93:22:@3479.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@3521.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@3521.4]
  wire [31:0] RetimeWrapper_1_io_in; // @[package.scala 93:22:@3521.4]
  wire [31:0] RetimeWrapper_1_io_out; // @[package.scala 93:22:@3521.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@3530.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@3530.4]
  wire [31:0] RetimeWrapper_2_io_in; // @[package.scala 93:22:@3530.4]
  wire [31:0] RetimeWrapper_2_io_out; // @[package.scala 93:22:@3530.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@3539.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@3539.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@3539.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@3539.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@3539.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@3550.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@3550.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@3550.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@3550.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@3550.4]
  wire  b456; // @[sm_x465_inr_Foreach.scala 62:18:@3473.4]
  wire [31:0] b455_number; // @[Math.scala 712:22:@3470.4 Math.scala 713:14:@3471.4]
  wire [31:0] _T_654; // @[Math.scala 406:49:@3493.4]
  wire [31:0] _T_656; // @[Math.scala 406:56:@3495.4]
  wire [31:0] _T_657; // @[Math.scala 406:56:@3496.4]
  wire [31:0] x780_number; // @[implicits.scala 133:21:@3497.4]
  wire [31:0] _T_667; // @[Math.scala 406:49:@3504.4]
  wire [31:0] _T_669; // @[Math.scala 406:56:@3506.4]
  wire [31:0] _T_670; // @[Math.scala 406:56:@3507.4]
  wire  _T_676; // @[FixedPoint.scala 50:25:@3513.4]
  wire [2:0] _T_680; // @[Bitwise.scala 72:12:@3515.4]
  wire [28:0] _T_681; // @[FixedPoint.scala 18:52:@3516.4]
  wire  _T_692; // @[sm_x465_inr_Foreach.scala 86:96:@3547.4]
  wire  _T_696; // @[package.scala 96:25:@3555.4 package.scala 96:25:@3556.4]
  wire  _T_698; // @[implicits.scala 55:10:@3557.4]
  wire  _T_699; // @[sm_x465_inr_Foreach.scala 86:113:@3558.4]
  wire  _T_701; // @[sm_x465_inr_Foreach.scala 86:200:@3560.4]
  wire  x785_b456_D1; // @[package.scala 96:25:@3544.4 package.scala 96:25:@3545.4]
  wire [368:0] x782_x457_D1_0; // @[package.scala 96:25:@3484.4 package.scala 96:25:@3485.4]
  wire [31:0] x783_x781_D1_number; // @[package.scala 96:25:@3526.4 package.scala 96:25:@3527.4]
  wire [31:0] x784_x461_D1_number; // @[package.scala 96:25:@3535.4 package.scala 96:25:@3536.4]
  _ _ ( // @[Math.scala 709:24:@3465.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  RetimeWrapper_36 RetimeWrapper ( // @[package.scala 93:22:@3479.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_37 RetimeWrapper_1 ( // @[package.scala 93:22:@3521.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_37 RetimeWrapper_2 ( // @[package.scala 93:22:@3530.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@3539.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@3550.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign b456 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x465_inr_Foreach.scala 62:18:@3473.4]
  assign b455_number = __io_result; // @[Math.scala 712:22:@3470.4 Math.scala 713:14:@3471.4]
  assign _T_654 = $signed(b455_number); // @[Math.scala 406:49:@3493.4]
  assign _T_656 = $signed(_T_654) & $signed(32'sh1f); // @[Math.scala 406:56:@3495.4]
  assign _T_657 = $signed(_T_656); // @[Math.scala 406:56:@3496.4]
  assign x780_number = $unsigned(_T_657); // @[implicits.scala 133:21:@3497.4]
  assign _T_667 = $signed(x780_number); // @[Math.scala 406:49:@3504.4]
  assign _T_669 = $signed(_T_667) & $signed(32'sh7); // @[Math.scala 406:56:@3506.4]
  assign _T_670 = $signed(_T_669); // @[Math.scala 406:56:@3507.4]
  assign _T_676 = x780_number[31]; // @[FixedPoint.scala 50:25:@3513.4]
  assign _T_680 = _T_676 ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12:@3515.4]
  assign _T_681 = x780_number[31:3]; // @[FixedPoint.scala 18:52:@3516.4]
  assign _T_692 = ~ io_sigsIn_break; // @[sm_x465_inr_Foreach.scala 86:96:@3547.4]
  assign _T_696 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@3555.4 package.scala 96:25:@3556.4]
  assign _T_698 = io_rr ? _T_696 : 1'h0; // @[implicits.scala 55:10:@3557.4]
  assign _T_699 = _T_692 & _T_698; // @[sm_x465_inr_Foreach.scala 86:113:@3558.4]
  assign _T_701 = _T_699 & _T_692; // @[sm_x465_inr_Foreach.scala 86:200:@3560.4]
  assign x785_b456_D1 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@3544.4 package.scala 96:25:@3545.4]
  assign x782_x457_D1_0 = RetimeWrapper_io_out; // @[package.scala 96:25:@3484.4 package.scala 96:25:@3485.4]
  assign x783_x781_D1_number = RetimeWrapper_1_io_out; // @[package.scala 96:25:@3526.4 package.scala 96:25:@3527.4]
  assign x784_x461_D1_number = RetimeWrapper_2_io_out; // @[package.scala 96:25:@3535.4 package.scala 96:25:@3536.4]
  assign io_in_x416_TREADY = b456 & io_sigsIn_datapathEn; // @[sm_x465_inr_Foreach.scala 64:18:@3476.4]
  assign io_in_x452_a_0_wPort_0_banks_0 = x783_x781_D1_number[3:0]; // @[MemInterfaceType.scala 88:58:@3563.4]
  assign io_in_x452_a_0_wPort_0_ofs_0 = x784_x461_D1_number[2:0]; // @[MemInterfaceType.scala 89:54:@3564.4]
  assign io_in_x452_a_0_wPort_0_data_0 = x782_x457_D1_0[63:0]; // @[MemInterfaceType.scala 90:56:@3565.4]
  assign io_in_x452_a_0_wPort_0_en_0 = _T_701 & x785_b456_D1; // @[MemInterfaceType.scala 93:57:@3567.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 710:17:@3468.4]
  assign RetimeWrapper_clock = clock; // @[:@3480.4]
  assign RetimeWrapper_reset = reset; // @[:@3481.4]
  assign RetimeWrapper_io_in = {{113'd0}, io_in_x416_TDATA}; // @[package.scala 94:16:@3482.4]
  assign RetimeWrapper_1_clock = clock; // @[:@3522.4]
  assign RetimeWrapper_1_reset = reset; // @[:@3523.4]
  assign RetimeWrapper_1_io_in = $unsigned(_T_670); // @[package.scala 94:16:@3524.4]
  assign RetimeWrapper_2_clock = clock; // @[:@3531.4]
  assign RetimeWrapper_2_reset = reset; // @[:@3532.4]
  assign RetimeWrapper_2_io_in = {_T_680,_T_681}; // @[package.scala 94:16:@3533.4]
  assign RetimeWrapper_3_clock = clock; // @[:@3540.4]
  assign RetimeWrapper_3_reset = reset; // @[:@3541.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@3543.4]
  assign RetimeWrapper_3_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@3542.4]
  assign RetimeWrapper_4_clock = clock; // @[:@3551.4]
  assign RetimeWrapper_4_reset = reset; // @[:@3552.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@3554.4]
  assign RetimeWrapper_4_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@3553.4]
endmodule
module x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1( // @[:@3569.2]
  input          clock, // @[:@3570.4]
  input          reset, // @[:@3571.4]
  input          io_in_x416_TVALID, // @[:@3572.4]
  output         io_in_x416_TREADY, // @[:@3572.4]
  input  [255:0] io_in_x416_TDATA, // @[:@3572.4]
  output [3:0]   io_in_x452_a_0_wPort_0_banks_0, // @[:@3572.4]
  output [2:0]   io_in_x452_a_0_wPort_0_ofs_0, // @[:@3572.4]
  output [63:0]  io_in_x452_a_0_wPort_0_data_0, // @[:@3572.4]
  output         io_in_x452_a_0_wPort_0_en_0, // @[:@3572.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@3572.4]
  input          io_sigsIn_smChildAcks_0, // @[:@3572.4]
  output         io_sigsOut_smDoneIn_0, // @[:@3572.4]
  output         io_sigsOut_smCtrCopyDone_0, // @[:@3572.4]
  input          io_rr // @[:@3572.4]
);
  wire  x454_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@3630.4]
  wire  x454_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@3630.4]
  wire  x454_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@3630.4]
  wire  x454_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@3630.4]
  wire [31:0] x454_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@3630.4]
  wire  x454_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@3630.4]
  wire  x454_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@3630.4]
  wire  x465_inr_Foreach_sm_clock; // @[sm_x465_inr_Foreach.scala 33:18:@3682.4]
  wire  x465_inr_Foreach_sm_reset; // @[sm_x465_inr_Foreach.scala 33:18:@3682.4]
  wire  x465_inr_Foreach_sm_io_enable; // @[sm_x465_inr_Foreach.scala 33:18:@3682.4]
  wire  x465_inr_Foreach_sm_io_done; // @[sm_x465_inr_Foreach.scala 33:18:@3682.4]
  wire  x465_inr_Foreach_sm_io_doneLatch; // @[sm_x465_inr_Foreach.scala 33:18:@3682.4]
  wire  x465_inr_Foreach_sm_io_ctrDone; // @[sm_x465_inr_Foreach.scala 33:18:@3682.4]
  wire  x465_inr_Foreach_sm_io_datapathEn; // @[sm_x465_inr_Foreach.scala 33:18:@3682.4]
  wire  x465_inr_Foreach_sm_io_ctrInc; // @[sm_x465_inr_Foreach.scala 33:18:@3682.4]
  wire  x465_inr_Foreach_sm_io_ctrRst; // @[sm_x465_inr_Foreach.scala 33:18:@3682.4]
  wire  x465_inr_Foreach_sm_io_parentAck; // @[sm_x465_inr_Foreach.scala 33:18:@3682.4]
  wire  x465_inr_Foreach_sm_io_break; // @[sm_x465_inr_Foreach.scala 33:18:@3682.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3710.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3710.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3710.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@3710.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@3710.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@3750.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@3750.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@3750.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@3750.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@3750.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@3758.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@3758.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@3758.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@3758.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@3758.4]
  wire  x465_inr_Foreach_kernelx465_inr_Foreach_concrete1_clock; // @[sm_x465_inr_Foreach.scala 88:24:@3790.4]
  wire  x465_inr_Foreach_kernelx465_inr_Foreach_concrete1_reset; // @[sm_x465_inr_Foreach.scala 88:24:@3790.4]
  wire  x465_inr_Foreach_kernelx465_inr_Foreach_concrete1_io_in_x416_TREADY; // @[sm_x465_inr_Foreach.scala 88:24:@3790.4]
  wire [255:0] x465_inr_Foreach_kernelx465_inr_Foreach_concrete1_io_in_x416_TDATA; // @[sm_x465_inr_Foreach.scala 88:24:@3790.4]
  wire [3:0] x465_inr_Foreach_kernelx465_inr_Foreach_concrete1_io_in_x452_a_0_wPort_0_banks_0; // @[sm_x465_inr_Foreach.scala 88:24:@3790.4]
  wire [2:0] x465_inr_Foreach_kernelx465_inr_Foreach_concrete1_io_in_x452_a_0_wPort_0_ofs_0; // @[sm_x465_inr_Foreach.scala 88:24:@3790.4]
  wire [63:0] x465_inr_Foreach_kernelx465_inr_Foreach_concrete1_io_in_x452_a_0_wPort_0_data_0; // @[sm_x465_inr_Foreach.scala 88:24:@3790.4]
  wire  x465_inr_Foreach_kernelx465_inr_Foreach_concrete1_io_in_x452_a_0_wPort_0_en_0; // @[sm_x465_inr_Foreach.scala 88:24:@3790.4]
  wire  x465_inr_Foreach_kernelx465_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x465_inr_Foreach.scala 88:24:@3790.4]
  wire  x465_inr_Foreach_kernelx465_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x465_inr_Foreach.scala 88:24:@3790.4]
  wire [31:0] x465_inr_Foreach_kernelx465_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x465_inr_Foreach.scala 88:24:@3790.4]
  wire  x465_inr_Foreach_kernelx465_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x465_inr_Foreach.scala 88:24:@3790.4]
  wire  x465_inr_Foreach_kernelx465_inr_Foreach_concrete1_io_rr; // @[sm_x465_inr_Foreach.scala 88:24:@3790.4]
  wire  _T_683; // @[package.scala 96:25:@3715.4 package.scala 96:25:@3716.4]
  wire  x465_inr_Foreach_sigsIn_forwardpressure; // @[sm_x466_outr_UnitPipe.scala 68:54:@3721.4]
  wire  _T_697; // @[package.scala 96:25:@3755.4 package.scala 96:25:@3756.4]
  wire  _T_703; // @[package.scala 96:25:@3763.4 package.scala 96:25:@3764.4]
  wire  _T_706; // @[SpatialBlocks.scala 110:93:@3766.4]
  wire  x465_inr_Foreach_sigsIn_baseEn; // @[SpatialBlocks.scala 110:90:@3767.4]
  wire  _T_708; // @[SpatialBlocks.scala 128:36:@3775.4]
  wire  _T_709; // @[SpatialBlocks.scala 128:78:@3776.4]
  wire  _T_714; // @[SpatialBlocks.scala 130:61:@3785.4]
  x454_ctrchain x454_ctrchain ( // @[SpatialBlocks.scala 37:22:@3630.4]
    .clock(x454_ctrchain_clock),
    .reset(x454_ctrchain_reset),
    .io_input_reset(x454_ctrchain_io_input_reset),
    .io_input_enable(x454_ctrchain_io_input_enable),
    .io_output_counts_0(x454_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x454_ctrchain_io_output_oobs_0),
    .io_output_done(x454_ctrchain_io_output_done)
  );
  x465_inr_Foreach_sm x465_inr_Foreach_sm ( // @[sm_x465_inr_Foreach.scala 33:18:@3682.4]
    .clock(x465_inr_Foreach_sm_clock),
    .reset(x465_inr_Foreach_sm_reset),
    .io_enable(x465_inr_Foreach_sm_io_enable),
    .io_done(x465_inr_Foreach_sm_io_done),
    .io_doneLatch(x465_inr_Foreach_sm_io_doneLatch),
    .io_ctrDone(x465_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x465_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x465_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x465_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x465_inr_Foreach_sm_io_parentAck),
    .io_break(x465_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@3710.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@3750.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@3758.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x465_inr_Foreach_kernelx465_inr_Foreach_concrete1 x465_inr_Foreach_kernelx465_inr_Foreach_concrete1 ( // @[sm_x465_inr_Foreach.scala 88:24:@3790.4]
    .clock(x465_inr_Foreach_kernelx465_inr_Foreach_concrete1_clock),
    .reset(x465_inr_Foreach_kernelx465_inr_Foreach_concrete1_reset),
    .io_in_x416_TREADY(x465_inr_Foreach_kernelx465_inr_Foreach_concrete1_io_in_x416_TREADY),
    .io_in_x416_TDATA(x465_inr_Foreach_kernelx465_inr_Foreach_concrete1_io_in_x416_TDATA),
    .io_in_x452_a_0_wPort_0_banks_0(x465_inr_Foreach_kernelx465_inr_Foreach_concrete1_io_in_x452_a_0_wPort_0_banks_0),
    .io_in_x452_a_0_wPort_0_ofs_0(x465_inr_Foreach_kernelx465_inr_Foreach_concrete1_io_in_x452_a_0_wPort_0_ofs_0),
    .io_in_x452_a_0_wPort_0_data_0(x465_inr_Foreach_kernelx465_inr_Foreach_concrete1_io_in_x452_a_0_wPort_0_data_0),
    .io_in_x452_a_0_wPort_0_en_0(x465_inr_Foreach_kernelx465_inr_Foreach_concrete1_io_in_x452_a_0_wPort_0_en_0),
    .io_sigsIn_datapathEn(x465_inr_Foreach_kernelx465_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x465_inr_Foreach_kernelx465_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_0(x465_inr_Foreach_kernelx465_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x465_inr_Foreach_kernelx465_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_rr(x465_inr_Foreach_kernelx465_inr_Foreach_concrete1_io_rr)
  );
  assign _T_683 = RetimeWrapper_io_out; // @[package.scala 96:25:@3715.4 package.scala 96:25:@3716.4]
  assign x465_inr_Foreach_sigsIn_forwardpressure = io_in_x416_TVALID | x465_inr_Foreach_sm_io_doneLatch; // @[sm_x466_outr_UnitPipe.scala 68:54:@3721.4]
  assign _T_697 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@3755.4 package.scala 96:25:@3756.4]
  assign _T_703 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@3763.4 package.scala 96:25:@3764.4]
  assign _T_706 = ~ _T_703; // @[SpatialBlocks.scala 110:93:@3766.4]
  assign x465_inr_Foreach_sigsIn_baseEn = _T_697 & _T_706; // @[SpatialBlocks.scala 110:90:@3767.4]
  assign _T_708 = x465_inr_Foreach_sm_io_datapathEn; // @[SpatialBlocks.scala 128:36:@3775.4]
  assign _T_709 = ~ x465_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 128:78:@3776.4]
  assign _T_714 = x465_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 130:61:@3785.4]
  assign io_in_x416_TREADY = x465_inr_Foreach_kernelx465_inr_Foreach_concrete1_io_in_x416_TREADY; // @[sm_x465_inr_Foreach.scala 49:23:@3882.4]
  assign io_in_x452_a_0_wPort_0_banks_0 = x465_inr_Foreach_kernelx465_inr_Foreach_concrete1_io_in_x452_a_0_wPort_0_banks_0; // @[MemInterfaceType.scala 67:44:@3890.4]
  assign io_in_x452_a_0_wPort_0_ofs_0 = x465_inr_Foreach_kernelx465_inr_Foreach_concrete1_io_in_x452_a_0_wPort_0_ofs_0; // @[MemInterfaceType.scala 67:44:@3889.4]
  assign io_in_x452_a_0_wPort_0_data_0 = x465_inr_Foreach_kernelx465_inr_Foreach_concrete1_io_in_x452_a_0_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@3888.4]
  assign io_in_x452_a_0_wPort_0_en_0 = x465_inr_Foreach_kernelx465_inr_Foreach_concrete1_io_in_x452_a_0_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@3884.4]
  assign io_sigsOut_smDoneIn_0 = x465_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 127:53:@3773.4]
  assign io_sigsOut_smCtrCopyDone_0 = x465_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 139:125:@3789.4]
  assign x454_ctrchain_clock = clock; // @[:@3631.4]
  assign x454_ctrchain_reset = reset; // @[:@3632.4]
  assign x454_ctrchain_io_input_reset = x465_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 130:103:@3788.4]
  assign x454_ctrchain_io_input_enable = _T_714 & x465_inr_Foreach_sigsIn_forwardpressure; // @[SpatialBlocks.scala 104:75:@3743.4 SpatialBlocks.scala 130:45:@3787.4]
  assign x465_inr_Foreach_sm_clock = clock; // @[:@3683.4]
  assign x465_inr_Foreach_sm_reset = reset; // @[:@3684.4]
  assign x465_inr_Foreach_sm_io_enable = x465_inr_Foreach_sigsIn_baseEn & x465_inr_Foreach_sigsIn_forwardpressure; // @[SpatialBlocks.scala 112:18:@3770.4]
  assign x465_inr_Foreach_sm_io_ctrDone = io_rr ? _T_683 : 1'h0; // @[sm_x466_outr_UnitPipe.scala 66:38:@3718.4]
  assign x465_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 114:21:@3772.4]
  assign x465_inr_Foreach_sm_io_break = 1'h0; // @[sm_x466_outr_UnitPipe.scala 70:36:@3724.4]
  assign RetimeWrapper_clock = clock; // @[:@3711.4]
  assign RetimeWrapper_reset = reset; // @[:@3712.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@3714.4]
  assign RetimeWrapper_io_in = x454_ctrchain_io_output_done; // @[package.scala 94:16:@3713.4]
  assign RetimeWrapper_1_clock = clock; // @[:@3751.4]
  assign RetimeWrapper_1_reset = reset; // @[:@3752.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@3754.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@3753.4]
  assign RetimeWrapper_2_clock = clock; // @[:@3759.4]
  assign RetimeWrapper_2_reset = reset; // @[:@3760.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@3762.4]
  assign RetimeWrapper_2_io_in = x465_inr_Foreach_sm_io_done; // @[package.scala 94:16:@3761.4]
  assign x465_inr_Foreach_kernelx465_inr_Foreach_concrete1_clock = clock; // @[:@3791.4]
  assign x465_inr_Foreach_kernelx465_inr_Foreach_concrete1_reset = reset; // @[:@3792.4]
  assign x465_inr_Foreach_kernelx465_inr_Foreach_concrete1_io_in_x416_TDATA = io_in_x416_TDATA; // @[sm_x465_inr_Foreach.scala 49:23:@3881.4]
  assign x465_inr_Foreach_kernelx465_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_708 & _T_709; // @[sm_x465_inr_Foreach.scala 92:22:@3903.4]
  assign x465_inr_Foreach_kernelx465_inr_Foreach_concrete1_io_sigsIn_break = x465_inr_Foreach_sm_io_break; // @[sm_x465_inr_Foreach.scala 92:22:@3901.4]
  assign x465_inr_Foreach_kernelx465_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = x454_ctrchain_io_output_counts_0; // @[sm_x465_inr_Foreach.scala 92:22:@3896.4]
  assign x465_inr_Foreach_kernelx465_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x454_ctrchain_io_output_oobs_0; // @[sm_x465_inr_Foreach.scala 92:22:@3895.4]
  assign x465_inr_Foreach_kernelx465_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x465_inr_Foreach.scala 91:18:@3891.4]
endmodule
module RetimeWrapper_41( // @[:@3956.2]
  input   clock, // @[:@3957.4]
  input   reset, // @[:@3958.4]
  input   io_in, // @[:@3959.4]
  output  io_out // @[:@3959.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@3961.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@3961.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@3961.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3961.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3961.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3961.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@3961.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3974.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3973.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@3972.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@3971.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3970.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3968.4]
endmodule
module x555_inr_UnitPipe_sm( // @[:@4104.2]
  input   clock, // @[:@4105.4]
  input   reset, // @[:@4106.4]
  input   io_enable, // @[:@4107.4]
  output  io_done, // @[:@4107.4]
  input   io_ctrDone, // @[:@4107.4]
  output  io_datapathEn, // @[:@4107.4]
  output  io_ctrInc, // @[:@4107.4]
  input   io_parentAck, // @[:@4107.4]
  input   io_break // @[:@4107.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@4109.4]
  wire  active_reset; // @[Controllers.scala 261:22:@4109.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@4109.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@4109.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@4109.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@4109.4]
  wire  done_clock; // @[Controllers.scala 262:20:@4112.4]
  wire  done_reset; // @[Controllers.scala 262:20:@4112.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@4112.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@4112.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@4112.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@4112.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@4146.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@4146.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@4146.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@4146.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@4168.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@4168.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@4168.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@4168.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@4180.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@4180.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@4180.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@4180.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@4180.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@4188.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@4188.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@4188.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@4188.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@4188.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@4204.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@4204.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@4204.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@4204.4]
  wire  _T_80; // @[Controllers.scala 264:48:@4117.4]
  wire  _T_81; // @[Controllers.scala 264:46:@4118.4]
  wire  _T_82; // @[Controllers.scala 264:62:@4119.4]
  wire  _T_100; // @[package.scala 100:49:@4137.4]
  reg  _T_103; // @[package.scala 48:56:@4138.4]
  reg [31:0] _RAND_0;
  wire  _T_118; // @[Controllers.scala 283:41:@4161.4]
  wire  _T_124; // @[package.scala 96:25:@4173.4 package.scala 96:25:@4174.4]
  wire  _T_126; // @[package.scala 100:49:@4175.4]
  reg  _T_129; // @[package.scala 48:56:@4176.4]
  reg [31:0] _RAND_1;
  wire  _T_150; // @[package.scala 100:49:@4200.4]
  reg  _T_153; // @[package.scala 48:56:@4201.4]
  reg [31:0] _RAND_2;
  SRFF active ( // @[Controllers.scala 261:22:@4109.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@4112.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_41 RetimeWrapper ( // @[package.scala 93:22:@4146.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_41 RetimeWrapper_1 ( // @[package.scala 93:22:@4168.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@4180.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@4188.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_13 RetimeWrapper_4 ( // @[package.scala 93:22:@4204.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@4117.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@4118.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@4119.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@4137.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@4161.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@4173.4 package.scala 96:25:@4174.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@4175.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@4200.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@4179.4]
  assign io_datapathEn = _T_118 & io_enable; // @[Controllers.scala 283:21:@4164.4]
  assign io_ctrInc = active_io_output & io_enable; // @[Controllers.scala 284:17:@4167.4]
  assign active_clock = clock; // @[:@4110.4]
  assign active_reset = reset; // @[:@4111.4]
  assign active_io_input_set = _T_81 & _T_82; // @[Controllers.scala 264:23:@4122.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@4126.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@4127.4]
  assign done_clock = clock; // @[:@4113.4]
  assign done_reset = reset; // @[:@4114.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@4142.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@4135.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@4136.4]
  assign RetimeWrapper_clock = clock; // @[:@4147.4]
  assign RetimeWrapper_reset = reset; // @[:@4148.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@4149.4]
  assign RetimeWrapper_1_clock = clock; // @[:@4169.4]
  assign RetimeWrapper_1_reset = reset; // @[:@4170.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@4171.4]
  assign RetimeWrapper_2_clock = clock; // @[:@4181.4]
  assign RetimeWrapper_2_reset = reset; // @[:@4182.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@4184.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@4183.4]
  assign RetimeWrapper_3_clock = clock; // @[:@4189.4]
  assign RetimeWrapper_3_reset = reset; // @[:@4190.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@4192.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@4191.4]
  assign RetimeWrapper_4_clock = clock; // @[:@4205.4]
  assign RetimeWrapper_4_reset = reset; // @[:@4206.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@4207.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_129 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_153 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1( // @[:@5312.2]
  input         clock, // @[:@5313.4]
  input         reset, // @[:@5314.4]
  output        io_in_x449_argOut_port_0_valid, // @[:@5315.4]
  output [63:0] io_in_x449_argOut_port_0_bits, // @[:@5315.4]
  output        io_in_x440_argOut_port_0_valid, // @[:@5315.4]
  output [63:0] io_in_x440_argOut_port_0_bits, // @[:@5315.4]
  output        io_in_x436_argOut_port_0_valid, // @[:@5315.4]
  output [63:0] io_in_x436_argOut_port_0_bits, // @[:@5315.4]
  output        io_in_x421_argOut_port_0_valid, // @[:@5315.4]
  output [63:0] io_in_x421_argOut_port_0_bits, // @[:@5315.4]
  output        io_in_x448_argOut_port_0_valid, // @[:@5315.4]
  output [63:0] io_in_x448_argOut_port_0_bits, // @[:@5315.4]
  output        io_in_x443_argOut_port_0_valid, // @[:@5315.4]
  output [63:0] io_in_x443_argOut_port_0_bits, // @[:@5315.4]
  output        io_in_x428_argOut_port_0_valid, // @[:@5315.4]
  output [63:0] io_in_x428_argOut_port_0_bits, // @[:@5315.4]
  output        io_in_x452_a_0_rPort_7_en_0, // @[:@5315.4]
  input  [63:0] io_in_x452_a_0_rPort_7_output_0, // @[:@5315.4]
  output        io_in_x452_a_0_rPort_6_en_0, // @[:@5315.4]
  input  [63:0] io_in_x452_a_0_rPort_6_output_0, // @[:@5315.4]
  output        io_in_x452_a_0_rPort_5_en_0, // @[:@5315.4]
  input  [63:0] io_in_x452_a_0_rPort_5_output_0, // @[:@5315.4]
  output        io_in_x452_a_0_rPort_4_en_0, // @[:@5315.4]
  input  [63:0] io_in_x452_a_0_rPort_4_output_0, // @[:@5315.4]
  output        io_in_x452_a_0_rPort_3_en_0, // @[:@5315.4]
  input  [63:0] io_in_x452_a_0_rPort_3_output_0, // @[:@5315.4]
  output        io_in_x452_a_0_rPort_2_en_0, // @[:@5315.4]
  input  [63:0] io_in_x452_a_0_rPort_2_output_0, // @[:@5315.4]
  output        io_in_x452_a_0_rPort_1_en_0, // @[:@5315.4]
  input  [63:0] io_in_x452_a_0_rPort_1_output_0, // @[:@5315.4]
  output        io_in_x452_a_0_rPort_0_en_0, // @[:@5315.4]
  input  [63:0] io_in_x452_a_0_rPort_0_output_0, // @[:@5315.4]
  output        io_in_x439_argOut_port_0_valid, // @[:@5315.4]
  output [63:0] io_in_x439_argOut_port_0_bits, // @[:@5315.4]
  output        io_in_x424_argOut_port_0_valid, // @[:@5315.4]
  output [63:0] io_in_x424_argOut_port_0_bits, // @[:@5315.4]
  output        io_in_x429_argOut_port_0_valid, // @[:@5315.4]
  output [63:0] io_in_x429_argOut_port_0_bits, // @[:@5315.4]
  output        io_in_x435_argOut_port_0_valid, // @[:@5315.4]
  output [63:0] io_in_x435_argOut_port_0_bits, // @[:@5315.4]
  output        io_in_x420_argOut_port_0_valid, // @[:@5315.4]
  output [63:0] io_in_x420_argOut_port_0_bits, // @[:@5315.4]
  output        io_in_x425_argOut_port_0_valid, // @[:@5315.4]
  output [63:0] io_in_x425_argOut_port_0_bits, // @[:@5315.4]
  output        io_in_x430_argOut_port_0_valid, // @[:@5315.4]
  output [63:0] io_in_x430_argOut_port_0_bits, // @[:@5315.4]
  output        io_in_x444_argOut_port_0_valid, // @[:@5315.4]
  output [63:0] io_in_x444_argOut_port_0_bits, // @[:@5315.4]
  output        io_in_x423_argOut_port_0_valid, // @[:@5315.4]
  output [63:0] io_in_x423_argOut_port_0_bits, // @[:@5315.4]
  output        io_in_x445_argOut_port_0_valid, // @[:@5315.4]
  output [63:0] io_in_x445_argOut_port_0_bits, // @[:@5315.4]
  output        io_in_x451_argOut_port_0_valid, // @[:@5315.4]
  output [63:0] io_in_x451_argOut_port_0_bits, // @[:@5315.4]
  output        io_in_x434_argOut_port_0_valid, // @[:@5315.4]
  output [63:0] io_in_x434_argOut_port_0_bits, // @[:@5315.4]
  output        io_in_x438_argOut_port_0_valid, // @[:@5315.4]
  output [63:0] io_in_x438_argOut_port_0_bits, // @[:@5315.4]
  output        io_in_x431_argOut_port_0_valid, // @[:@5315.4]
  output [63:0] io_in_x431_argOut_port_0_bits, // @[:@5315.4]
  output        io_in_x426_argOut_port_0_valid, // @[:@5315.4]
  output [63:0] io_in_x426_argOut_port_0_bits, // @[:@5315.4]
  output        io_in_x441_argOut_port_0_valid, // @[:@5315.4]
  output [63:0] io_in_x441_argOut_port_0_bits, // @[:@5315.4]
  output        io_in_x446_argOut_port_0_valid, // @[:@5315.4]
  output [63:0] io_in_x446_argOut_port_0_bits, // @[:@5315.4]
  output        io_in_x450_argOut_port_0_valid, // @[:@5315.4]
  output [63:0] io_in_x450_argOut_port_0_bits, // @[:@5315.4]
  output        io_in_x433_argOut_port_0_valid, // @[:@5315.4]
  output [63:0] io_in_x433_argOut_port_0_bits, // @[:@5315.4]
  output        io_in_x447_argOut_port_0_valid, // @[:@5315.4]
  output [63:0] io_in_x447_argOut_port_0_bits, // @[:@5315.4]
  output        io_in_x432_argOut_port_0_valid, // @[:@5315.4]
  output [63:0] io_in_x432_argOut_port_0_bits, // @[:@5315.4]
  output        io_in_x422_argOut_port_0_valid, // @[:@5315.4]
  output [63:0] io_in_x422_argOut_port_0_bits, // @[:@5315.4]
  output        io_in_x437_argOut_port_0_valid, // @[:@5315.4]
  output [63:0] io_in_x437_argOut_port_0_bits, // @[:@5315.4]
  output        io_in_x427_argOut_port_0_valid, // @[:@5315.4]
  output [63:0] io_in_x427_argOut_port_0_bits, // @[:@5315.4]
  output        io_in_x442_argOut_port_0_valid, // @[:@5315.4]
  output [63:0] io_in_x442_argOut_port_0_bits, // @[:@5315.4]
  input         io_sigsIn_datapathEn, // @[:@5315.4]
  input         io_sigsIn_break, // @[:@5315.4]
  input         io_rr // @[:@5315.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@5531.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@5531.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@5531.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@5531.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@5544.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@5544.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@5544.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@5544.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@5557.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@5557.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@5557.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@5557.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@5570.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@5570.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@5570.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@5570.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@5610.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@5610.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@5610.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@5610.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@5623.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@5623.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@5623.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@5623.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@5636.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@5636.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@5636.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@5636.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@5649.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@5649.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@5649.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@5649.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@5689.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@5689.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@5689.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@5689.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@5702.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@5702.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@5702.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@5702.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@5715.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@5715.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@5715.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@5715.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@5728.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@5728.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@5728.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@5728.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@5768.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@5768.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@5768.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@5768.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@5781.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@5781.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@5781.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@5781.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@5794.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@5794.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@5794.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@5794.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@5807.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@5807.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@5807.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@5807.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@5847.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@5847.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@5847.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@5847.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@5860.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@5860.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@5860.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@5860.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@5873.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@5873.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@5873.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@5873.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@5886.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@5886.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@5886.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@5886.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@5926.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@5926.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@5926.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@5926.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@5939.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@5939.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@5939.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@5939.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@5952.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@5952.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@5952.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@5952.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@5965.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@5965.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@5965.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@5965.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@6005.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@6005.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@6005.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@6005.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@6018.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@6018.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@6018.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@6018.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@6031.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@6031.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@6031.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@6031.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@6044.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@6044.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@6044.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@6044.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@6084.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@6084.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@6084.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@6084.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@6097.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@6097.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@6097.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@6097.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@6110.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@6110.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@6110.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@6110.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@6123.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@6123.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@6123.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@6123.4]
  wire  _T_1262; // @[sm_x555_inr_UnitPipe.scala 223:128:@5506.4]
  wire  _T_1266; // @[implicits.scala 55:10:@5509.4]
  wire [15:0] x469_0_number; // @[FixedPoint.scala 18:52:@5520.4]
  wire [15:0] x469_1_number; // @[FixedPoint.scala 18:52:@5522.4]
  wire [15:0] x469_2_number; // @[FixedPoint.scala 18:52:@5524.4]
  wire [15:0] x469_3_number; // @[FixedPoint.scala 18:52:@5526.4]
  wire [15:0] x480_0_number; // @[FixedPoint.scala 18:52:@5599.4]
  wire [15:0] x480_1_number; // @[FixedPoint.scala 18:52:@5601.4]
  wire [15:0] x480_2_number; // @[FixedPoint.scala 18:52:@5603.4]
  wire [15:0] x480_3_number; // @[FixedPoint.scala 18:52:@5605.4]
  wire [15:0] x491_0_number; // @[FixedPoint.scala 18:52:@5678.4]
  wire [15:0] x491_1_number; // @[FixedPoint.scala 18:52:@5680.4]
  wire [15:0] x491_2_number; // @[FixedPoint.scala 18:52:@5682.4]
  wire [15:0] x491_3_number; // @[FixedPoint.scala 18:52:@5684.4]
  wire [15:0] x502_0_number; // @[FixedPoint.scala 18:52:@5757.4]
  wire [15:0] x502_1_number; // @[FixedPoint.scala 18:52:@5759.4]
  wire [15:0] x502_2_number; // @[FixedPoint.scala 18:52:@5761.4]
  wire [15:0] x502_3_number; // @[FixedPoint.scala 18:52:@5763.4]
  wire [15:0] x513_0_number; // @[FixedPoint.scala 18:52:@5836.4]
  wire [15:0] x513_1_number; // @[FixedPoint.scala 18:52:@5838.4]
  wire [15:0] x513_2_number; // @[FixedPoint.scala 18:52:@5840.4]
  wire [15:0] x513_3_number; // @[FixedPoint.scala 18:52:@5842.4]
  wire [15:0] x524_0_number; // @[FixedPoint.scala 18:52:@5915.4]
  wire [15:0] x524_1_number; // @[FixedPoint.scala 18:52:@5917.4]
  wire [15:0] x524_2_number; // @[FixedPoint.scala 18:52:@5919.4]
  wire [15:0] x524_3_number; // @[FixedPoint.scala 18:52:@5921.4]
  wire [15:0] x535_0_number; // @[FixedPoint.scala 18:52:@5994.4]
  wire [15:0] x535_1_number; // @[FixedPoint.scala 18:52:@5996.4]
  wire [15:0] x535_2_number; // @[FixedPoint.scala 18:52:@5998.4]
  wire [15:0] x535_3_number; // @[FixedPoint.scala 18:52:@6000.4]
  wire [15:0] x546_0_number; // @[FixedPoint.scala 18:52:@6073.4]
  wire [15:0] x546_1_number; // @[FixedPoint.scala 18:52:@6075.4]
  wire [15:0] x546_2_number; // @[FixedPoint.scala 18:52:@6077.4]
  wire [15:0] x546_3_number; // @[FixedPoint.scala 18:52:@6079.4]
  RetimeWrapper_13 RetimeWrapper ( // @[package.scala 93:22:@5531.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_13 RetimeWrapper_1 ( // @[package.scala 93:22:@5544.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_13 RetimeWrapper_2 ( // @[package.scala 93:22:@5557.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_13 RetimeWrapper_3 ( // @[package.scala 93:22:@5570.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_13 RetimeWrapper_4 ( // @[package.scala 93:22:@5610.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_13 RetimeWrapper_5 ( // @[package.scala 93:22:@5623.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_13 RetimeWrapper_6 ( // @[package.scala 93:22:@5636.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_13 RetimeWrapper_7 ( // @[package.scala 93:22:@5649.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_13 RetimeWrapper_8 ( // @[package.scala 93:22:@5689.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_13 RetimeWrapper_9 ( // @[package.scala 93:22:@5702.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_13 RetimeWrapper_10 ( // @[package.scala 93:22:@5715.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_13 RetimeWrapper_11 ( // @[package.scala 93:22:@5728.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_13 RetimeWrapper_12 ( // @[package.scala 93:22:@5768.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_13 RetimeWrapper_13 ( // @[package.scala 93:22:@5781.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_13 RetimeWrapper_14 ( // @[package.scala 93:22:@5794.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_13 RetimeWrapper_15 ( // @[package.scala 93:22:@5807.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_13 RetimeWrapper_16 ( // @[package.scala 93:22:@5847.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_13 RetimeWrapper_17 ( // @[package.scala 93:22:@5860.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_13 RetimeWrapper_18 ( // @[package.scala 93:22:@5873.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_13 RetimeWrapper_19 ( // @[package.scala 93:22:@5886.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_13 RetimeWrapper_20 ( // @[package.scala 93:22:@5926.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_13 RetimeWrapper_21 ( // @[package.scala 93:22:@5939.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_13 RetimeWrapper_22 ( // @[package.scala 93:22:@5952.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_13 RetimeWrapper_23 ( // @[package.scala 93:22:@5965.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_13 RetimeWrapper_24 ( // @[package.scala 93:22:@6005.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper_13 RetimeWrapper_25 ( // @[package.scala 93:22:@6018.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_13 RetimeWrapper_26 ( // @[package.scala 93:22:@6031.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_13 RetimeWrapper_27 ( // @[package.scala 93:22:@6044.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper_13 RetimeWrapper_28 ( // @[package.scala 93:22:@6084.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper_13 RetimeWrapper_29 ( // @[package.scala 93:22:@6097.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_13 RetimeWrapper_30 ( // @[package.scala 93:22:@6110.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_13 RetimeWrapper_31 ( // @[package.scala 93:22:@6123.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  assign _T_1262 = ~ io_sigsIn_break; // @[sm_x555_inr_UnitPipe.scala 223:128:@5506.4]
  assign _T_1266 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 55:10:@5509.4]
  assign x469_0_number = io_in_x452_a_0_rPort_3_output_0[15:0]; // @[FixedPoint.scala 18:52:@5520.4]
  assign x469_1_number = io_in_x452_a_0_rPort_3_output_0[31:16]; // @[FixedPoint.scala 18:52:@5522.4]
  assign x469_2_number = io_in_x452_a_0_rPort_3_output_0[47:32]; // @[FixedPoint.scala 18:52:@5524.4]
  assign x469_3_number = io_in_x452_a_0_rPort_3_output_0[63:48]; // @[FixedPoint.scala 18:52:@5526.4]
  assign x480_0_number = io_in_x452_a_0_rPort_7_output_0[15:0]; // @[FixedPoint.scala 18:52:@5599.4]
  assign x480_1_number = io_in_x452_a_0_rPort_7_output_0[31:16]; // @[FixedPoint.scala 18:52:@5601.4]
  assign x480_2_number = io_in_x452_a_0_rPort_7_output_0[47:32]; // @[FixedPoint.scala 18:52:@5603.4]
  assign x480_3_number = io_in_x452_a_0_rPort_7_output_0[63:48]; // @[FixedPoint.scala 18:52:@5605.4]
  assign x491_0_number = io_in_x452_a_0_rPort_5_output_0[15:0]; // @[FixedPoint.scala 18:52:@5678.4]
  assign x491_1_number = io_in_x452_a_0_rPort_5_output_0[31:16]; // @[FixedPoint.scala 18:52:@5680.4]
  assign x491_2_number = io_in_x452_a_0_rPort_5_output_0[47:32]; // @[FixedPoint.scala 18:52:@5682.4]
  assign x491_3_number = io_in_x452_a_0_rPort_5_output_0[63:48]; // @[FixedPoint.scala 18:52:@5684.4]
  assign x502_0_number = io_in_x452_a_0_rPort_2_output_0[15:0]; // @[FixedPoint.scala 18:52:@5757.4]
  assign x502_1_number = io_in_x452_a_0_rPort_2_output_0[31:16]; // @[FixedPoint.scala 18:52:@5759.4]
  assign x502_2_number = io_in_x452_a_0_rPort_2_output_0[47:32]; // @[FixedPoint.scala 18:52:@5761.4]
  assign x502_3_number = io_in_x452_a_0_rPort_2_output_0[63:48]; // @[FixedPoint.scala 18:52:@5763.4]
  assign x513_0_number = io_in_x452_a_0_rPort_0_output_0[15:0]; // @[FixedPoint.scala 18:52:@5836.4]
  assign x513_1_number = io_in_x452_a_0_rPort_0_output_0[31:16]; // @[FixedPoint.scala 18:52:@5838.4]
  assign x513_2_number = io_in_x452_a_0_rPort_0_output_0[47:32]; // @[FixedPoint.scala 18:52:@5840.4]
  assign x513_3_number = io_in_x452_a_0_rPort_0_output_0[63:48]; // @[FixedPoint.scala 18:52:@5842.4]
  assign x524_0_number = io_in_x452_a_0_rPort_4_output_0[15:0]; // @[FixedPoint.scala 18:52:@5915.4]
  assign x524_1_number = io_in_x452_a_0_rPort_4_output_0[31:16]; // @[FixedPoint.scala 18:52:@5917.4]
  assign x524_2_number = io_in_x452_a_0_rPort_4_output_0[47:32]; // @[FixedPoint.scala 18:52:@5919.4]
  assign x524_3_number = io_in_x452_a_0_rPort_4_output_0[63:48]; // @[FixedPoint.scala 18:52:@5921.4]
  assign x535_0_number = io_in_x452_a_0_rPort_1_output_0[15:0]; // @[FixedPoint.scala 18:52:@5994.4]
  assign x535_1_number = io_in_x452_a_0_rPort_1_output_0[31:16]; // @[FixedPoint.scala 18:52:@5996.4]
  assign x535_2_number = io_in_x452_a_0_rPort_1_output_0[47:32]; // @[FixedPoint.scala 18:52:@5998.4]
  assign x535_3_number = io_in_x452_a_0_rPort_1_output_0[63:48]; // @[FixedPoint.scala 18:52:@6000.4]
  assign x546_0_number = io_in_x452_a_0_rPort_6_output_0[15:0]; // @[FixedPoint.scala 18:52:@6073.4]
  assign x546_1_number = io_in_x452_a_0_rPort_6_output_0[31:16]; // @[FixedPoint.scala 18:52:@6075.4]
  assign x546_2_number = io_in_x452_a_0_rPort_6_output_0[47:32]; // @[FixedPoint.scala 18:52:@6077.4]
  assign x546_3_number = io_in_x452_a_0_rPort_6_output_0[63:48]; // @[FixedPoint.scala 18:52:@6079.4]
  assign io_in_x449_argOut_port_0_valid = RetimeWrapper_29_io_out; // @[MemInterfaceType.scala 311:132:@6106.4]
  assign io_in_x449_argOut_port_0_bits = {{48'd0}, x546_1_number}; // @[MemInterfaceType.scala 311:109:@6105.4]
  assign io_in_x440_argOut_port_0_valid = RetimeWrapper_20_io_out; // @[MemInterfaceType.scala 311:132:@5935.4]
  assign io_in_x440_argOut_port_0_bits = {{48'd0}, x524_0_number}; // @[MemInterfaceType.scala 311:109:@5934.4]
  assign io_in_x436_argOut_port_0_valid = RetimeWrapper_16_io_out; // @[MemInterfaceType.scala 311:132:@5856.4]
  assign io_in_x436_argOut_port_0_bits = {{48'd0}, x513_0_number}; // @[MemInterfaceType.scala 311:109:@5855.4]
  assign io_in_x421_argOut_port_0_valid = RetimeWrapper_1_io_out; // @[MemInterfaceType.scala 311:132:@5553.4]
  assign io_in_x421_argOut_port_0_bits = {{48'd0}, x469_1_number}; // @[MemInterfaceType.scala 311:109:@5552.4]
  assign io_in_x448_argOut_port_0_valid = RetimeWrapper_28_io_out; // @[MemInterfaceType.scala 311:132:@6093.4]
  assign io_in_x448_argOut_port_0_bits = {{48'd0}, x546_0_number}; // @[MemInterfaceType.scala 311:109:@6092.4]
  assign io_in_x443_argOut_port_0_valid = RetimeWrapper_23_io_out; // @[MemInterfaceType.scala 311:132:@5974.4]
  assign io_in_x443_argOut_port_0_bits = {{48'd0}, x524_3_number}; // @[MemInterfaceType.scala 311:109:@5973.4]
  assign io_in_x428_argOut_port_0_valid = RetimeWrapper_8_io_out; // @[MemInterfaceType.scala 311:132:@5698.4]
  assign io_in_x428_argOut_port_0_bits = {{48'd0}, x491_0_number}; // @[MemInterfaceType.scala 311:109:@5697.4]
  assign io_in_x452_a_0_rPort_7_en_0 = _T_1262 & _T_1266; // @[MemInterfaceType.scala 110:79:@5594.4]
  assign io_in_x452_a_0_rPort_6_en_0 = _T_1262 & _T_1266; // @[MemInterfaceType.scala 110:79:@6068.4]
  assign io_in_x452_a_0_rPort_5_en_0 = _T_1262 & _T_1266; // @[MemInterfaceType.scala 110:79:@5673.4]
  assign io_in_x452_a_0_rPort_4_en_0 = _T_1262 & _T_1266; // @[MemInterfaceType.scala 110:79:@5910.4]
  assign io_in_x452_a_0_rPort_3_en_0 = _T_1262 & _T_1266; // @[MemInterfaceType.scala 110:79:@5515.4]
  assign io_in_x452_a_0_rPort_2_en_0 = _T_1262 & _T_1266; // @[MemInterfaceType.scala 110:79:@5752.4]
  assign io_in_x452_a_0_rPort_1_en_0 = _T_1262 & _T_1266; // @[MemInterfaceType.scala 110:79:@5989.4]
  assign io_in_x452_a_0_rPort_0_en_0 = _T_1262 & _T_1266; // @[MemInterfaceType.scala 110:79:@5831.4]
  assign io_in_x439_argOut_port_0_valid = RetimeWrapper_19_io_out; // @[MemInterfaceType.scala 311:132:@5895.4]
  assign io_in_x439_argOut_port_0_bits = {{48'd0}, x513_3_number}; // @[MemInterfaceType.scala 311:109:@5894.4]
  assign io_in_x424_argOut_port_0_valid = RetimeWrapper_4_io_out; // @[MemInterfaceType.scala 311:132:@5619.4]
  assign io_in_x424_argOut_port_0_bits = {{48'd0}, x480_0_number}; // @[MemInterfaceType.scala 311:109:@5618.4]
  assign io_in_x429_argOut_port_0_valid = RetimeWrapper_9_io_out; // @[MemInterfaceType.scala 311:132:@5711.4]
  assign io_in_x429_argOut_port_0_bits = {{48'd0}, x491_1_number}; // @[MemInterfaceType.scala 311:109:@5710.4]
  assign io_in_x435_argOut_port_0_valid = RetimeWrapper_15_io_out; // @[MemInterfaceType.scala 311:132:@5816.4]
  assign io_in_x435_argOut_port_0_bits = {{48'd0}, x502_3_number}; // @[MemInterfaceType.scala 311:109:@5815.4]
  assign io_in_x420_argOut_port_0_valid = RetimeWrapper_io_out; // @[MemInterfaceType.scala 311:132:@5540.4]
  assign io_in_x420_argOut_port_0_bits = {{48'd0}, x469_0_number}; // @[MemInterfaceType.scala 311:109:@5539.4]
  assign io_in_x425_argOut_port_0_valid = RetimeWrapper_5_io_out; // @[MemInterfaceType.scala 311:132:@5632.4]
  assign io_in_x425_argOut_port_0_bits = {{48'd0}, x480_1_number}; // @[MemInterfaceType.scala 311:109:@5631.4]
  assign io_in_x430_argOut_port_0_valid = RetimeWrapper_10_io_out; // @[MemInterfaceType.scala 311:132:@5724.4]
  assign io_in_x430_argOut_port_0_bits = {{48'd0}, x491_2_number}; // @[MemInterfaceType.scala 311:109:@5723.4]
  assign io_in_x444_argOut_port_0_valid = RetimeWrapper_24_io_out; // @[MemInterfaceType.scala 311:132:@6014.4]
  assign io_in_x444_argOut_port_0_bits = {{48'd0}, x535_0_number}; // @[MemInterfaceType.scala 311:109:@6013.4]
  assign io_in_x423_argOut_port_0_valid = RetimeWrapper_3_io_out; // @[MemInterfaceType.scala 311:132:@5579.4]
  assign io_in_x423_argOut_port_0_bits = {{48'd0}, x469_3_number}; // @[MemInterfaceType.scala 311:109:@5578.4]
  assign io_in_x445_argOut_port_0_valid = RetimeWrapper_25_io_out; // @[MemInterfaceType.scala 311:132:@6027.4]
  assign io_in_x445_argOut_port_0_bits = {{48'd0}, x535_1_number}; // @[MemInterfaceType.scala 311:109:@6026.4]
  assign io_in_x451_argOut_port_0_valid = RetimeWrapper_31_io_out; // @[MemInterfaceType.scala 311:132:@6132.4]
  assign io_in_x451_argOut_port_0_bits = {{48'd0}, x546_3_number}; // @[MemInterfaceType.scala 311:109:@6131.4]
  assign io_in_x434_argOut_port_0_valid = RetimeWrapper_14_io_out; // @[MemInterfaceType.scala 311:132:@5803.4]
  assign io_in_x434_argOut_port_0_bits = {{48'd0}, x502_2_number}; // @[MemInterfaceType.scala 311:109:@5802.4]
  assign io_in_x438_argOut_port_0_valid = RetimeWrapper_18_io_out; // @[MemInterfaceType.scala 311:132:@5882.4]
  assign io_in_x438_argOut_port_0_bits = {{48'd0}, x513_2_number}; // @[MemInterfaceType.scala 311:109:@5881.4]
  assign io_in_x431_argOut_port_0_valid = RetimeWrapper_11_io_out; // @[MemInterfaceType.scala 311:132:@5737.4]
  assign io_in_x431_argOut_port_0_bits = {{48'd0}, x491_3_number}; // @[MemInterfaceType.scala 311:109:@5736.4]
  assign io_in_x426_argOut_port_0_valid = RetimeWrapper_6_io_out; // @[MemInterfaceType.scala 311:132:@5645.4]
  assign io_in_x426_argOut_port_0_bits = {{48'd0}, x480_2_number}; // @[MemInterfaceType.scala 311:109:@5644.4]
  assign io_in_x441_argOut_port_0_valid = RetimeWrapper_21_io_out; // @[MemInterfaceType.scala 311:132:@5948.4]
  assign io_in_x441_argOut_port_0_bits = {{48'd0}, x524_1_number}; // @[MemInterfaceType.scala 311:109:@5947.4]
  assign io_in_x446_argOut_port_0_valid = RetimeWrapper_26_io_out; // @[MemInterfaceType.scala 311:132:@6040.4]
  assign io_in_x446_argOut_port_0_bits = {{48'd0}, x535_2_number}; // @[MemInterfaceType.scala 311:109:@6039.4]
  assign io_in_x450_argOut_port_0_valid = RetimeWrapper_30_io_out; // @[MemInterfaceType.scala 311:132:@6119.4]
  assign io_in_x450_argOut_port_0_bits = {{48'd0}, x546_2_number}; // @[MemInterfaceType.scala 311:109:@6118.4]
  assign io_in_x433_argOut_port_0_valid = RetimeWrapper_13_io_out; // @[MemInterfaceType.scala 311:132:@5790.4]
  assign io_in_x433_argOut_port_0_bits = {{48'd0}, x502_1_number}; // @[MemInterfaceType.scala 311:109:@5789.4]
  assign io_in_x447_argOut_port_0_valid = RetimeWrapper_27_io_out; // @[MemInterfaceType.scala 311:132:@6053.4]
  assign io_in_x447_argOut_port_0_bits = {{48'd0}, x535_3_number}; // @[MemInterfaceType.scala 311:109:@6052.4]
  assign io_in_x432_argOut_port_0_valid = RetimeWrapper_12_io_out; // @[MemInterfaceType.scala 311:132:@5777.4]
  assign io_in_x432_argOut_port_0_bits = {{48'd0}, x502_0_number}; // @[MemInterfaceType.scala 311:109:@5776.4]
  assign io_in_x422_argOut_port_0_valid = RetimeWrapper_2_io_out; // @[MemInterfaceType.scala 311:132:@5566.4]
  assign io_in_x422_argOut_port_0_bits = {{48'd0}, x469_2_number}; // @[MemInterfaceType.scala 311:109:@5565.4]
  assign io_in_x437_argOut_port_0_valid = RetimeWrapper_17_io_out; // @[MemInterfaceType.scala 311:132:@5869.4]
  assign io_in_x437_argOut_port_0_bits = {{48'd0}, x513_1_number}; // @[MemInterfaceType.scala 311:109:@5868.4]
  assign io_in_x427_argOut_port_0_valid = RetimeWrapper_7_io_out; // @[MemInterfaceType.scala 311:132:@5658.4]
  assign io_in_x427_argOut_port_0_bits = {{48'd0}, x480_3_number}; // @[MemInterfaceType.scala 311:109:@5657.4]
  assign io_in_x442_argOut_port_0_valid = RetimeWrapper_22_io_out; // @[MemInterfaceType.scala 311:132:@5961.4]
  assign io_in_x442_argOut_port_0_bits = {{48'd0}, x524_2_number}; // @[MemInterfaceType.scala 311:109:@5960.4]
  assign RetimeWrapper_clock = clock; // @[:@5532.4]
  assign RetimeWrapper_reset = reset; // @[:@5533.4]
  assign RetimeWrapper_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@5534.4]
  assign RetimeWrapper_1_clock = clock; // @[:@5545.4]
  assign RetimeWrapper_1_reset = reset; // @[:@5546.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@5547.4]
  assign RetimeWrapper_2_clock = clock; // @[:@5558.4]
  assign RetimeWrapper_2_reset = reset; // @[:@5559.4]
  assign RetimeWrapper_2_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@5560.4]
  assign RetimeWrapper_3_clock = clock; // @[:@5571.4]
  assign RetimeWrapper_3_reset = reset; // @[:@5572.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@5573.4]
  assign RetimeWrapper_4_clock = clock; // @[:@5611.4]
  assign RetimeWrapper_4_reset = reset; // @[:@5612.4]
  assign RetimeWrapper_4_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@5613.4]
  assign RetimeWrapper_5_clock = clock; // @[:@5624.4]
  assign RetimeWrapper_5_reset = reset; // @[:@5625.4]
  assign RetimeWrapper_5_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@5626.4]
  assign RetimeWrapper_6_clock = clock; // @[:@5637.4]
  assign RetimeWrapper_6_reset = reset; // @[:@5638.4]
  assign RetimeWrapper_6_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@5639.4]
  assign RetimeWrapper_7_clock = clock; // @[:@5650.4]
  assign RetimeWrapper_7_reset = reset; // @[:@5651.4]
  assign RetimeWrapper_7_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@5652.4]
  assign RetimeWrapper_8_clock = clock; // @[:@5690.4]
  assign RetimeWrapper_8_reset = reset; // @[:@5691.4]
  assign RetimeWrapper_8_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@5692.4]
  assign RetimeWrapper_9_clock = clock; // @[:@5703.4]
  assign RetimeWrapper_9_reset = reset; // @[:@5704.4]
  assign RetimeWrapper_9_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@5705.4]
  assign RetimeWrapper_10_clock = clock; // @[:@5716.4]
  assign RetimeWrapper_10_reset = reset; // @[:@5717.4]
  assign RetimeWrapper_10_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@5718.4]
  assign RetimeWrapper_11_clock = clock; // @[:@5729.4]
  assign RetimeWrapper_11_reset = reset; // @[:@5730.4]
  assign RetimeWrapper_11_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@5731.4]
  assign RetimeWrapper_12_clock = clock; // @[:@5769.4]
  assign RetimeWrapper_12_reset = reset; // @[:@5770.4]
  assign RetimeWrapper_12_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@5771.4]
  assign RetimeWrapper_13_clock = clock; // @[:@5782.4]
  assign RetimeWrapper_13_reset = reset; // @[:@5783.4]
  assign RetimeWrapper_13_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@5784.4]
  assign RetimeWrapper_14_clock = clock; // @[:@5795.4]
  assign RetimeWrapper_14_reset = reset; // @[:@5796.4]
  assign RetimeWrapper_14_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@5797.4]
  assign RetimeWrapper_15_clock = clock; // @[:@5808.4]
  assign RetimeWrapper_15_reset = reset; // @[:@5809.4]
  assign RetimeWrapper_15_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@5810.4]
  assign RetimeWrapper_16_clock = clock; // @[:@5848.4]
  assign RetimeWrapper_16_reset = reset; // @[:@5849.4]
  assign RetimeWrapper_16_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@5850.4]
  assign RetimeWrapper_17_clock = clock; // @[:@5861.4]
  assign RetimeWrapper_17_reset = reset; // @[:@5862.4]
  assign RetimeWrapper_17_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@5863.4]
  assign RetimeWrapper_18_clock = clock; // @[:@5874.4]
  assign RetimeWrapper_18_reset = reset; // @[:@5875.4]
  assign RetimeWrapper_18_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@5876.4]
  assign RetimeWrapper_19_clock = clock; // @[:@5887.4]
  assign RetimeWrapper_19_reset = reset; // @[:@5888.4]
  assign RetimeWrapper_19_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@5889.4]
  assign RetimeWrapper_20_clock = clock; // @[:@5927.4]
  assign RetimeWrapper_20_reset = reset; // @[:@5928.4]
  assign RetimeWrapper_20_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@5929.4]
  assign RetimeWrapper_21_clock = clock; // @[:@5940.4]
  assign RetimeWrapper_21_reset = reset; // @[:@5941.4]
  assign RetimeWrapper_21_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@5942.4]
  assign RetimeWrapper_22_clock = clock; // @[:@5953.4]
  assign RetimeWrapper_22_reset = reset; // @[:@5954.4]
  assign RetimeWrapper_22_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@5955.4]
  assign RetimeWrapper_23_clock = clock; // @[:@5966.4]
  assign RetimeWrapper_23_reset = reset; // @[:@5967.4]
  assign RetimeWrapper_23_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@5968.4]
  assign RetimeWrapper_24_clock = clock; // @[:@6006.4]
  assign RetimeWrapper_24_reset = reset; // @[:@6007.4]
  assign RetimeWrapper_24_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@6008.4]
  assign RetimeWrapper_25_clock = clock; // @[:@6019.4]
  assign RetimeWrapper_25_reset = reset; // @[:@6020.4]
  assign RetimeWrapper_25_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@6021.4]
  assign RetimeWrapper_26_clock = clock; // @[:@6032.4]
  assign RetimeWrapper_26_reset = reset; // @[:@6033.4]
  assign RetimeWrapper_26_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@6034.4]
  assign RetimeWrapper_27_clock = clock; // @[:@6045.4]
  assign RetimeWrapper_27_reset = reset; // @[:@6046.4]
  assign RetimeWrapper_27_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@6047.4]
  assign RetimeWrapper_28_clock = clock; // @[:@6085.4]
  assign RetimeWrapper_28_reset = reset; // @[:@6086.4]
  assign RetimeWrapper_28_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@6087.4]
  assign RetimeWrapper_29_clock = clock; // @[:@6098.4]
  assign RetimeWrapper_29_reset = reset; // @[:@6099.4]
  assign RetimeWrapper_29_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@6100.4]
  assign RetimeWrapper_30_clock = clock; // @[:@6111.4]
  assign RetimeWrapper_30_reset = reset; // @[:@6112.4]
  assign RetimeWrapper_30_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@6113.4]
  assign RetimeWrapper_31_clock = clock; // @[:@6124.4]
  assign RetimeWrapper_31_reset = reset; // @[:@6125.4]
  assign RetimeWrapper_31_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@6126.4]
endmodule
module RootController_kernelRootController_concrete1( // @[:@6134.2]
  input          clock, // @[:@6135.4]
  input          reset, // @[:@6136.4]
  output         io_in_x449_argOut_port_0_valid, // @[:@6137.4]
  output [63:0]  io_in_x449_argOut_port_0_bits, // @[:@6137.4]
  output         io_in_x440_argOut_port_0_valid, // @[:@6137.4]
  output [63:0]  io_in_x440_argOut_port_0_bits, // @[:@6137.4]
  output         io_in_x436_argOut_port_0_valid, // @[:@6137.4]
  output [63:0]  io_in_x436_argOut_port_0_bits, // @[:@6137.4]
  output         io_in_x421_argOut_port_0_valid, // @[:@6137.4]
  output [63:0]  io_in_x421_argOut_port_0_bits, // @[:@6137.4]
  input          io_in_x416_TVALID, // @[:@6137.4]
  output         io_in_x416_TREADY, // @[:@6137.4]
  input  [255:0] io_in_x416_TDATA, // @[:@6137.4]
  output         io_in_x448_argOut_port_0_valid, // @[:@6137.4]
  output [63:0]  io_in_x448_argOut_port_0_bits, // @[:@6137.4]
  output         io_in_x443_argOut_port_0_valid, // @[:@6137.4]
  output [63:0]  io_in_x443_argOut_port_0_bits, // @[:@6137.4]
  output         io_in_x428_argOut_port_0_valid, // @[:@6137.4]
  output [63:0]  io_in_x428_argOut_port_0_bits, // @[:@6137.4]
  output         io_in_x439_argOut_port_0_valid, // @[:@6137.4]
  output [63:0]  io_in_x439_argOut_port_0_bits, // @[:@6137.4]
  output         io_in_x424_argOut_port_0_valid, // @[:@6137.4]
  output [63:0]  io_in_x424_argOut_port_0_bits, // @[:@6137.4]
  output         io_in_x429_argOut_port_0_valid, // @[:@6137.4]
  output [63:0]  io_in_x429_argOut_port_0_bits, // @[:@6137.4]
  output         io_in_x435_argOut_port_0_valid, // @[:@6137.4]
  output [63:0]  io_in_x435_argOut_port_0_bits, // @[:@6137.4]
  output         io_in_x420_argOut_port_0_valid, // @[:@6137.4]
  output [63:0]  io_in_x420_argOut_port_0_bits, // @[:@6137.4]
  output         io_in_x425_argOut_port_0_valid, // @[:@6137.4]
  output [63:0]  io_in_x425_argOut_port_0_bits, // @[:@6137.4]
  output         io_in_x430_argOut_port_0_valid, // @[:@6137.4]
  output [63:0]  io_in_x430_argOut_port_0_bits, // @[:@6137.4]
  output         io_in_x444_argOut_port_0_valid, // @[:@6137.4]
  output [63:0]  io_in_x444_argOut_port_0_bits, // @[:@6137.4]
  output         io_in_x423_argOut_port_0_valid, // @[:@6137.4]
  output [63:0]  io_in_x423_argOut_port_0_bits, // @[:@6137.4]
  output         io_in_x445_argOut_port_0_valid, // @[:@6137.4]
  output [63:0]  io_in_x445_argOut_port_0_bits, // @[:@6137.4]
  output         io_in_x451_argOut_port_0_valid, // @[:@6137.4]
  output [63:0]  io_in_x451_argOut_port_0_bits, // @[:@6137.4]
  output         io_in_x434_argOut_port_0_valid, // @[:@6137.4]
  output [63:0]  io_in_x434_argOut_port_0_bits, // @[:@6137.4]
  output         io_in_x438_argOut_port_0_valid, // @[:@6137.4]
  output [63:0]  io_in_x438_argOut_port_0_bits, // @[:@6137.4]
  output         io_in_x431_argOut_port_0_valid, // @[:@6137.4]
  output [63:0]  io_in_x431_argOut_port_0_bits, // @[:@6137.4]
  output         io_in_x426_argOut_port_0_valid, // @[:@6137.4]
  output [63:0]  io_in_x426_argOut_port_0_bits, // @[:@6137.4]
  output         io_in_x441_argOut_port_0_valid, // @[:@6137.4]
  output [63:0]  io_in_x441_argOut_port_0_bits, // @[:@6137.4]
  output         io_in_x446_argOut_port_0_valid, // @[:@6137.4]
  output [63:0]  io_in_x446_argOut_port_0_bits, // @[:@6137.4]
  output         io_in_x450_argOut_port_0_valid, // @[:@6137.4]
  output [63:0]  io_in_x450_argOut_port_0_bits, // @[:@6137.4]
  output         io_in_x433_argOut_port_0_valid, // @[:@6137.4]
  output [63:0]  io_in_x433_argOut_port_0_bits, // @[:@6137.4]
  output         io_in_x447_argOut_port_0_valid, // @[:@6137.4]
  output [63:0]  io_in_x447_argOut_port_0_bits, // @[:@6137.4]
  output         io_in_x432_argOut_port_0_valid, // @[:@6137.4]
  output [63:0]  io_in_x432_argOut_port_0_bits, // @[:@6137.4]
  output         io_in_x422_argOut_port_0_valid, // @[:@6137.4]
  output [63:0]  io_in_x422_argOut_port_0_bits, // @[:@6137.4]
  output         io_in_x437_argOut_port_0_valid, // @[:@6137.4]
  output [63:0]  io_in_x437_argOut_port_0_bits, // @[:@6137.4]
  output         io_in_x427_argOut_port_0_valid, // @[:@6137.4]
  output [63:0]  io_in_x427_argOut_port_0_bits, // @[:@6137.4]
  output         io_in_x442_argOut_port_0_valid, // @[:@6137.4]
  output [63:0]  io_in_x442_argOut_port_0_bits, // @[:@6137.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@6137.4]
  input          io_sigsIn_smEnableOuts_1, // @[:@6137.4]
  input          io_sigsIn_smChildAcks_0, // @[:@6137.4]
  input          io_sigsIn_smChildAcks_1, // @[:@6137.4]
  output         io_sigsOut_smDoneIn_0, // @[:@6137.4]
  output         io_sigsOut_smDoneIn_1, // @[:@6137.4]
  input          io_rr // @[:@6137.4]
);
  wire  x452_a_0_clock; // @[m_x452_a_0.scala 34:17:@6277.4]
  wire  x452_a_0_reset; // @[m_x452_a_0.scala 34:17:@6277.4]
  wire  x452_a_0_io_rPort_7_en_0; // @[m_x452_a_0.scala 34:17:@6277.4]
  wire [63:0] x452_a_0_io_rPort_7_output_0; // @[m_x452_a_0.scala 34:17:@6277.4]
  wire  x452_a_0_io_rPort_6_en_0; // @[m_x452_a_0.scala 34:17:@6277.4]
  wire [63:0] x452_a_0_io_rPort_6_output_0; // @[m_x452_a_0.scala 34:17:@6277.4]
  wire  x452_a_0_io_rPort_5_en_0; // @[m_x452_a_0.scala 34:17:@6277.4]
  wire [63:0] x452_a_0_io_rPort_5_output_0; // @[m_x452_a_0.scala 34:17:@6277.4]
  wire  x452_a_0_io_rPort_4_en_0; // @[m_x452_a_0.scala 34:17:@6277.4]
  wire [63:0] x452_a_0_io_rPort_4_output_0; // @[m_x452_a_0.scala 34:17:@6277.4]
  wire  x452_a_0_io_rPort_3_en_0; // @[m_x452_a_0.scala 34:17:@6277.4]
  wire [63:0] x452_a_0_io_rPort_3_output_0; // @[m_x452_a_0.scala 34:17:@6277.4]
  wire  x452_a_0_io_rPort_2_en_0; // @[m_x452_a_0.scala 34:17:@6277.4]
  wire [63:0] x452_a_0_io_rPort_2_output_0; // @[m_x452_a_0.scala 34:17:@6277.4]
  wire  x452_a_0_io_rPort_1_en_0; // @[m_x452_a_0.scala 34:17:@6277.4]
  wire [63:0] x452_a_0_io_rPort_1_output_0; // @[m_x452_a_0.scala 34:17:@6277.4]
  wire  x452_a_0_io_rPort_0_en_0; // @[m_x452_a_0.scala 34:17:@6277.4]
  wire [63:0] x452_a_0_io_rPort_0_output_0; // @[m_x452_a_0.scala 34:17:@6277.4]
  wire [3:0] x452_a_0_io_wPort_0_banks_0; // @[m_x452_a_0.scala 34:17:@6277.4]
  wire [2:0] x452_a_0_io_wPort_0_ofs_0; // @[m_x452_a_0.scala 34:17:@6277.4]
  wire [63:0] x452_a_0_io_wPort_0_data_0; // @[m_x452_a_0.scala 34:17:@6277.4]
  wire  x452_a_0_io_wPort_0_en_0; // @[m_x452_a_0.scala 34:17:@6277.4]
  wire  x466_outr_UnitPipe_sm_clock; // @[sm_x466_outr_UnitPipe.scala 33:18:@6364.4]
  wire  x466_outr_UnitPipe_sm_reset; // @[sm_x466_outr_UnitPipe.scala 33:18:@6364.4]
  wire  x466_outr_UnitPipe_sm_io_enable; // @[sm_x466_outr_UnitPipe.scala 33:18:@6364.4]
  wire  x466_outr_UnitPipe_sm_io_done; // @[sm_x466_outr_UnitPipe.scala 33:18:@6364.4]
  wire  x466_outr_UnitPipe_sm_io_parentAck; // @[sm_x466_outr_UnitPipe.scala 33:18:@6364.4]
  wire  x466_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x466_outr_UnitPipe.scala 33:18:@6364.4]
  wire  x466_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x466_outr_UnitPipe.scala 33:18:@6364.4]
  wire  x466_outr_UnitPipe_sm_io_childAck_0; // @[sm_x466_outr_UnitPipe.scala 33:18:@6364.4]
  wire  x466_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x466_outr_UnitPipe.scala 33:18:@6364.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@6416.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@6416.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@6416.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@6416.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@6416.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@6424.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@6424.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@6424.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@6424.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@6424.4]
  wire  x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_clock; // @[sm_x466_outr_UnitPipe.scala 75:24:@6451.4]
  wire  x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_reset; // @[sm_x466_outr_UnitPipe.scala 75:24:@6451.4]
  wire  x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_in_x416_TVALID; // @[sm_x466_outr_UnitPipe.scala 75:24:@6451.4]
  wire  x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_in_x416_TREADY; // @[sm_x466_outr_UnitPipe.scala 75:24:@6451.4]
  wire [255:0] x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_in_x416_TDATA; // @[sm_x466_outr_UnitPipe.scala 75:24:@6451.4]
  wire [3:0] x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_in_x452_a_0_wPort_0_banks_0; // @[sm_x466_outr_UnitPipe.scala 75:24:@6451.4]
  wire [2:0] x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_in_x452_a_0_wPort_0_ofs_0; // @[sm_x466_outr_UnitPipe.scala 75:24:@6451.4]
  wire [63:0] x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_in_x452_a_0_wPort_0_data_0; // @[sm_x466_outr_UnitPipe.scala 75:24:@6451.4]
  wire  x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_in_x452_a_0_wPort_0_en_0; // @[sm_x466_outr_UnitPipe.scala 75:24:@6451.4]
  wire  x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x466_outr_UnitPipe.scala 75:24:@6451.4]
  wire  x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x466_outr_UnitPipe.scala 75:24:@6451.4]
  wire  x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x466_outr_UnitPipe.scala 75:24:@6451.4]
  wire  x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x466_outr_UnitPipe.scala 75:24:@6451.4]
  wire  x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_rr; // @[sm_x466_outr_UnitPipe.scala 75:24:@6451.4]
  wire  x555_inr_UnitPipe_sm_clock; // @[sm_x555_inr_UnitPipe.scala 33:18:@6613.4]
  wire  x555_inr_UnitPipe_sm_reset; // @[sm_x555_inr_UnitPipe.scala 33:18:@6613.4]
  wire  x555_inr_UnitPipe_sm_io_enable; // @[sm_x555_inr_UnitPipe.scala 33:18:@6613.4]
  wire  x555_inr_UnitPipe_sm_io_done; // @[sm_x555_inr_UnitPipe.scala 33:18:@6613.4]
  wire  x555_inr_UnitPipe_sm_io_ctrDone; // @[sm_x555_inr_UnitPipe.scala 33:18:@6613.4]
  wire  x555_inr_UnitPipe_sm_io_datapathEn; // @[sm_x555_inr_UnitPipe.scala 33:18:@6613.4]
  wire  x555_inr_UnitPipe_sm_io_ctrInc; // @[sm_x555_inr_UnitPipe.scala 33:18:@6613.4]
  wire  x555_inr_UnitPipe_sm_io_parentAck; // @[sm_x555_inr_UnitPipe.scala 33:18:@6613.4]
  wire  x555_inr_UnitPipe_sm_io_break; // @[sm_x555_inr_UnitPipe.scala 33:18:@6613.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@6670.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@6670.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@6670.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@6670.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@6670.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@6678.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@6678.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@6678.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@6678.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@6678.4]
  wire  x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_clock; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire  x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_reset; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire  x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x449_argOut_port_0_valid; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire [63:0] x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x449_argOut_port_0_bits; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire  x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x440_argOut_port_0_valid; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire [63:0] x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x440_argOut_port_0_bits; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire  x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x436_argOut_port_0_valid; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire [63:0] x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x436_argOut_port_0_bits; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire  x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x421_argOut_port_0_valid; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire [63:0] x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x421_argOut_port_0_bits; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire  x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x448_argOut_port_0_valid; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire [63:0] x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x448_argOut_port_0_bits; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire  x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x443_argOut_port_0_valid; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire [63:0] x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x443_argOut_port_0_bits; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire  x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x428_argOut_port_0_valid; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire [63:0] x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x428_argOut_port_0_bits; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire  x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x452_a_0_rPort_7_en_0; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire [63:0] x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x452_a_0_rPort_7_output_0; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire  x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x452_a_0_rPort_6_en_0; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire [63:0] x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x452_a_0_rPort_6_output_0; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire  x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x452_a_0_rPort_5_en_0; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire [63:0] x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x452_a_0_rPort_5_output_0; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire  x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x452_a_0_rPort_4_en_0; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire [63:0] x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x452_a_0_rPort_4_output_0; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire  x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x452_a_0_rPort_3_en_0; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire [63:0] x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x452_a_0_rPort_3_output_0; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire  x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x452_a_0_rPort_2_en_0; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire [63:0] x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x452_a_0_rPort_2_output_0; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire  x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x452_a_0_rPort_1_en_0; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire [63:0] x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x452_a_0_rPort_1_output_0; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire  x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x452_a_0_rPort_0_en_0; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire [63:0] x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x452_a_0_rPort_0_output_0; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire  x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x439_argOut_port_0_valid; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire [63:0] x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x439_argOut_port_0_bits; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire  x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x424_argOut_port_0_valid; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire [63:0] x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x424_argOut_port_0_bits; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire  x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x429_argOut_port_0_valid; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire [63:0] x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x429_argOut_port_0_bits; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire  x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x435_argOut_port_0_valid; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire [63:0] x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x435_argOut_port_0_bits; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire  x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x420_argOut_port_0_valid; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire [63:0] x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x420_argOut_port_0_bits; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire  x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x425_argOut_port_0_valid; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire [63:0] x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x425_argOut_port_0_bits; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire  x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x430_argOut_port_0_valid; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire [63:0] x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x430_argOut_port_0_bits; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire  x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x444_argOut_port_0_valid; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire [63:0] x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x444_argOut_port_0_bits; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire  x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x423_argOut_port_0_valid; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire [63:0] x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x423_argOut_port_0_bits; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire  x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x445_argOut_port_0_valid; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire [63:0] x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x445_argOut_port_0_bits; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire  x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x451_argOut_port_0_valid; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire [63:0] x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x451_argOut_port_0_bits; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire  x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x434_argOut_port_0_valid; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire [63:0] x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x434_argOut_port_0_bits; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire  x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x438_argOut_port_0_valid; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire [63:0] x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x438_argOut_port_0_bits; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire  x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x431_argOut_port_0_valid; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire [63:0] x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x431_argOut_port_0_bits; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire  x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x426_argOut_port_0_valid; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire [63:0] x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x426_argOut_port_0_bits; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire  x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x441_argOut_port_0_valid; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire [63:0] x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x441_argOut_port_0_bits; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire  x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x446_argOut_port_0_valid; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire [63:0] x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x446_argOut_port_0_bits; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire  x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x450_argOut_port_0_valid; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire [63:0] x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x450_argOut_port_0_bits; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire  x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x433_argOut_port_0_valid; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire [63:0] x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x433_argOut_port_0_bits; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire  x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x447_argOut_port_0_valid; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire [63:0] x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x447_argOut_port_0_bits; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire  x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x432_argOut_port_0_valid; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire [63:0] x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x432_argOut_port_0_bits; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire  x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x422_argOut_port_0_valid; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire [63:0] x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x422_argOut_port_0_bits; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire  x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x437_argOut_port_0_valid; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire [63:0] x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x437_argOut_port_0_bits; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire  x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x427_argOut_port_0_valid; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire [63:0] x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x427_argOut_port_0_bits; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire  x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x442_argOut_port_0_valid; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire [63:0] x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x442_argOut_port_0_bits; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire  x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_sigsIn_datapathEn; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire  x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_sigsIn_break; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire  x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_rr; // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
  wire  _T_843; // @[package.scala 96:25:@6421.4 package.scala 96:25:@6422.4]
  wire  _T_849; // @[package.scala 96:25:@6429.4 package.scala 96:25:@6430.4]
  wire  _T_852; // @[SpatialBlocks.scala 110:93:@6432.4]
  wire  _T_918; // @[package.scala 100:49:@6641.4]
  reg  _T_921; // @[package.scala 48:56:@6642.4]
  reg [31:0] _RAND_0;
  wire  _T_935; // @[package.scala 96:25:@6675.4 package.scala 96:25:@6676.4]
  wire  _T_941; // @[package.scala 96:25:@6683.4 package.scala 96:25:@6684.4]
  wire  _T_944; // @[SpatialBlocks.scala 110:93:@6686.4]
  x452_a_0 x452_a_0 ( // @[m_x452_a_0.scala 34:17:@6277.4]
    .clock(x452_a_0_clock),
    .reset(x452_a_0_reset),
    .io_rPort_7_en_0(x452_a_0_io_rPort_7_en_0),
    .io_rPort_7_output_0(x452_a_0_io_rPort_7_output_0),
    .io_rPort_6_en_0(x452_a_0_io_rPort_6_en_0),
    .io_rPort_6_output_0(x452_a_0_io_rPort_6_output_0),
    .io_rPort_5_en_0(x452_a_0_io_rPort_5_en_0),
    .io_rPort_5_output_0(x452_a_0_io_rPort_5_output_0),
    .io_rPort_4_en_0(x452_a_0_io_rPort_4_en_0),
    .io_rPort_4_output_0(x452_a_0_io_rPort_4_output_0),
    .io_rPort_3_en_0(x452_a_0_io_rPort_3_en_0),
    .io_rPort_3_output_0(x452_a_0_io_rPort_3_output_0),
    .io_rPort_2_en_0(x452_a_0_io_rPort_2_en_0),
    .io_rPort_2_output_0(x452_a_0_io_rPort_2_output_0),
    .io_rPort_1_en_0(x452_a_0_io_rPort_1_en_0),
    .io_rPort_1_output_0(x452_a_0_io_rPort_1_output_0),
    .io_rPort_0_en_0(x452_a_0_io_rPort_0_en_0),
    .io_rPort_0_output_0(x452_a_0_io_rPort_0_output_0),
    .io_wPort_0_banks_0(x452_a_0_io_wPort_0_banks_0),
    .io_wPort_0_ofs_0(x452_a_0_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x452_a_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x452_a_0_io_wPort_0_en_0)
  );
  x466_outr_UnitPipe_sm x466_outr_UnitPipe_sm ( // @[sm_x466_outr_UnitPipe.scala 33:18:@6364.4]
    .clock(x466_outr_UnitPipe_sm_clock),
    .reset(x466_outr_UnitPipe_sm_reset),
    .io_enable(x466_outr_UnitPipe_sm_io_enable),
    .io_done(x466_outr_UnitPipe_sm_io_done),
    .io_parentAck(x466_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x466_outr_UnitPipe_sm_io_doneIn_0),
    .io_enableOut_0(x466_outr_UnitPipe_sm_io_enableOut_0),
    .io_childAck_0(x466_outr_UnitPipe_sm_io_childAck_0),
    .io_ctrCopyDone_0(x466_outr_UnitPipe_sm_io_ctrCopyDone_0)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@6416.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@6424.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1 x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1 ( // @[sm_x466_outr_UnitPipe.scala 75:24:@6451.4]
    .clock(x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_clock),
    .reset(x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_reset),
    .io_in_x416_TVALID(x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_in_x416_TVALID),
    .io_in_x416_TREADY(x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_in_x416_TREADY),
    .io_in_x416_TDATA(x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_in_x416_TDATA),
    .io_in_x452_a_0_wPort_0_banks_0(x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_in_x452_a_0_wPort_0_banks_0),
    .io_in_x452_a_0_wPort_0_ofs_0(x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_in_x452_a_0_wPort_0_ofs_0),
    .io_in_x452_a_0_wPort_0_data_0(x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_in_x452_a_0_wPort_0_data_0),
    .io_in_x452_a_0_wPort_0_en_0(x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_in_x452_a_0_wPort_0_en_0),
    .io_sigsIn_smEnableOuts_0(x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smCtrCopyDone_0(x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_rr(x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_rr)
  );
  x555_inr_UnitPipe_sm x555_inr_UnitPipe_sm ( // @[sm_x555_inr_UnitPipe.scala 33:18:@6613.4]
    .clock(x555_inr_UnitPipe_sm_clock),
    .reset(x555_inr_UnitPipe_sm_reset),
    .io_enable(x555_inr_UnitPipe_sm_io_enable),
    .io_done(x555_inr_UnitPipe_sm_io_done),
    .io_ctrDone(x555_inr_UnitPipe_sm_io_ctrDone),
    .io_datapathEn(x555_inr_UnitPipe_sm_io_datapathEn),
    .io_ctrInc(x555_inr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x555_inr_UnitPipe_sm_io_parentAck),
    .io_break(x555_inr_UnitPipe_sm_io_break)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@6670.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@6678.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1 x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1 ( // @[sm_x555_inr_UnitPipe.scala 398:24:@6704.4]
    .clock(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_clock),
    .reset(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_reset),
    .io_in_x449_argOut_port_0_valid(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x449_argOut_port_0_valid),
    .io_in_x449_argOut_port_0_bits(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x449_argOut_port_0_bits),
    .io_in_x440_argOut_port_0_valid(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x440_argOut_port_0_valid),
    .io_in_x440_argOut_port_0_bits(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x440_argOut_port_0_bits),
    .io_in_x436_argOut_port_0_valid(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x436_argOut_port_0_valid),
    .io_in_x436_argOut_port_0_bits(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x436_argOut_port_0_bits),
    .io_in_x421_argOut_port_0_valid(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x421_argOut_port_0_valid),
    .io_in_x421_argOut_port_0_bits(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x421_argOut_port_0_bits),
    .io_in_x448_argOut_port_0_valid(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x448_argOut_port_0_valid),
    .io_in_x448_argOut_port_0_bits(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x448_argOut_port_0_bits),
    .io_in_x443_argOut_port_0_valid(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x443_argOut_port_0_valid),
    .io_in_x443_argOut_port_0_bits(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x443_argOut_port_0_bits),
    .io_in_x428_argOut_port_0_valid(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x428_argOut_port_0_valid),
    .io_in_x428_argOut_port_0_bits(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x428_argOut_port_0_bits),
    .io_in_x452_a_0_rPort_7_en_0(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x452_a_0_rPort_7_en_0),
    .io_in_x452_a_0_rPort_7_output_0(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x452_a_0_rPort_7_output_0),
    .io_in_x452_a_0_rPort_6_en_0(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x452_a_0_rPort_6_en_0),
    .io_in_x452_a_0_rPort_6_output_0(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x452_a_0_rPort_6_output_0),
    .io_in_x452_a_0_rPort_5_en_0(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x452_a_0_rPort_5_en_0),
    .io_in_x452_a_0_rPort_5_output_0(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x452_a_0_rPort_5_output_0),
    .io_in_x452_a_0_rPort_4_en_0(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x452_a_0_rPort_4_en_0),
    .io_in_x452_a_0_rPort_4_output_0(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x452_a_0_rPort_4_output_0),
    .io_in_x452_a_0_rPort_3_en_0(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x452_a_0_rPort_3_en_0),
    .io_in_x452_a_0_rPort_3_output_0(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x452_a_0_rPort_3_output_0),
    .io_in_x452_a_0_rPort_2_en_0(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x452_a_0_rPort_2_en_0),
    .io_in_x452_a_0_rPort_2_output_0(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x452_a_0_rPort_2_output_0),
    .io_in_x452_a_0_rPort_1_en_0(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x452_a_0_rPort_1_en_0),
    .io_in_x452_a_0_rPort_1_output_0(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x452_a_0_rPort_1_output_0),
    .io_in_x452_a_0_rPort_0_en_0(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x452_a_0_rPort_0_en_0),
    .io_in_x452_a_0_rPort_0_output_0(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x452_a_0_rPort_0_output_0),
    .io_in_x439_argOut_port_0_valid(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x439_argOut_port_0_valid),
    .io_in_x439_argOut_port_0_bits(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x439_argOut_port_0_bits),
    .io_in_x424_argOut_port_0_valid(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x424_argOut_port_0_valid),
    .io_in_x424_argOut_port_0_bits(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x424_argOut_port_0_bits),
    .io_in_x429_argOut_port_0_valid(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x429_argOut_port_0_valid),
    .io_in_x429_argOut_port_0_bits(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x429_argOut_port_0_bits),
    .io_in_x435_argOut_port_0_valid(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x435_argOut_port_0_valid),
    .io_in_x435_argOut_port_0_bits(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x435_argOut_port_0_bits),
    .io_in_x420_argOut_port_0_valid(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x420_argOut_port_0_valid),
    .io_in_x420_argOut_port_0_bits(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x420_argOut_port_0_bits),
    .io_in_x425_argOut_port_0_valid(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x425_argOut_port_0_valid),
    .io_in_x425_argOut_port_0_bits(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x425_argOut_port_0_bits),
    .io_in_x430_argOut_port_0_valid(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x430_argOut_port_0_valid),
    .io_in_x430_argOut_port_0_bits(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x430_argOut_port_0_bits),
    .io_in_x444_argOut_port_0_valid(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x444_argOut_port_0_valid),
    .io_in_x444_argOut_port_0_bits(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x444_argOut_port_0_bits),
    .io_in_x423_argOut_port_0_valid(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x423_argOut_port_0_valid),
    .io_in_x423_argOut_port_0_bits(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x423_argOut_port_0_bits),
    .io_in_x445_argOut_port_0_valid(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x445_argOut_port_0_valid),
    .io_in_x445_argOut_port_0_bits(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x445_argOut_port_0_bits),
    .io_in_x451_argOut_port_0_valid(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x451_argOut_port_0_valid),
    .io_in_x451_argOut_port_0_bits(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x451_argOut_port_0_bits),
    .io_in_x434_argOut_port_0_valid(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x434_argOut_port_0_valid),
    .io_in_x434_argOut_port_0_bits(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x434_argOut_port_0_bits),
    .io_in_x438_argOut_port_0_valid(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x438_argOut_port_0_valid),
    .io_in_x438_argOut_port_0_bits(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x438_argOut_port_0_bits),
    .io_in_x431_argOut_port_0_valid(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x431_argOut_port_0_valid),
    .io_in_x431_argOut_port_0_bits(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x431_argOut_port_0_bits),
    .io_in_x426_argOut_port_0_valid(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x426_argOut_port_0_valid),
    .io_in_x426_argOut_port_0_bits(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x426_argOut_port_0_bits),
    .io_in_x441_argOut_port_0_valid(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x441_argOut_port_0_valid),
    .io_in_x441_argOut_port_0_bits(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x441_argOut_port_0_bits),
    .io_in_x446_argOut_port_0_valid(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x446_argOut_port_0_valid),
    .io_in_x446_argOut_port_0_bits(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x446_argOut_port_0_bits),
    .io_in_x450_argOut_port_0_valid(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x450_argOut_port_0_valid),
    .io_in_x450_argOut_port_0_bits(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x450_argOut_port_0_bits),
    .io_in_x433_argOut_port_0_valid(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x433_argOut_port_0_valid),
    .io_in_x433_argOut_port_0_bits(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x433_argOut_port_0_bits),
    .io_in_x447_argOut_port_0_valid(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x447_argOut_port_0_valid),
    .io_in_x447_argOut_port_0_bits(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x447_argOut_port_0_bits),
    .io_in_x432_argOut_port_0_valid(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x432_argOut_port_0_valid),
    .io_in_x432_argOut_port_0_bits(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x432_argOut_port_0_bits),
    .io_in_x422_argOut_port_0_valid(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x422_argOut_port_0_valid),
    .io_in_x422_argOut_port_0_bits(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x422_argOut_port_0_bits),
    .io_in_x437_argOut_port_0_valid(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x437_argOut_port_0_valid),
    .io_in_x437_argOut_port_0_bits(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x437_argOut_port_0_bits),
    .io_in_x427_argOut_port_0_valid(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x427_argOut_port_0_valid),
    .io_in_x427_argOut_port_0_bits(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x427_argOut_port_0_bits),
    .io_in_x442_argOut_port_0_valid(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x442_argOut_port_0_valid),
    .io_in_x442_argOut_port_0_bits(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x442_argOut_port_0_bits),
    .io_sigsIn_datapathEn(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_sigsIn_break),
    .io_rr(x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_rr)
  );
  assign _T_843 = RetimeWrapper_io_out; // @[package.scala 96:25:@6421.4 package.scala 96:25:@6422.4]
  assign _T_849 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@6429.4 package.scala 96:25:@6430.4]
  assign _T_852 = ~ _T_849; // @[SpatialBlocks.scala 110:93:@6432.4]
  assign _T_918 = x555_inr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@6641.4]
  assign _T_935 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@6675.4 package.scala 96:25:@6676.4]
  assign _T_941 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@6683.4 package.scala 96:25:@6684.4]
  assign _T_944 = ~ _T_941; // @[SpatialBlocks.scala 110:93:@6686.4]
  assign io_in_x449_argOut_port_0_valid = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x449_argOut_port_0_valid; // @[MemInterfaceType.scala 317:38:@6911.4]
  assign io_in_x449_argOut_port_0_bits = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x449_argOut_port_0_bits; // @[MemInterfaceType.scala 317:38:@6910.4]
  assign io_in_x440_argOut_port_0_valid = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x440_argOut_port_0_valid; // @[MemInterfaceType.scala 317:38:@6916.4]
  assign io_in_x440_argOut_port_0_bits = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x440_argOut_port_0_bits; // @[MemInterfaceType.scala 317:38:@6915.4]
  assign io_in_x436_argOut_port_0_valid = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x436_argOut_port_0_valid; // @[MemInterfaceType.scala 317:38:@6921.4]
  assign io_in_x436_argOut_port_0_bits = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x436_argOut_port_0_bits; // @[MemInterfaceType.scala 317:38:@6920.4]
  assign io_in_x421_argOut_port_0_valid = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x421_argOut_port_0_valid; // @[MemInterfaceType.scala 317:38:@6926.4]
  assign io_in_x421_argOut_port_0_bits = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x421_argOut_port_0_bits; // @[MemInterfaceType.scala 317:38:@6925.4]
  assign io_in_x416_TREADY = x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_in_x416_TREADY; // @[sm_x466_outr_UnitPipe.scala 49:23:@6543.4]
  assign io_in_x448_argOut_port_0_valid = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x448_argOut_port_0_valid; // @[MemInterfaceType.scala 317:38:@6931.4]
  assign io_in_x448_argOut_port_0_bits = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x448_argOut_port_0_bits; // @[MemInterfaceType.scala 317:38:@6930.4]
  assign io_in_x443_argOut_port_0_valid = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x443_argOut_port_0_valid; // @[MemInterfaceType.scala 317:38:@6936.4]
  assign io_in_x443_argOut_port_0_bits = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x443_argOut_port_0_bits; // @[MemInterfaceType.scala 317:38:@6935.4]
  assign io_in_x428_argOut_port_0_valid = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x428_argOut_port_0_valid; // @[MemInterfaceType.scala 317:38:@6941.4]
  assign io_in_x428_argOut_port_0_bits = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x428_argOut_port_0_bits; // @[MemInterfaceType.scala 317:38:@6940.4]
  assign io_in_x439_argOut_port_0_valid = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x439_argOut_port_0_valid; // @[MemInterfaceType.scala 317:38:@6986.4]
  assign io_in_x439_argOut_port_0_bits = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x439_argOut_port_0_bits; // @[MemInterfaceType.scala 317:38:@6985.4]
  assign io_in_x424_argOut_port_0_valid = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x424_argOut_port_0_valid; // @[MemInterfaceType.scala 317:38:@6991.4]
  assign io_in_x424_argOut_port_0_bits = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x424_argOut_port_0_bits; // @[MemInterfaceType.scala 317:38:@6990.4]
  assign io_in_x429_argOut_port_0_valid = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x429_argOut_port_0_valid; // @[MemInterfaceType.scala 317:38:@6996.4]
  assign io_in_x429_argOut_port_0_bits = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x429_argOut_port_0_bits; // @[MemInterfaceType.scala 317:38:@6995.4]
  assign io_in_x435_argOut_port_0_valid = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x435_argOut_port_0_valid; // @[MemInterfaceType.scala 317:38:@7001.4]
  assign io_in_x435_argOut_port_0_bits = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x435_argOut_port_0_bits; // @[MemInterfaceType.scala 317:38:@7000.4]
  assign io_in_x420_argOut_port_0_valid = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x420_argOut_port_0_valid; // @[MemInterfaceType.scala 317:38:@7006.4]
  assign io_in_x420_argOut_port_0_bits = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x420_argOut_port_0_bits; // @[MemInterfaceType.scala 317:38:@7005.4]
  assign io_in_x425_argOut_port_0_valid = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x425_argOut_port_0_valid; // @[MemInterfaceType.scala 317:38:@7011.4]
  assign io_in_x425_argOut_port_0_bits = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x425_argOut_port_0_bits; // @[MemInterfaceType.scala 317:38:@7010.4]
  assign io_in_x430_argOut_port_0_valid = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x430_argOut_port_0_valid; // @[MemInterfaceType.scala 317:38:@7016.4]
  assign io_in_x430_argOut_port_0_bits = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x430_argOut_port_0_bits; // @[MemInterfaceType.scala 317:38:@7015.4]
  assign io_in_x444_argOut_port_0_valid = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x444_argOut_port_0_valid; // @[MemInterfaceType.scala 317:38:@7021.4]
  assign io_in_x444_argOut_port_0_bits = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x444_argOut_port_0_bits; // @[MemInterfaceType.scala 317:38:@7020.4]
  assign io_in_x423_argOut_port_0_valid = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x423_argOut_port_0_valid; // @[MemInterfaceType.scala 317:38:@7026.4]
  assign io_in_x423_argOut_port_0_bits = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x423_argOut_port_0_bits; // @[MemInterfaceType.scala 317:38:@7025.4]
  assign io_in_x445_argOut_port_0_valid = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x445_argOut_port_0_valid; // @[MemInterfaceType.scala 317:38:@7031.4]
  assign io_in_x445_argOut_port_0_bits = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x445_argOut_port_0_bits; // @[MemInterfaceType.scala 317:38:@7030.4]
  assign io_in_x451_argOut_port_0_valid = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x451_argOut_port_0_valid; // @[MemInterfaceType.scala 317:38:@7036.4]
  assign io_in_x451_argOut_port_0_bits = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x451_argOut_port_0_bits; // @[MemInterfaceType.scala 317:38:@7035.4]
  assign io_in_x434_argOut_port_0_valid = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x434_argOut_port_0_valid; // @[MemInterfaceType.scala 317:38:@7041.4]
  assign io_in_x434_argOut_port_0_bits = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x434_argOut_port_0_bits; // @[MemInterfaceType.scala 317:38:@7040.4]
  assign io_in_x438_argOut_port_0_valid = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x438_argOut_port_0_valid; // @[MemInterfaceType.scala 317:38:@7046.4]
  assign io_in_x438_argOut_port_0_bits = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x438_argOut_port_0_bits; // @[MemInterfaceType.scala 317:38:@7045.4]
  assign io_in_x431_argOut_port_0_valid = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x431_argOut_port_0_valid; // @[MemInterfaceType.scala 317:38:@7051.4]
  assign io_in_x431_argOut_port_0_bits = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x431_argOut_port_0_bits; // @[MemInterfaceType.scala 317:38:@7050.4]
  assign io_in_x426_argOut_port_0_valid = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x426_argOut_port_0_valid; // @[MemInterfaceType.scala 317:38:@7056.4]
  assign io_in_x426_argOut_port_0_bits = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x426_argOut_port_0_bits; // @[MemInterfaceType.scala 317:38:@7055.4]
  assign io_in_x441_argOut_port_0_valid = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x441_argOut_port_0_valid; // @[MemInterfaceType.scala 317:38:@7061.4]
  assign io_in_x441_argOut_port_0_bits = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x441_argOut_port_0_bits; // @[MemInterfaceType.scala 317:38:@7060.4]
  assign io_in_x446_argOut_port_0_valid = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x446_argOut_port_0_valid; // @[MemInterfaceType.scala 317:38:@7066.4]
  assign io_in_x446_argOut_port_0_bits = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x446_argOut_port_0_bits; // @[MemInterfaceType.scala 317:38:@7065.4]
  assign io_in_x450_argOut_port_0_valid = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x450_argOut_port_0_valid; // @[MemInterfaceType.scala 317:38:@7071.4]
  assign io_in_x450_argOut_port_0_bits = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x450_argOut_port_0_bits; // @[MemInterfaceType.scala 317:38:@7070.4]
  assign io_in_x433_argOut_port_0_valid = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x433_argOut_port_0_valid; // @[MemInterfaceType.scala 317:38:@7076.4]
  assign io_in_x433_argOut_port_0_bits = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x433_argOut_port_0_bits; // @[MemInterfaceType.scala 317:38:@7075.4]
  assign io_in_x447_argOut_port_0_valid = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x447_argOut_port_0_valid; // @[MemInterfaceType.scala 317:38:@7081.4]
  assign io_in_x447_argOut_port_0_bits = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x447_argOut_port_0_bits; // @[MemInterfaceType.scala 317:38:@7080.4]
  assign io_in_x432_argOut_port_0_valid = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x432_argOut_port_0_valid; // @[MemInterfaceType.scala 317:38:@7086.4]
  assign io_in_x432_argOut_port_0_bits = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x432_argOut_port_0_bits; // @[MemInterfaceType.scala 317:38:@7085.4]
  assign io_in_x422_argOut_port_0_valid = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x422_argOut_port_0_valid; // @[MemInterfaceType.scala 317:38:@7091.4]
  assign io_in_x422_argOut_port_0_bits = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x422_argOut_port_0_bits; // @[MemInterfaceType.scala 317:38:@7090.4]
  assign io_in_x437_argOut_port_0_valid = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x437_argOut_port_0_valid; // @[MemInterfaceType.scala 317:38:@7096.4]
  assign io_in_x437_argOut_port_0_bits = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x437_argOut_port_0_bits; // @[MemInterfaceType.scala 317:38:@7095.4]
  assign io_in_x427_argOut_port_0_valid = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x427_argOut_port_0_valid; // @[MemInterfaceType.scala 317:38:@7101.4]
  assign io_in_x427_argOut_port_0_bits = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x427_argOut_port_0_bits; // @[MemInterfaceType.scala 317:38:@7100.4]
  assign io_in_x442_argOut_port_0_valid = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x442_argOut_port_0_valid; // @[MemInterfaceType.scala 317:38:@7106.4]
  assign io_in_x442_argOut_port_0_bits = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x442_argOut_port_0_bits; // @[MemInterfaceType.scala 317:38:@7105.4]
  assign io_sigsOut_smDoneIn_0 = x466_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 127:53:@6439.4]
  assign io_sigsOut_smDoneIn_1 = x555_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 127:53:@6693.4]
  assign x452_a_0_clock = clock; // @[:@6278.4]
  assign x452_a_0_reset = reset; // @[:@6279.4]
  assign x452_a_0_io_rPort_7_en_0 = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x452_a_0_rPort_7_en_0; // @[MemInterfaceType.scala 66:44:@6952.4]
  assign x452_a_0_io_rPort_6_en_0 = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x452_a_0_rPort_6_en_0; // @[MemInterfaceType.scala 66:44:@6982.4]
  assign x452_a_0_io_rPort_5_en_0 = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x452_a_0_rPort_5_en_0; // @[MemInterfaceType.scala 66:44:@6957.4]
  assign x452_a_0_io_rPort_4_en_0 = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x452_a_0_rPort_4_en_0; // @[MemInterfaceType.scala 66:44:@6972.4]
  assign x452_a_0_io_rPort_3_en_0 = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x452_a_0_rPort_3_en_0; // @[MemInterfaceType.scala 66:44:@6947.4]
  assign x452_a_0_io_rPort_2_en_0 = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x452_a_0_rPort_2_en_0; // @[MemInterfaceType.scala 66:44:@6962.4]
  assign x452_a_0_io_rPort_1_en_0 = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x452_a_0_rPort_1_en_0; // @[MemInterfaceType.scala 66:44:@6977.4]
  assign x452_a_0_io_rPort_0_en_0 = x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x452_a_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@6967.4]
  assign x452_a_0_io_wPort_0_banks_0 = x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_in_x452_a_0_wPort_0_banks_0; // @[MemInterfaceType.scala 67:44:@6551.4]
  assign x452_a_0_io_wPort_0_ofs_0 = x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_in_x452_a_0_wPort_0_ofs_0; // @[MemInterfaceType.scala 67:44:@6550.4]
  assign x452_a_0_io_wPort_0_data_0 = x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_in_x452_a_0_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@6549.4]
  assign x452_a_0_io_wPort_0_en_0 = x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_in_x452_a_0_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@6545.4]
  assign x466_outr_UnitPipe_sm_clock = clock; // @[:@6365.4]
  assign x466_outr_UnitPipe_sm_reset = reset; // @[:@6366.4]
  assign x466_outr_UnitPipe_sm_io_enable = _T_843 & _T_852; // @[SpatialBlocks.scala 112:18:@6436.4]
  assign x466_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 114:21:@6438.4]
  assign x466_outr_UnitPipe_sm_io_doneIn_0 = x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 102:67:@6408.4]
  assign x466_outr_UnitPipe_sm_io_ctrCopyDone_0 = x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 132:80:@6450.4]
  assign RetimeWrapper_clock = clock; // @[:@6417.4]
  assign RetimeWrapper_reset = reset; // @[:@6418.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@6420.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@6419.4]
  assign RetimeWrapper_1_clock = clock; // @[:@6425.4]
  assign RetimeWrapper_1_reset = reset; // @[:@6426.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@6428.4]
  assign RetimeWrapper_1_io_in = x466_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@6427.4]
  assign x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_clock = clock; // @[:@6452.4]
  assign x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_reset = reset; // @[:@6453.4]
  assign x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_in_x416_TVALID = io_in_x416_TVALID; // @[sm_x466_outr_UnitPipe.scala 49:23:@6544.4]
  assign x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_in_x416_TDATA = io_in_x416_TDATA; // @[sm_x466_outr_UnitPipe.scala 49:23:@6542.4]
  assign x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x466_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x466_outr_UnitPipe.scala 79:22:@6560.4]
  assign x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x466_outr_UnitPipe_sm_io_childAck_0; // @[sm_x466_outr_UnitPipe.scala 79:22:@6558.4]
  assign x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x466_outr_UnitPipe.scala 78:18:@6552.4]
  assign x555_inr_UnitPipe_sm_clock = clock; // @[:@6614.4]
  assign x555_inr_UnitPipe_sm_reset = reset; // @[:@6615.4]
  assign x555_inr_UnitPipe_sm_io_enable = _T_935 & _T_944; // @[SpatialBlocks.scala 112:18:@6690.4]
  assign x555_inr_UnitPipe_sm_io_ctrDone = x555_inr_UnitPipe_sm_io_ctrInc & _T_921; // @[sm_RootController.scala 227:39:@6645.4]
  assign x555_inr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 114:21:@6692.4]
  assign x555_inr_UnitPipe_sm_io_break = 1'h0; // @[sm_RootController.scala 231:37:@6651.4]
  assign RetimeWrapper_2_clock = clock; // @[:@6671.4]
  assign RetimeWrapper_2_reset = reset; // @[:@6672.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@6674.4]
  assign RetimeWrapper_2_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@6673.4]
  assign RetimeWrapper_3_clock = clock; // @[:@6679.4]
  assign RetimeWrapper_3_reset = reset; // @[:@6680.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@6682.4]
  assign RetimeWrapper_3_io_in = x555_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@6681.4]
  assign x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_clock = clock; // @[:@6705.4]
  assign x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_reset = reset; // @[:@6706.4]
  assign x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x452_a_0_rPort_7_output_0 = x452_a_0_io_rPort_7_output_0; // @[MemInterfaceType.scala 66:44:@6950.4]
  assign x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x452_a_0_rPort_6_output_0 = x452_a_0_io_rPort_6_output_0; // @[MemInterfaceType.scala 66:44:@6980.4]
  assign x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x452_a_0_rPort_5_output_0 = x452_a_0_io_rPort_5_output_0; // @[MemInterfaceType.scala 66:44:@6955.4]
  assign x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x452_a_0_rPort_4_output_0 = x452_a_0_io_rPort_4_output_0; // @[MemInterfaceType.scala 66:44:@6970.4]
  assign x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x452_a_0_rPort_3_output_0 = x452_a_0_io_rPort_3_output_0; // @[MemInterfaceType.scala 66:44:@6945.4]
  assign x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x452_a_0_rPort_2_output_0 = x452_a_0_io_rPort_2_output_0; // @[MemInterfaceType.scala 66:44:@6960.4]
  assign x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x452_a_0_rPort_1_output_0 = x452_a_0_io_rPort_1_output_0; // @[MemInterfaceType.scala 66:44:@6975.4]
  assign x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_in_x452_a_0_rPort_0_output_0 = x452_a_0_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@6965.4]
  assign x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_sigsIn_datapathEn = x555_inr_UnitPipe_sm_io_datapathEn; // @[sm_x555_inr_UnitPipe.scala 402:22:@7122.4]
  assign x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_sigsIn_break = x555_inr_UnitPipe_sm_io_break; // @[sm_x555_inr_UnitPipe.scala 402:22:@7120.4]
  assign x555_inr_UnitPipe_kernelx555_inr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x555_inr_UnitPipe.scala 401:18:@7110.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_921 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_921 <= 1'h0;
    end else begin
      _T_921 <= _T_918;
    end
  end
endmodule
module AccelUnit( // @[:@7137.2]
  input          clock, // @[:@7138.4]
  input          reset, // @[:@7139.4]
  input          io_enable, // @[:@7140.4]
  output         io_done, // @[:@7140.4]
  input          io_reset, // @[:@7140.4]
  input          io_memStreams_loads_0_cmd_ready, // @[:@7140.4]
  output         io_memStreams_loads_0_cmd_valid, // @[:@7140.4]
  output [63:0]  io_memStreams_loads_0_cmd_bits_addr, // @[:@7140.4]
  output [31:0]  io_memStreams_loads_0_cmd_bits_size, // @[:@7140.4]
  output         io_memStreams_loads_0_data_ready, // @[:@7140.4]
  input          io_memStreams_loads_0_data_valid, // @[:@7140.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_0, // @[:@7140.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_1, // @[:@7140.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_2, // @[:@7140.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_3, // @[:@7140.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_4, // @[:@7140.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_5, // @[:@7140.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_6, // @[:@7140.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_7, // @[:@7140.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_8, // @[:@7140.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_9, // @[:@7140.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_10, // @[:@7140.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_11, // @[:@7140.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_12, // @[:@7140.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_13, // @[:@7140.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_14, // @[:@7140.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_15, // @[:@7140.4]
  input          io_memStreams_stores_0_cmd_ready, // @[:@7140.4]
  output         io_memStreams_stores_0_cmd_valid, // @[:@7140.4]
  output [63:0]  io_memStreams_stores_0_cmd_bits_addr, // @[:@7140.4]
  output [31:0]  io_memStreams_stores_0_cmd_bits_size, // @[:@7140.4]
  input          io_memStreams_stores_0_data_ready, // @[:@7140.4]
  output         io_memStreams_stores_0_data_valid, // @[:@7140.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_0, // @[:@7140.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_1, // @[:@7140.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_2, // @[:@7140.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_3, // @[:@7140.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_4, // @[:@7140.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_5, // @[:@7140.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_6, // @[:@7140.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_7, // @[:@7140.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_8, // @[:@7140.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_9, // @[:@7140.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_10, // @[:@7140.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_11, // @[:@7140.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_12, // @[:@7140.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_13, // @[:@7140.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_14, // @[:@7140.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_15, // @[:@7140.4]
  output [15:0]  io_memStreams_stores_0_data_bits_wstrb, // @[:@7140.4]
  output         io_memStreams_stores_0_wresp_ready, // @[:@7140.4]
  input          io_memStreams_stores_0_wresp_valid, // @[:@7140.4]
  input          io_memStreams_stores_0_wresp_bits, // @[:@7140.4]
  input          io_memStreams_gathers_0_cmd_ready, // @[:@7140.4]
  output         io_memStreams_gathers_0_cmd_valid, // @[:@7140.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_0, // @[:@7140.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_1, // @[:@7140.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_2, // @[:@7140.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_3, // @[:@7140.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_4, // @[:@7140.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_5, // @[:@7140.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_6, // @[:@7140.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_7, // @[:@7140.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_8, // @[:@7140.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_9, // @[:@7140.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_10, // @[:@7140.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_11, // @[:@7140.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_12, // @[:@7140.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_13, // @[:@7140.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_14, // @[:@7140.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_15, // @[:@7140.4]
  output         io_memStreams_gathers_0_data_ready, // @[:@7140.4]
  input          io_memStreams_gathers_0_data_valid, // @[:@7140.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_0, // @[:@7140.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_1, // @[:@7140.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_2, // @[:@7140.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_3, // @[:@7140.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_4, // @[:@7140.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_5, // @[:@7140.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_6, // @[:@7140.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_7, // @[:@7140.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_8, // @[:@7140.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_9, // @[:@7140.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_10, // @[:@7140.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_11, // @[:@7140.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_12, // @[:@7140.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_13, // @[:@7140.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_14, // @[:@7140.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_15, // @[:@7140.4]
  input          io_memStreams_scatters_0_cmd_ready, // @[:@7140.4]
  output         io_memStreams_scatters_0_cmd_valid, // @[:@7140.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_0, // @[:@7140.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_1, // @[:@7140.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_2, // @[:@7140.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_3, // @[:@7140.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_4, // @[:@7140.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_5, // @[:@7140.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_6, // @[:@7140.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_7, // @[:@7140.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_8, // @[:@7140.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_9, // @[:@7140.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_10, // @[:@7140.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_11, // @[:@7140.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_12, // @[:@7140.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_13, // @[:@7140.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_14, // @[:@7140.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_15, // @[:@7140.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_0, // @[:@7140.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_1, // @[:@7140.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_2, // @[:@7140.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_3, // @[:@7140.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_4, // @[:@7140.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_5, // @[:@7140.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_6, // @[:@7140.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_7, // @[:@7140.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_8, // @[:@7140.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_9, // @[:@7140.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_10, // @[:@7140.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_11, // @[:@7140.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_12, // @[:@7140.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_13, // @[:@7140.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_14, // @[:@7140.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_15, // @[:@7140.4]
  output         io_memStreams_scatters_0_wresp_ready, // @[:@7140.4]
  input          io_memStreams_scatters_0_wresp_valid, // @[:@7140.4]
  input          io_memStreams_scatters_0_wresp_bits, // @[:@7140.4]
  input          io_axiStreamsIn_0_TVALID, // @[:@7140.4]
  output         io_axiStreamsIn_0_TREADY, // @[:@7140.4]
  input  [255:0] io_axiStreamsIn_0_TDATA, // @[:@7140.4]
  input  [31:0]  io_axiStreamsIn_0_TSTRB, // @[:@7140.4]
  input  [31:0]  io_axiStreamsIn_0_TKEEP, // @[:@7140.4]
  input          io_axiStreamsIn_0_TLAST, // @[:@7140.4]
  input  [7:0]   io_axiStreamsIn_0_TID, // @[:@7140.4]
  input  [7:0]   io_axiStreamsIn_0_TDEST, // @[:@7140.4]
  output         io_axiStreamsOut_0_TVALID, // @[:@7140.4]
  input          io_axiStreamsOut_0_TREADY, // @[:@7140.4]
  output [255:0] io_axiStreamsOut_0_TDATA, // @[:@7140.4]
  output [31:0]  io_axiStreamsOut_0_TSTRB, // @[:@7140.4]
  output [31:0]  io_axiStreamsOut_0_TKEEP, // @[:@7140.4]
  output         io_axiStreamsOut_0_TLAST, // @[:@7140.4]
  output [7:0]   io_axiStreamsOut_0_TID, // @[:@7140.4]
  output [7:0]   io_axiStreamsOut_0_TDEST, // @[:@7140.4]
  output         io_heap_0_req_valid, // @[:@7140.4]
  output         io_heap_0_req_bits_allocDealloc, // @[:@7140.4]
  output [63:0]  io_heap_0_req_bits_sizeAddr, // @[:@7140.4]
  input          io_heap_0_resp_valid, // @[:@7140.4]
  input          io_heap_0_resp_bits_allocDealloc, // @[:@7140.4]
  input  [63:0]  io_heap_0_resp_bits_sizeAddr, // @[:@7140.4]
  input  [63:0]  io_argIns_0, // @[:@7140.4]
  input          io_argOuts_0_port_ready, // @[:@7140.4]
  output         io_argOuts_0_port_valid, // @[:@7140.4]
  output [63:0]  io_argOuts_0_port_bits, // @[:@7140.4]
  input  [63:0]  io_argOuts_0_echo, // @[:@7140.4]
  input          io_argOuts_1_port_ready, // @[:@7140.4]
  output         io_argOuts_1_port_valid, // @[:@7140.4]
  output [63:0]  io_argOuts_1_port_bits, // @[:@7140.4]
  input  [63:0]  io_argOuts_1_echo, // @[:@7140.4]
  input          io_argOuts_2_port_ready, // @[:@7140.4]
  output         io_argOuts_2_port_valid, // @[:@7140.4]
  output [63:0]  io_argOuts_2_port_bits, // @[:@7140.4]
  input  [63:0]  io_argOuts_2_echo, // @[:@7140.4]
  input          io_argOuts_3_port_ready, // @[:@7140.4]
  output         io_argOuts_3_port_valid, // @[:@7140.4]
  output [63:0]  io_argOuts_3_port_bits, // @[:@7140.4]
  input  [63:0]  io_argOuts_3_echo, // @[:@7140.4]
  input          io_argOuts_4_port_ready, // @[:@7140.4]
  output         io_argOuts_4_port_valid, // @[:@7140.4]
  output [63:0]  io_argOuts_4_port_bits, // @[:@7140.4]
  input  [63:0]  io_argOuts_4_echo, // @[:@7140.4]
  input          io_argOuts_5_port_ready, // @[:@7140.4]
  output         io_argOuts_5_port_valid, // @[:@7140.4]
  output [63:0]  io_argOuts_5_port_bits, // @[:@7140.4]
  input  [63:0]  io_argOuts_5_echo, // @[:@7140.4]
  input          io_argOuts_6_port_ready, // @[:@7140.4]
  output         io_argOuts_6_port_valid, // @[:@7140.4]
  output [63:0]  io_argOuts_6_port_bits, // @[:@7140.4]
  input  [63:0]  io_argOuts_6_echo, // @[:@7140.4]
  input          io_argOuts_7_port_ready, // @[:@7140.4]
  output         io_argOuts_7_port_valid, // @[:@7140.4]
  output [63:0]  io_argOuts_7_port_bits, // @[:@7140.4]
  input  [63:0]  io_argOuts_7_echo, // @[:@7140.4]
  input          io_argOuts_8_port_ready, // @[:@7140.4]
  output         io_argOuts_8_port_valid, // @[:@7140.4]
  output [63:0]  io_argOuts_8_port_bits, // @[:@7140.4]
  input  [63:0]  io_argOuts_8_echo, // @[:@7140.4]
  input          io_argOuts_9_port_ready, // @[:@7140.4]
  output         io_argOuts_9_port_valid, // @[:@7140.4]
  output [63:0]  io_argOuts_9_port_bits, // @[:@7140.4]
  input  [63:0]  io_argOuts_9_echo, // @[:@7140.4]
  input          io_argOuts_10_port_ready, // @[:@7140.4]
  output         io_argOuts_10_port_valid, // @[:@7140.4]
  output [63:0]  io_argOuts_10_port_bits, // @[:@7140.4]
  input  [63:0]  io_argOuts_10_echo, // @[:@7140.4]
  input          io_argOuts_11_port_ready, // @[:@7140.4]
  output         io_argOuts_11_port_valid, // @[:@7140.4]
  output [63:0]  io_argOuts_11_port_bits, // @[:@7140.4]
  input  [63:0]  io_argOuts_11_echo, // @[:@7140.4]
  input          io_argOuts_12_port_ready, // @[:@7140.4]
  output         io_argOuts_12_port_valid, // @[:@7140.4]
  output [63:0]  io_argOuts_12_port_bits, // @[:@7140.4]
  input  [63:0]  io_argOuts_12_echo, // @[:@7140.4]
  input          io_argOuts_13_port_ready, // @[:@7140.4]
  output         io_argOuts_13_port_valid, // @[:@7140.4]
  output [63:0]  io_argOuts_13_port_bits, // @[:@7140.4]
  input  [63:0]  io_argOuts_13_echo, // @[:@7140.4]
  input          io_argOuts_14_port_ready, // @[:@7140.4]
  output         io_argOuts_14_port_valid, // @[:@7140.4]
  output [63:0]  io_argOuts_14_port_bits, // @[:@7140.4]
  input  [63:0]  io_argOuts_14_echo, // @[:@7140.4]
  input          io_argOuts_15_port_ready, // @[:@7140.4]
  output         io_argOuts_15_port_valid, // @[:@7140.4]
  output [63:0]  io_argOuts_15_port_bits, // @[:@7140.4]
  input  [63:0]  io_argOuts_15_echo, // @[:@7140.4]
  input          io_argOuts_16_port_ready, // @[:@7140.4]
  output         io_argOuts_16_port_valid, // @[:@7140.4]
  output [63:0]  io_argOuts_16_port_bits, // @[:@7140.4]
  input  [63:0]  io_argOuts_16_echo, // @[:@7140.4]
  input          io_argOuts_17_port_ready, // @[:@7140.4]
  output         io_argOuts_17_port_valid, // @[:@7140.4]
  output [63:0]  io_argOuts_17_port_bits, // @[:@7140.4]
  input  [63:0]  io_argOuts_17_echo, // @[:@7140.4]
  input          io_argOuts_18_port_ready, // @[:@7140.4]
  output         io_argOuts_18_port_valid, // @[:@7140.4]
  output [63:0]  io_argOuts_18_port_bits, // @[:@7140.4]
  input  [63:0]  io_argOuts_18_echo, // @[:@7140.4]
  input          io_argOuts_19_port_ready, // @[:@7140.4]
  output         io_argOuts_19_port_valid, // @[:@7140.4]
  output [63:0]  io_argOuts_19_port_bits, // @[:@7140.4]
  input  [63:0]  io_argOuts_19_echo, // @[:@7140.4]
  input          io_argOuts_20_port_ready, // @[:@7140.4]
  output         io_argOuts_20_port_valid, // @[:@7140.4]
  output [63:0]  io_argOuts_20_port_bits, // @[:@7140.4]
  input  [63:0]  io_argOuts_20_echo, // @[:@7140.4]
  input          io_argOuts_21_port_ready, // @[:@7140.4]
  output         io_argOuts_21_port_valid, // @[:@7140.4]
  output [63:0]  io_argOuts_21_port_bits, // @[:@7140.4]
  input  [63:0]  io_argOuts_21_echo, // @[:@7140.4]
  input          io_argOuts_22_port_ready, // @[:@7140.4]
  output         io_argOuts_22_port_valid, // @[:@7140.4]
  output [63:0]  io_argOuts_22_port_bits, // @[:@7140.4]
  input  [63:0]  io_argOuts_22_echo, // @[:@7140.4]
  input          io_argOuts_23_port_ready, // @[:@7140.4]
  output         io_argOuts_23_port_valid, // @[:@7140.4]
  output [63:0]  io_argOuts_23_port_bits, // @[:@7140.4]
  input  [63:0]  io_argOuts_23_echo, // @[:@7140.4]
  input          io_argOuts_24_port_ready, // @[:@7140.4]
  output         io_argOuts_24_port_valid, // @[:@7140.4]
  output [63:0]  io_argOuts_24_port_bits, // @[:@7140.4]
  input  [63:0]  io_argOuts_24_echo, // @[:@7140.4]
  input          io_argOuts_25_port_ready, // @[:@7140.4]
  output         io_argOuts_25_port_valid, // @[:@7140.4]
  output [63:0]  io_argOuts_25_port_bits, // @[:@7140.4]
  input  [63:0]  io_argOuts_25_echo, // @[:@7140.4]
  input          io_argOuts_26_port_ready, // @[:@7140.4]
  output         io_argOuts_26_port_valid, // @[:@7140.4]
  output [63:0]  io_argOuts_26_port_bits, // @[:@7140.4]
  input  [63:0]  io_argOuts_26_echo, // @[:@7140.4]
  input          io_argOuts_27_port_ready, // @[:@7140.4]
  output         io_argOuts_27_port_valid, // @[:@7140.4]
  output [63:0]  io_argOuts_27_port_bits, // @[:@7140.4]
  input  [63:0]  io_argOuts_27_echo, // @[:@7140.4]
  input          io_argOuts_28_port_ready, // @[:@7140.4]
  output         io_argOuts_28_port_valid, // @[:@7140.4]
  output [63:0]  io_argOuts_28_port_bits, // @[:@7140.4]
  input  [63:0]  io_argOuts_28_echo, // @[:@7140.4]
  input          io_argOuts_29_port_ready, // @[:@7140.4]
  output         io_argOuts_29_port_valid, // @[:@7140.4]
  output [63:0]  io_argOuts_29_port_bits, // @[:@7140.4]
  input  [63:0]  io_argOuts_29_echo, // @[:@7140.4]
  input          io_argOuts_30_port_ready, // @[:@7140.4]
  output         io_argOuts_30_port_valid, // @[:@7140.4]
  output [63:0]  io_argOuts_30_port_bits, // @[:@7140.4]
  input  [63:0]  io_argOuts_30_echo, // @[:@7140.4]
  input          io_argOuts_31_port_ready, // @[:@7140.4]
  output         io_argOuts_31_port_valid, // @[:@7140.4]
  output [63:0]  io_argOuts_31_port_bits, // @[:@7140.4]
  input  [63:0]  io_argOuts_31_echo // @[:@7140.4]
);
  wire  SingleCounter_clock; // @[Main.scala 188:32:@7676.4]
  wire  SingleCounter_reset; // @[Main.scala 188:32:@7676.4]
  wire  SingleCounter_io_input_reset; // @[Main.scala 188:32:@7676.4]
  wire  SingleCounter_io_output_done; // @[Main.scala 188:32:@7676.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@7694.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@7694.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@7694.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@7694.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@7694.4]
  wire  SRFF_clock; // @[Main.scala 192:28:@7703.4]
  wire  SRFF_reset; // @[Main.scala 192:28:@7703.4]
  wire  SRFF_io_input_set; // @[Main.scala 192:28:@7703.4]
  wire  SRFF_io_input_reset; // @[Main.scala 192:28:@7703.4]
  wire  SRFF_io_input_asyn_reset; // @[Main.scala 192:28:@7703.4]
  wire  SRFF_io_output; // @[Main.scala 192:28:@7703.4]
  wire  RootController_sm_clock; // @[sm_RootController.scala 33:18:@7746.4]
  wire  RootController_sm_reset; // @[sm_RootController.scala 33:18:@7746.4]
  wire  RootController_sm_io_enable; // @[sm_RootController.scala 33:18:@7746.4]
  wire  RootController_sm_io_done; // @[sm_RootController.scala 33:18:@7746.4]
  wire  RootController_sm_io_rst; // @[sm_RootController.scala 33:18:@7746.4]
  wire  RootController_sm_io_ctrDone; // @[sm_RootController.scala 33:18:@7746.4]
  wire  RootController_sm_io_ctrInc; // @[sm_RootController.scala 33:18:@7746.4]
  wire  RootController_sm_io_doneIn_0; // @[sm_RootController.scala 33:18:@7746.4]
  wire  RootController_sm_io_doneIn_1; // @[sm_RootController.scala 33:18:@7746.4]
  wire  RootController_sm_io_enableOut_0; // @[sm_RootController.scala 33:18:@7746.4]
  wire  RootController_sm_io_enableOut_1; // @[sm_RootController.scala 33:18:@7746.4]
  wire  RootController_sm_io_childAck_0; // @[sm_RootController.scala 33:18:@7746.4]
  wire  RootController_sm_io_childAck_1; // @[sm_RootController.scala 33:18:@7746.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@7783.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@7783.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@7783.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@7783.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@7783.4]
  wire  RootController_kernelRootController_concrete1_clock; // @[sm_RootController.scala 236:24:@7847.4]
  wire  RootController_kernelRootController_concrete1_reset; // @[sm_RootController.scala 236:24:@7847.4]
  wire  RootController_kernelRootController_concrete1_io_in_x449_argOut_port_0_valid; // @[sm_RootController.scala 236:24:@7847.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x449_argOut_port_0_bits; // @[sm_RootController.scala 236:24:@7847.4]
  wire  RootController_kernelRootController_concrete1_io_in_x440_argOut_port_0_valid; // @[sm_RootController.scala 236:24:@7847.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x440_argOut_port_0_bits; // @[sm_RootController.scala 236:24:@7847.4]
  wire  RootController_kernelRootController_concrete1_io_in_x436_argOut_port_0_valid; // @[sm_RootController.scala 236:24:@7847.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x436_argOut_port_0_bits; // @[sm_RootController.scala 236:24:@7847.4]
  wire  RootController_kernelRootController_concrete1_io_in_x421_argOut_port_0_valid; // @[sm_RootController.scala 236:24:@7847.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x421_argOut_port_0_bits; // @[sm_RootController.scala 236:24:@7847.4]
  wire  RootController_kernelRootController_concrete1_io_in_x416_TVALID; // @[sm_RootController.scala 236:24:@7847.4]
  wire  RootController_kernelRootController_concrete1_io_in_x416_TREADY; // @[sm_RootController.scala 236:24:@7847.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x416_TDATA; // @[sm_RootController.scala 236:24:@7847.4]
  wire  RootController_kernelRootController_concrete1_io_in_x448_argOut_port_0_valid; // @[sm_RootController.scala 236:24:@7847.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x448_argOut_port_0_bits; // @[sm_RootController.scala 236:24:@7847.4]
  wire  RootController_kernelRootController_concrete1_io_in_x443_argOut_port_0_valid; // @[sm_RootController.scala 236:24:@7847.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x443_argOut_port_0_bits; // @[sm_RootController.scala 236:24:@7847.4]
  wire  RootController_kernelRootController_concrete1_io_in_x428_argOut_port_0_valid; // @[sm_RootController.scala 236:24:@7847.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x428_argOut_port_0_bits; // @[sm_RootController.scala 236:24:@7847.4]
  wire  RootController_kernelRootController_concrete1_io_in_x439_argOut_port_0_valid; // @[sm_RootController.scala 236:24:@7847.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x439_argOut_port_0_bits; // @[sm_RootController.scala 236:24:@7847.4]
  wire  RootController_kernelRootController_concrete1_io_in_x424_argOut_port_0_valid; // @[sm_RootController.scala 236:24:@7847.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x424_argOut_port_0_bits; // @[sm_RootController.scala 236:24:@7847.4]
  wire  RootController_kernelRootController_concrete1_io_in_x429_argOut_port_0_valid; // @[sm_RootController.scala 236:24:@7847.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x429_argOut_port_0_bits; // @[sm_RootController.scala 236:24:@7847.4]
  wire  RootController_kernelRootController_concrete1_io_in_x435_argOut_port_0_valid; // @[sm_RootController.scala 236:24:@7847.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x435_argOut_port_0_bits; // @[sm_RootController.scala 236:24:@7847.4]
  wire  RootController_kernelRootController_concrete1_io_in_x420_argOut_port_0_valid; // @[sm_RootController.scala 236:24:@7847.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x420_argOut_port_0_bits; // @[sm_RootController.scala 236:24:@7847.4]
  wire  RootController_kernelRootController_concrete1_io_in_x425_argOut_port_0_valid; // @[sm_RootController.scala 236:24:@7847.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x425_argOut_port_0_bits; // @[sm_RootController.scala 236:24:@7847.4]
  wire  RootController_kernelRootController_concrete1_io_in_x430_argOut_port_0_valid; // @[sm_RootController.scala 236:24:@7847.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x430_argOut_port_0_bits; // @[sm_RootController.scala 236:24:@7847.4]
  wire  RootController_kernelRootController_concrete1_io_in_x444_argOut_port_0_valid; // @[sm_RootController.scala 236:24:@7847.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x444_argOut_port_0_bits; // @[sm_RootController.scala 236:24:@7847.4]
  wire  RootController_kernelRootController_concrete1_io_in_x423_argOut_port_0_valid; // @[sm_RootController.scala 236:24:@7847.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x423_argOut_port_0_bits; // @[sm_RootController.scala 236:24:@7847.4]
  wire  RootController_kernelRootController_concrete1_io_in_x445_argOut_port_0_valid; // @[sm_RootController.scala 236:24:@7847.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x445_argOut_port_0_bits; // @[sm_RootController.scala 236:24:@7847.4]
  wire  RootController_kernelRootController_concrete1_io_in_x451_argOut_port_0_valid; // @[sm_RootController.scala 236:24:@7847.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x451_argOut_port_0_bits; // @[sm_RootController.scala 236:24:@7847.4]
  wire  RootController_kernelRootController_concrete1_io_in_x434_argOut_port_0_valid; // @[sm_RootController.scala 236:24:@7847.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x434_argOut_port_0_bits; // @[sm_RootController.scala 236:24:@7847.4]
  wire  RootController_kernelRootController_concrete1_io_in_x438_argOut_port_0_valid; // @[sm_RootController.scala 236:24:@7847.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x438_argOut_port_0_bits; // @[sm_RootController.scala 236:24:@7847.4]
  wire  RootController_kernelRootController_concrete1_io_in_x431_argOut_port_0_valid; // @[sm_RootController.scala 236:24:@7847.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x431_argOut_port_0_bits; // @[sm_RootController.scala 236:24:@7847.4]
  wire  RootController_kernelRootController_concrete1_io_in_x426_argOut_port_0_valid; // @[sm_RootController.scala 236:24:@7847.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x426_argOut_port_0_bits; // @[sm_RootController.scala 236:24:@7847.4]
  wire  RootController_kernelRootController_concrete1_io_in_x441_argOut_port_0_valid; // @[sm_RootController.scala 236:24:@7847.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x441_argOut_port_0_bits; // @[sm_RootController.scala 236:24:@7847.4]
  wire  RootController_kernelRootController_concrete1_io_in_x446_argOut_port_0_valid; // @[sm_RootController.scala 236:24:@7847.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x446_argOut_port_0_bits; // @[sm_RootController.scala 236:24:@7847.4]
  wire  RootController_kernelRootController_concrete1_io_in_x450_argOut_port_0_valid; // @[sm_RootController.scala 236:24:@7847.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x450_argOut_port_0_bits; // @[sm_RootController.scala 236:24:@7847.4]
  wire  RootController_kernelRootController_concrete1_io_in_x433_argOut_port_0_valid; // @[sm_RootController.scala 236:24:@7847.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x433_argOut_port_0_bits; // @[sm_RootController.scala 236:24:@7847.4]
  wire  RootController_kernelRootController_concrete1_io_in_x447_argOut_port_0_valid; // @[sm_RootController.scala 236:24:@7847.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x447_argOut_port_0_bits; // @[sm_RootController.scala 236:24:@7847.4]
  wire  RootController_kernelRootController_concrete1_io_in_x432_argOut_port_0_valid; // @[sm_RootController.scala 236:24:@7847.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x432_argOut_port_0_bits; // @[sm_RootController.scala 236:24:@7847.4]
  wire  RootController_kernelRootController_concrete1_io_in_x422_argOut_port_0_valid; // @[sm_RootController.scala 236:24:@7847.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x422_argOut_port_0_bits; // @[sm_RootController.scala 236:24:@7847.4]
  wire  RootController_kernelRootController_concrete1_io_in_x437_argOut_port_0_valid; // @[sm_RootController.scala 236:24:@7847.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x437_argOut_port_0_bits; // @[sm_RootController.scala 236:24:@7847.4]
  wire  RootController_kernelRootController_concrete1_io_in_x427_argOut_port_0_valid; // @[sm_RootController.scala 236:24:@7847.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x427_argOut_port_0_bits; // @[sm_RootController.scala 236:24:@7847.4]
  wire  RootController_kernelRootController_concrete1_io_in_x442_argOut_port_0_valid; // @[sm_RootController.scala 236:24:@7847.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x442_argOut_port_0_bits; // @[sm_RootController.scala 236:24:@7847.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_RootController.scala 236:24:@7847.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_RootController.scala 236:24:@7847.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0; // @[sm_RootController.scala 236:24:@7847.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_1; // @[sm_RootController.scala 236:24:@7847.4]
  wire  RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[sm_RootController.scala 236:24:@7847.4]
  wire  RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_1; // @[sm_RootController.scala 236:24:@7847.4]
  wire  RootController_kernelRootController_concrete1_io_rr; // @[sm_RootController.scala 236:24:@7847.4]
  wire  _T_1539; // @[package.scala 96:25:@7699.4 package.scala 96:25:@7700.4]
  wire  _T_1604; // @[Main.scala 194:50:@7779.4]
  wire  _T_1605; // @[Main.scala 194:59:@7780.4]
  wire  _T_1617; // @[package.scala 100:49:@7800.4]
  reg  _T_1620; // @[package.scala 48:56:@7801.4]
  reg [31:0] _RAND_0;
  SingleCounter SingleCounter ( // @[Main.scala 188:32:@7676.4]
    .clock(SingleCounter_clock),
    .reset(SingleCounter_reset),
    .io_input_reset(SingleCounter_io_input_reset),
    .io_output_done(SingleCounter_io_output_done)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@7694.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  SRFF SRFF ( // @[Main.scala 192:28:@7703.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  RootController_sm RootController_sm ( // @[sm_RootController.scala 33:18:@7746.4]
    .clock(RootController_sm_clock),
    .reset(RootController_sm_reset),
    .io_enable(RootController_sm_io_enable),
    .io_done(RootController_sm_io_done),
    .io_rst(RootController_sm_io_rst),
    .io_ctrDone(RootController_sm_io_ctrDone),
    .io_ctrInc(RootController_sm_io_ctrInc),
    .io_doneIn_0(RootController_sm_io_doneIn_0),
    .io_doneIn_1(RootController_sm_io_doneIn_1),
    .io_enableOut_0(RootController_sm_io_enableOut_0),
    .io_enableOut_1(RootController_sm_io_enableOut_1),
    .io_childAck_0(RootController_sm_io_childAck_0),
    .io_childAck_1(RootController_sm_io_childAck_1)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@7783.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RootController_kernelRootController_concrete1 RootController_kernelRootController_concrete1 ( // @[sm_RootController.scala 236:24:@7847.4]
    .clock(RootController_kernelRootController_concrete1_clock),
    .reset(RootController_kernelRootController_concrete1_reset),
    .io_in_x449_argOut_port_0_valid(RootController_kernelRootController_concrete1_io_in_x449_argOut_port_0_valid),
    .io_in_x449_argOut_port_0_bits(RootController_kernelRootController_concrete1_io_in_x449_argOut_port_0_bits),
    .io_in_x440_argOut_port_0_valid(RootController_kernelRootController_concrete1_io_in_x440_argOut_port_0_valid),
    .io_in_x440_argOut_port_0_bits(RootController_kernelRootController_concrete1_io_in_x440_argOut_port_0_bits),
    .io_in_x436_argOut_port_0_valid(RootController_kernelRootController_concrete1_io_in_x436_argOut_port_0_valid),
    .io_in_x436_argOut_port_0_bits(RootController_kernelRootController_concrete1_io_in_x436_argOut_port_0_bits),
    .io_in_x421_argOut_port_0_valid(RootController_kernelRootController_concrete1_io_in_x421_argOut_port_0_valid),
    .io_in_x421_argOut_port_0_bits(RootController_kernelRootController_concrete1_io_in_x421_argOut_port_0_bits),
    .io_in_x416_TVALID(RootController_kernelRootController_concrete1_io_in_x416_TVALID),
    .io_in_x416_TREADY(RootController_kernelRootController_concrete1_io_in_x416_TREADY),
    .io_in_x416_TDATA(RootController_kernelRootController_concrete1_io_in_x416_TDATA),
    .io_in_x448_argOut_port_0_valid(RootController_kernelRootController_concrete1_io_in_x448_argOut_port_0_valid),
    .io_in_x448_argOut_port_0_bits(RootController_kernelRootController_concrete1_io_in_x448_argOut_port_0_bits),
    .io_in_x443_argOut_port_0_valid(RootController_kernelRootController_concrete1_io_in_x443_argOut_port_0_valid),
    .io_in_x443_argOut_port_0_bits(RootController_kernelRootController_concrete1_io_in_x443_argOut_port_0_bits),
    .io_in_x428_argOut_port_0_valid(RootController_kernelRootController_concrete1_io_in_x428_argOut_port_0_valid),
    .io_in_x428_argOut_port_0_bits(RootController_kernelRootController_concrete1_io_in_x428_argOut_port_0_bits),
    .io_in_x439_argOut_port_0_valid(RootController_kernelRootController_concrete1_io_in_x439_argOut_port_0_valid),
    .io_in_x439_argOut_port_0_bits(RootController_kernelRootController_concrete1_io_in_x439_argOut_port_0_bits),
    .io_in_x424_argOut_port_0_valid(RootController_kernelRootController_concrete1_io_in_x424_argOut_port_0_valid),
    .io_in_x424_argOut_port_0_bits(RootController_kernelRootController_concrete1_io_in_x424_argOut_port_0_bits),
    .io_in_x429_argOut_port_0_valid(RootController_kernelRootController_concrete1_io_in_x429_argOut_port_0_valid),
    .io_in_x429_argOut_port_0_bits(RootController_kernelRootController_concrete1_io_in_x429_argOut_port_0_bits),
    .io_in_x435_argOut_port_0_valid(RootController_kernelRootController_concrete1_io_in_x435_argOut_port_0_valid),
    .io_in_x435_argOut_port_0_bits(RootController_kernelRootController_concrete1_io_in_x435_argOut_port_0_bits),
    .io_in_x420_argOut_port_0_valid(RootController_kernelRootController_concrete1_io_in_x420_argOut_port_0_valid),
    .io_in_x420_argOut_port_0_bits(RootController_kernelRootController_concrete1_io_in_x420_argOut_port_0_bits),
    .io_in_x425_argOut_port_0_valid(RootController_kernelRootController_concrete1_io_in_x425_argOut_port_0_valid),
    .io_in_x425_argOut_port_0_bits(RootController_kernelRootController_concrete1_io_in_x425_argOut_port_0_bits),
    .io_in_x430_argOut_port_0_valid(RootController_kernelRootController_concrete1_io_in_x430_argOut_port_0_valid),
    .io_in_x430_argOut_port_0_bits(RootController_kernelRootController_concrete1_io_in_x430_argOut_port_0_bits),
    .io_in_x444_argOut_port_0_valid(RootController_kernelRootController_concrete1_io_in_x444_argOut_port_0_valid),
    .io_in_x444_argOut_port_0_bits(RootController_kernelRootController_concrete1_io_in_x444_argOut_port_0_bits),
    .io_in_x423_argOut_port_0_valid(RootController_kernelRootController_concrete1_io_in_x423_argOut_port_0_valid),
    .io_in_x423_argOut_port_0_bits(RootController_kernelRootController_concrete1_io_in_x423_argOut_port_0_bits),
    .io_in_x445_argOut_port_0_valid(RootController_kernelRootController_concrete1_io_in_x445_argOut_port_0_valid),
    .io_in_x445_argOut_port_0_bits(RootController_kernelRootController_concrete1_io_in_x445_argOut_port_0_bits),
    .io_in_x451_argOut_port_0_valid(RootController_kernelRootController_concrete1_io_in_x451_argOut_port_0_valid),
    .io_in_x451_argOut_port_0_bits(RootController_kernelRootController_concrete1_io_in_x451_argOut_port_0_bits),
    .io_in_x434_argOut_port_0_valid(RootController_kernelRootController_concrete1_io_in_x434_argOut_port_0_valid),
    .io_in_x434_argOut_port_0_bits(RootController_kernelRootController_concrete1_io_in_x434_argOut_port_0_bits),
    .io_in_x438_argOut_port_0_valid(RootController_kernelRootController_concrete1_io_in_x438_argOut_port_0_valid),
    .io_in_x438_argOut_port_0_bits(RootController_kernelRootController_concrete1_io_in_x438_argOut_port_0_bits),
    .io_in_x431_argOut_port_0_valid(RootController_kernelRootController_concrete1_io_in_x431_argOut_port_0_valid),
    .io_in_x431_argOut_port_0_bits(RootController_kernelRootController_concrete1_io_in_x431_argOut_port_0_bits),
    .io_in_x426_argOut_port_0_valid(RootController_kernelRootController_concrete1_io_in_x426_argOut_port_0_valid),
    .io_in_x426_argOut_port_0_bits(RootController_kernelRootController_concrete1_io_in_x426_argOut_port_0_bits),
    .io_in_x441_argOut_port_0_valid(RootController_kernelRootController_concrete1_io_in_x441_argOut_port_0_valid),
    .io_in_x441_argOut_port_0_bits(RootController_kernelRootController_concrete1_io_in_x441_argOut_port_0_bits),
    .io_in_x446_argOut_port_0_valid(RootController_kernelRootController_concrete1_io_in_x446_argOut_port_0_valid),
    .io_in_x446_argOut_port_0_bits(RootController_kernelRootController_concrete1_io_in_x446_argOut_port_0_bits),
    .io_in_x450_argOut_port_0_valid(RootController_kernelRootController_concrete1_io_in_x450_argOut_port_0_valid),
    .io_in_x450_argOut_port_0_bits(RootController_kernelRootController_concrete1_io_in_x450_argOut_port_0_bits),
    .io_in_x433_argOut_port_0_valid(RootController_kernelRootController_concrete1_io_in_x433_argOut_port_0_valid),
    .io_in_x433_argOut_port_0_bits(RootController_kernelRootController_concrete1_io_in_x433_argOut_port_0_bits),
    .io_in_x447_argOut_port_0_valid(RootController_kernelRootController_concrete1_io_in_x447_argOut_port_0_valid),
    .io_in_x447_argOut_port_0_bits(RootController_kernelRootController_concrete1_io_in_x447_argOut_port_0_bits),
    .io_in_x432_argOut_port_0_valid(RootController_kernelRootController_concrete1_io_in_x432_argOut_port_0_valid),
    .io_in_x432_argOut_port_0_bits(RootController_kernelRootController_concrete1_io_in_x432_argOut_port_0_bits),
    .io_in_x422_argOut_port_0_valid(RootController_kernelRootController_concrete1_io_in_x422_argOut_port_0_valid),
    .io_in_x422_argOut_port_0_bits(RootController_kernelRootController_concrete1_io_in_x422_argOut_port_0_bits),
    .io_in_x437_argOut_port_0_valid(RootController_kernelRootController_concrete1_io_in_x437_argOut_port_0_valid),
    .io_in_x437_argOut_port_0_bits(RootController_kernelRootController_concrete1_io_in_x437_argOut_port_0_bits),
    .io_in_x427_argOut_port_0_valid(RootController_kernelRootController_concrete1_io_in_x427_argOut_port_0_valid),
    .io_in_x427_argOut_port_0_bits(RootController_kernelRootController_concrete1_io_in_x427_argOut_port_0_bits),
    .io_in_x442_argOut_port_0_valid(RootController_kernelRootController_concrete1_io_in_x442_argOut_port_0_valid),
    .io_in_x442_argOut_port_0_bits(RootController_kernelRootController_concrete1_io_in_x442_argOut_port_0_bits),
    .io_sigsIn_smEnableOuts_0(RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smChildAcks_0(RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsOut_smDoneIn_0(RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_1),
    .io_rr(RootController_kernelRootController_concrete1_io_rr)
  );
  assign _T_1539 = RetimeWrapper_io_out; // @[package.scala 96:25:@7699.4 package.scala 96:25:@7700.4]
  assign _T_1604 = io_enable & _T_1539; // @[Main.scala 194:50:@7779.4]
  assign _T_1605 = ~ SRFF_io_output; // @[Main.scala 194:59:@7780.4]
  assign _T_1617 = RootController_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@7800.4]
  assign io_done = SRFF_io_output; // @[Main.scala 201:23:@7799.4]
  assign io_memStreams_loads_0_cmd_valid = 1'h0;
  assign io_memStreams_loads_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_loads_0_cmd_bits_size = 32'h0;
  assign io_memStreams_loads_0_data_ready = 1'h0;
  assign io_memStreams_stores_0_cmd_valid = 1'h0;
  assign io_memStreams_stores_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_stores_0_cmd_bits_size = 32'h0;
  assign io_memStreams_stores_0_data_valid = 1'h0;
  assign io_memStreams_stores_0_data_bits_wdata_0 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_1 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_2 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_3 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_4 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_5 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_6 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_7 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_8 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_9 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_10 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_11 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_12 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_13 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_14 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_15 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wstrb = 16'h0;
  assign io_memStreams_stores_0_wresp_ready = 1'h0;
  assign io_memStreams_gathers_0_cmd_valid = 1'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_0 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_1 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_2 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_3 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_4 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_5 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_6 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_7 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_8 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_9 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_10 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_11 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_12 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_13 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_14 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_15 = 64'h0;
  assign io_memStreams_gathers_0_data_ready = 1'h0;
  assign io_memStreams_scatters_0_cmd_valid = 1'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_0 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_1 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_2 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_3 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_4 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_5 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_6 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_7 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_8 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_9 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_10 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_11 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_12 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_13 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_14 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_15 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_0 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_1 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_2 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_3 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_4 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_5 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_6 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_7 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_8 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_9 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_10 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_11 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_12 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_13 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_14 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_15 = 32'h0;
  assign io_memStreams_scatters_0_wresp_ready = 1'h0;
  assign io_axiStreamsIn_0_TREADY = RootController_kernelRootController_concrete1_io_in_x416_TREADY; // @[sm_RootController.scala 119:23:@8044.4]
  assign io_axiStreamsOut_0_TVALID = 1'h0;
  assign io_axiStreamsOut_0_TDATA = 256'h0;
  assign io_axiStreamsOut_0_TSTRB = 32'h0;
  assign io_axiStreamsOut_0_TKEEP = 32'h0;
  assign io_axiStreamsOut_0_TLAST = 1'h0;
  assign io_axiStreamsOut_0_TID = 8'h0;
  assign io_axiStreamsOut_0_TDEST = 8'h0;
  assign io_heap_0_req_valid = 1'h0;
  assign io_heap_0_req_bits_allocDealloc = 1'h0;
  assign io_heap_0_req_bits_sizeAddr = 64'h0;
  assign io_argOuts_0_port_valid = RootController_kernelRootController_concrete1_io_in_x420_argOut_port_0_valid; // @[Main.scala 29:69:@7424.4]
  assign io_argOuts_0_port_bits = RootController_kernelRootController_concrete1_io_in_x420_argOut_port_0_bits; // @[Main.scala 30:68:@7425.4]
  assign io_argOuts_1_port_valid = RootController_kernelRootController_concrete1_io_in_x421_argOut_port_0_valid; // @[Main.scala 34:69:@7432.4]
  assign io_argOuts_1_port_bits = RootController_kernelRootController_concrete1_io_in_x421_argOut_port_0_bits; // @[Main.scala 35:68:@7433.4]
  assign io_argOuts_2_port_valid = RootController_kernelRootController_concrete1_io_in_x422_argOut_port_0_valid; // @[Main.scala 39:69:@7440.4]
  assign io_argOuts_2_port_bits = RootController_kernelRootController_concrete1_io_in_x422_argOut_port_0_bits; // @[Main.scala 40:68:@7441.4]
  assign io_argOuts_3_port_valid = RootController_kernelRootController_concrete1_io_in_x423_argOut_port_0_valid; // @[Main.scala 44:69:@7448.4]
  assign io_argOuts_3_port_bits = RootController_kernelRootController_concrete1_io_in_x423_argOut_port_0_bits; // @[Main.scala 45:68:@7449.4]
  assign io_argOuts_4_port_valid = RootController_kernelRootController_concrete1_io_in_x424_argOut_port_0_valid; // @[Main.scala 49:69:@7456.4]
  assign io_argOuts_4_port_bits = RootController_kernelRootController_concrete1_io_in_x424_argOut_port_0_bits; // @[Main.scala 50:68:@7457.4]
  assign io_argOuts_5_port_valid = RootController_kernelRootController_concrete1_io_in_x425_argOut_port_0_valid; // @[Main.scala 54:69:@7464.4]
  assign io_argOuts_5_port_bits = RootController_kernelRootController_concrete1_io_in_x425_argOut_port_0_bits; // @[Main.scala 55:68:@7465.4]
  assign io_argOuts_6_port_valid = RootController_kernelRootController_concrete1_io_in_x426_argOut_port_0_valid; // @[Main.scala 59:69:@7472.4]
  assign io_argOuts_6_port_bits = RootController_kernelRootController_concrete1_io_in_x426_argOut_port_0_bits; // @[Main.scala 60:68:@7473.4]
  assign io_argOuts_7_port_valid = RootController_kernelRootController_concrete1_io_in_x427_argOut_port_0_valid; // @[Main.scala 64:69:@7480.4]
  assign io_argOuts_7_port_bits = RootController_kernelRootController_concrete1_io_in_x427_argOut_port_0_bits; // @[Main.scala 65:68:@7481.4]
  assign io_argOuts_8_port_valid = RootController_kernelRootController_concrete1_io_in_x428_argOut_port_0_valid; // @[Main.scala 69:69:@7488.4]
  assign io_argOuts_8_port_bits = RootController_kernelRootController_concrete1_io_in_x428_argOut_port_0_bits; // @[Main.scala 70:68:@7489.4]
  assign io_argOuts_9_port_valid = RootController_kernelRootController_concrete1_io_in_x429_argOut_port_0_valid; // @[Main.scala 74:69:@7496.4]
  assign io_argOuts_9_port_bits = RootController_kernelRootController_concrete1_io_in_x429_argOut_port_0_bits; // @[Main.scala 75:68:@7497.4]
  assign io_argOuts_10_port_valid = RootController_kernelRootController_concrete1_io_in_x430_argOut_port_0_valid; // @[Main.scala 79:70:@7504.4]
  assign io_argOuts_10_port_bits = RootController_kernelRootController_concrete1_io_in_x430_argOut_port_0_bits; // @[Main.scala 80:69:@7505.4]
  assign io_argOuts_11_port_valid = RootController_kernelRootController_concrete1_io_in_x431_argOut_port_0_valid; // @[Main.scala 84:70:@7512.4]
  assign io_argOuts_11_port_bits = RootController_kernelRootController_concrete1_io_in_x431_argOut_port_0_bits; // @[Main.scala 85:69:@7513.4]
  assign io_argOuts_12_port_valid = RootController_kernelRootController_concrete1_io_in_x432_argOut_port_0_valid; // @[Main.scala 89:70:@7520.4]
  assign io_argOuts_12_port_bits = RootController_kernelRootController_concrete1_io_in_x432_argOut_port_0_bits; // @[Main.scala 90:69:@7521.4]
  assign io_argOuts_13_port_valid = RootController_kernelRootController_concrete1_io_in_x433_argOut_port_0_valid; // @[Main.scala 94:70:@7528.4]
  assign io_argOuts_13_port_bits = RootController_kernelRootController_concrete1_io_in_x433_argOut_port_0_bits; // @[Main.scala 95:69:@7529.4]
  assign io_argOuts_14_port_valid = RootController_kernelRootController_concrete1_io_in_x434_argOut_port_0_valid; // @[Main.scala 99:70:@7536.4]
  assign io_argOuts_14_port_bits = RootController_kernelRootController_concrete1_io_in_x434_argOut_port_0_bits; // @[Main.scala 100:69:@7537.4]
  assign io_argOuts_15_port_valid = RootController_kernelRootController_concrete1_io_in_x435_argOut_port_0_valid; // @[Main.scala 104:70:@7544.4]
  assign io_argOuts_15_port_bits = RootController_kernelRootController_concrete1_io_in_x435_argOut_port_0_bits; // @[Main.scala 105:69:@7545.4]
  assign io_argOuts_16_port_valid = RootController_kernelRootController_concrete1_io_in_x436_argOut_port_0_valid; // @[Main.scala 109:70:@7552.4]
  assign io_argOuts_16_port_bits = RootController_kernelRootController_concrete1_io_in_x436_argOut_port_0_bits; // @[Main.scala 110:69:@7553.4]
  assign io_argOuts_17_port_valid = RootController_kernelRootController_concrete1_io_in_x437_argOut_port_0_valid; // @[Main.scala 114:70:@7560.4]
  assign io_argOuts_17_port_bits = RootController_kernelRootController_concrete1_io_in_x437_argOut_port_0_bits; // @[Main.scala 115:69:@7561.4]
  assign io_argOuts_18_port_valid = RootController_kernelRootController_concrete1_io_in_x438_argOut_port_0_valid; // @[Main.scala 119:70:@7568.4]
  assign io_argOuts_18_port_bits = RootController_kernelRootController_concrete1_io_in_x438_argOut_port_0_bits; // @[Main.scala 120:69:@7569.4]
  assign io_argOuts_19_port_valid = RootController_kernelRootController_concrete1_io_in_x439_argOut_port_0_valid; // @[Main.scala 124:70:@7576.4]
  assign io_argOuts_19_port_bits = RootController_kernelRootController_concrete1_io_in_x439_argOut_port_0_bits; // @[Main.scala 125:69:@7577.4]
  assign io_argOuts_20_port_valid = RootController_kernelRootController_concrete1_io_in_x440_argOut_port_0_valid; // @[Main.scala 129:70:@7584.4]
  assign io_argOuts_20_port_bits = RootController_kernelRootController_concrete1_io_in_x440_argOut_port_0_bits; // @[Main.scala 130:69:@7585.4]
  assign io_argOuts_21_port_valid = RootController_kernelRootController_concrete1_io_in_x441_argOut_port_0_valid; // @[Main.scala 134:70:@7592.4]
  assign io_argOuts_21_port_bits = RootController_kernelRootController_concrete1_io_in_x441_argOut_port_0_bits; // @[Main.scala 135:69:@7593.4]
  assign io_argOuts_22_port_valid = RootController_kernelRootController_concrete1_io_in_x442_argOut_port_0_valid; // @[Main.scala 139:70:@7600.4]
  assign io_argOuts_22_port_bits = RootController_kernelRootController_concrete1_io_in_x442_argOut_port_0_bits; // @[Main.scala 140:69:@7601.4]
  assign io_argOuts_23_port_valid = RootController_kernelRootController_concrete1_io_in_x443_argOut_port_0_valid; // @[Main.scala 144:70:@7608.4]
  assign io_argOuts_23_port_bits = RootController_kernelRootController_concrete1_io_in_x443_argOut_port_0_bits; // @[Main.scala 145:69:@7609.4]
  assign io_argOuts_24_port_valid = RootController_kernelRootController_concrete1_io_in_x444_argOut_port_0_valid; // @[Main.scala 149:70:@7616.4]
  assign io_argOuts_24_port_bits = RootController_kernelRootController_concrete1_io_in_x444_argOut_port_0_bits; // @[Main.scala 150:69:@7617.4]
  assign io_argOuts_25_port_valid = RootController_kernelRootController_concrete1_io_in_x445_argOut_port_0_valid; // @[Main.scala 154:70:@7624.4]
  assign io_argOuts_25_port_bits = RootController_kernelRootController_concrete1_io_in_x445_argOut_port_0_bits; // @[Main.scala 155:69:@7625.4]
  assign io_argOuts_26_port_valid = RootController_kernelRootController_concrete1_io_in_x446_argOut_port_0_valid; // @[Main.scala 159:70:@7632.4]
  assign io_argOuts_26_port_bits = RootController_kernelRootController_concrete1_io_in_x446_argOut_port_0_bits; // @[Main.scala 160:69:@7633.4]
  assign io_argOuts_27_port_valid = RootController_kernelRootController_concrete1_io_in_x447_argOut_port_0_valid; // @[Main.scala 164:70:@7640.4]
  assign io_argOuts_27_port_bits = RootController_kernelRootController_concrete1_io_in_x447_argOut_port_0_bits; // @[Main.scala 165:69:@7641.4]
  assign io_argOuts_28_port_valid = RootController_kernelRootController_concrete1_io_in_x448_argOut_port_0_valid; // @[Main.scala 169:70:@7648.4]
  assign io_argOuts_28_port_bits = RootController_kernelRootController_concrete1_io_in_x448_argOut_port_0_bits; // @[Main.scala 170:69:@7649.4]
  assign io_argOuts_29_port_valid = RootController_kernelRootController_concrete1_io_in_x449_argOut_port_0_valid; // @[Main.scala 174:70:@7656.4]
  assign io_argOuts_29_port_bits = RootController_kernelRootController_concrete1_io_in_x449_argOut_port_0_bits; // @[Main.scala 175:69:@7657.4]
  assign io_argOuts_30_port_valid = RootController_kernelRootController_concrete1_io_in_x450_argOut_port_0_valid; // @[Main.scala 179:70:@7664.4]
  assign io_argOuts_30_port_bits = RootController_kernelRootController_concrete1_io_in_x450_argOut_port_0_bits; // @[Main.scala 180:69:@7665.4]
  assign io_argOuts_31_port_valid = RootController_kernelRootController_concrete1_io_in_x451_argOut_port_0_valid; // @[Main.scala 184:70:@7672.4]
  assign io_argOuts_31_port_bits = RootController_kernelRootController_concrete1_io_in_x451_argOut_port_0_bits; // @[Main.scala 185:69:@7673.4]
  assign SingleCounter_clock = clock; // @[:@7677.4]
  assign SingleCounter_reset = reset; // @[:@7678.4]
  assign SingleCounter_io_input_reset = reset; // @[Main.scala 189:79:@7692.4]
  assign RetimeWrapper_clock = clock; // @[:@7695.4]
  assign RetimeWrapper_reset = reset; // @[:@7696.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@7698.4]
  assign RetimeWrapper_io_in = SingleCounter_io_output_done; // @[package.scala 94:16:@7697.4]
  assign SRFF_clock = clock; // @[:@7704.4]
  assign SRFF_reset = reset; // @[:@7705.4]
  assign SRFF_io_input_set = RootController_sm_io_done; // @[Main.scala 210:29:@8217.4]
  assign SRFF_io_input_reset = RetimeWrapper_1_io_out; // @[Main.scala 199:31:@7797.4]
  assign SRFF_io_input_asyn_reset = RetimeWrapper_1_io_out; // @[Main.scala 200:36:@7798.4]
  assign RootController_sm_clock = clock; // @[:@7747.4]
  assign RootController_sm_reset = reset; // @[:@7748.4]
  assign RootController_sm_io_enable = _T_1604 & _T_1605; // @[Main.scala 198:33:@7796.4 SpatialBlocks.scala 112:18:@7835.4]
  assign RootController_sm_io_rst = RetimeWrapper_1_io_out; // @[SpatialBlocks.scala 106:15:@7829.4]
  assign RootController_sm_io_ctrDone = RootController_sm_io_ctrInc & _T_1620; // @[Main.scala 202:34:@7804.4]
  assign RootController_sm_io_doneIn_0 = RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 102:67:@7824.4]
  assign RootController_sm_io_doneIn_1 = RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 102:67:@7825.4]
  assign RetimeWrapper_1_clock = clock; // @[:@7784.4]
  assign RetimeWrapper_1_reset = reset; // @[:@7785.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@7787.4]
  assign RetimeWrapper_1_io_in = reset | io_reset; // @[package.scala 94:16:@7786.4]
  assign RootController_kernelRootController_concrete1_clock = clock; // @[:@7848.4]
  assign RootController_kernelRootController_concrete1_reset = reset; // @[:@7849.4]
  assign RootController_kernelRootController_concrete1_io_in_x416_TVALID = io_axiStreamsIn_0_TVALID; // @[sm_RootController.scala 119:23:@8045.4]
  assign RootController_kernelRootController_concrete1_io_in_x416_TDATA = io_axiStreamsIn_0_TDATA; // @[sm_RootController.scala 119:23:@8043.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0 = RootController_sm_io_enableOut_0; // @[sm_RootController.scala 240:22:@8196.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_1 = RootController_sm_io_enableOut_1; // @[sm_RootController.scala 240:22:@8197.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0 = RootController_sm_io_childAck_0; // @[sm_RootController.scala 240:22:@8192.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_1 = RootController_sm_io_childAck_1; // @[sm_RootController.scala 240:22:@8193.4]
  assign RootController_kernelRootController_concrete1_io_rr = RetimeWrapper_io_out; // @[sm_RootController.scala 239:18:@8186.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1620 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_1620 <= 1'h0;
    end else begin
      _T_1620 <= _T_1617;
    end
  end
endmodule
module DRAMHeap( // @[:@9124.2]
  input         io_accel_0_req_valid, // @[:@9127.4]
  input         io_accel_0_req_bits_allocDealloc, // @[:@9127.4]
  input  [63:0] io_accel_0_req_bits_sizeAddr, // @[:@9127.4]
  output        io_accel_0_resp_valid, // @[:@9127.4]
  output        io_accel_0_resp_bits_allocDealloc, // @[:@9127.4]
  output [63:0] io_accel_0_resp_bits_sizeAddr, // @[:@9127.4]
  output        io_host_0_req_valid, // @[:@9127.4]
  output        io_host_0_req_bits_allocDealloc, // @[:@9127.4]
  output [63:0] io_host_0_req_bits_sizeAddr, // @[:@9127.4]
  input         io_host_0_resp_valid, // @[:@9127.4]
  input         io_host_0_resp_bits_allocDealloc, // @[:@9127.4]
  input  [63:0] io_host_0_resp_bits_sizeAddr // @[:@9127.4]
);
  assign io_accel_0_resp_valid = io_host_0_resp_valid; // @[DRAMHeap.scala 24:18:@9134.4]
  assign io_accel_0_resp_bits_allocDealloc = io_host_0_resp_bits_allocDealloc; // @[DRAMHeap.scala 25:17:@9136.4]
  assign io_accel_0_resp_bits_sizeAddr = io_host_0_resp_bits_sizeAddr; // @[DRAMHeap.scala 25:17:@9135.4]
  assign io_host_0_req_valid = io_accel_0_req_valid; // @[DRAMHeap.scala 21:18:@9131.4]
  assign io_host_0_req_bits_allocDealloc = io_accel_0_req_bits_allocDealloc; // @[DRAMHeap.scala 21:18:@9130.4]
  assign io_host_0_req_bits_sizeAddr = io_accel_0_req_bits_sizeAddr; // @[DRAMHeap.scala 21:18:@9129.4]
endmodule
module RetimeWrapper_80( // @[:@9150.2]
  input         clock, // @[:@9151.4]
  input         reset, // @[:@9152.4]
  input         io_flow, // @[:@9153.4]
  input  [63:0] io_in, // @[:@9153.4]
  output [63:0] io_out // @[:@9153.4]
);
  wire [63:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@9155.4]
  wire [63:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@9155.4]
  wire [63:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@9155.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@9155.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@9155.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@9155.4]
  RetimeShiftRegister #(.WIDTH(64), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@9155.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@9168.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@9167.4]
  assign sr_init = 64'h0; // @[RetimeShiftRegister.scala 19:16:@9166.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@9165.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@9164.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@9162.4]
endmodule
module FringeFF( // @[:@9170.2]
  input         clock, // @[:@9171.4]
  input         reset, // @[:@9172.4]
  input  [63:0] io_in, // @[:@9173.4]
  input         io_reset, // @[:@9173.4]
  output [63:0] io_out, // @[:@9173.4]
  input         io_enable // @[:@9173.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@9176.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@9176.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@9176.4]
  wire [63:0] RetimeWrapper_io_in; // @[package.scala 93:22:@9176.4]
  wire [63:0] RetimeWrapper_io_out; // @[package.scala 93:22:@9176.4]
  wire [63:0] _T_18; // @[package.scala 96:25:@9181.4 package.scala 96:25:@9182.4]
  wire [63:0] _GEN_0; // @[FringeFF.scala 21:27:@9187.6]
  RetimeWrapper_80 RetimeWrapper ( // @[package.scala 93:22:@9176.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@9181.4 package.scala 96:25:@9182.4]
  assign _GEN_0 = io_reset ? 64'h0 : _T_18; // @[FringeFF.scala 21:27:@9187.6]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@9193.4]
  assign RetimeWrapper_clock = clock; // @[:@9177.4]
  assign RetimeWrapper_reset = reset; // @[:@9178.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@9180.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _GEN_0; // @[package.scala 94:16:@9179.4]
endmodule
module MuxN( // @[:@39576.2]
  input  [63:0] io_ins_0, // @[:@39579.4]
  input  [63:0] io_ins_1, // @[:@39579.4]
  input  [63:0] io_ins_2, // @[:@39579.4]
  input  [63:0] io_ins_3, // @[:@39579.4]
  input  [63:0] io_ins_4, // @[:@39579.4]
  input  [63:0] io_ins_5, // @[:@39579.4]
  input  [63:0] io_ins_6, // @[:@39579.4]
  input  [63:0] io_ins_7, // @[:@39579.4]
  input  [63:0] io_ins_8, // @[:@39579.4]
  input  [63:0] io_ins_9, // @[:@39579.4]
  input  [63:0] io_ins_10, // @[:@39579.4]
  input  [63:0] io_ins_11, // @[:@39579.4]
  input  [63:0] io_ins_12, // @[:@39579.4]
  input  [63:0] io_ins_13, // @[:@39579.4]
  input  [63:0] io_ins_14, // @[:@39579.4]
  input  [63:0] io_ins_15, // @[:@39579.4]
  input  [63:0] io_ins_16, // @[:@39579.4]
  input  [63:0] io_ins_17, // @[:@39579.4]
  input  [63:0] io_ins_18, // @[:@39579.4]
  input  [63:0] io_ins_19, // @[:@39579.4]
  input  [63:0] io_ins_20, // @[:@39579.4]
  input  [63:0] io_ins_21, // @[:@39579.4]
  input  [63:0] io_ins_22, // @[:@39579.4]
  input  [63:0] io_ins_23, // @[:@39579.4]
  input  [63:0] io_ins_24, // @[:@39579.4]
  input  [63:0] io_ins_25, // @[:@39579.4]
  input  [63:0] io_ins_26, // @[:@39579.4]
  input  [63:0] io_ins_27, // @[:@39579.4]
  input  [63:0] io_ins_28, // @[:@39579.4]
  input  [63:0] io_ins_29, // @[:@39579.4]
  input  [63:0] io_ins_30, // @[:@39579.4]
  input  [63:0] io_ins_31, // @[:@39579.4]
  input  [63:0] io_ins_32, // @[:@39579.4]
  input  [63:0] io_ins_33, // @[:@39579.4]
  input  [63:0] io_ins_34, // @[:@39579.4]
  input  [63:0] io_ins_35, // @[:@39579.4]
  input  [63:0] io_ins_36, // @[:@39579.4]
  input  [63:0] io_ins_37, // @[:@39579.4]
  input  [63:0] io_ins_38, // @[:@39579.4]
  input  [63:0] io_ins_39, // @[:@39579.4]
  input  [63:0] io_ins_40, // @[:@39579.4]
  input  [63:0] io_ins_41, // @[:@39579.4]
  input  [63:0] io_ins_42, // @[:@39579.4]
  input  [63:0] io_ins_43, // @[:@39579.4]
  input  [63:0] io_ins_44, // @[:@39579.4]
  input  [63:0] io_ins_45, // @[:@39579.4]
  input  [63:0] io_ins_46, // @[:@39579.4]
  input  [63:0] io_ins_47, // @[:@39579.4]
  input  [63:0] io_ins_48, // @[:@39579.4]
  input  [63:0] io_ins_49, // @[:@39579.4]
  input  [63:0] io_ins_50, // @[:@39579.4]
  input  [63:0] io_ins_51, // @[:@39579.4]
  input  [63:0] io_ins_52, // @[:@39579.4]
  input  [63:0] io_ins_53, // @[:@39579.4]
  input  [63:0] io_ins_54, // @[:@39579.4]
  input  [63:0] io_ins_55, // @[:@39579.4]
  input  [63:0] io_ins_56, // @[:@39579.4]
  input  [63:0] io_ins_57, // @[:@39579.4]
  input  [63:0] io_ins_58, // @[:@39579.4]
  input  [63:0] io_ins_59, // @[:@39579.4]
  input  [63:0] io_ins_60, // @[:@39579.4]
  input  [63:0] io_ins_61, // @[:@39579.4]
  input  [63:0] io_ins_62, // @[:@39579.4]
  input  [63:0] io_ins_63, // @[:@39579.4]
  input  [63:0] io_ins_64, // @[:@39579.4]
  input  [63:0] io_ins_65, // @[:@39579.4]
  input  [63:0] io_ins_66, // @[:@39579.4]
  input  [63:0] io_ins_67, // @[:@39579.4]
  input  [63:0] io_ins_68, // @[:@39579.4]
  input  [63:0] io_ins_69, // @[:@39579.4]
  input  [63:0] io_ins_70, // @[:@39579.4]
  input  [63:0] io_ins_71, // @[:@39579.4]
  input  [63:0] io_ins_72, // @[:@39579.4]
  input  [63:0] io_ins_73, // @[:@39579.4]
  input  [63:0] io_ins_74, // @[:@39579.4]
  input  [63:0] io_ins_75, // @[:@39579.4]
  input  [63:0] io_ins_76, // @[:@39579.4]
  input  [63:0] io_ins_77, // @[:@39579.4]
  input  [63:0] io_ins_78, // @[:@39579.4]
  input  [63:0] io_ins_79, // @[:@39579.4]
  input  [63:0] io_ins_80, // @[:@39579.4]
  input  [63:0] io_ins_81, // @[:@39579.4]
  input  [63:0] io_ins_82, // @[:@39579.4]
  input  [63:0] io_ins_83, // @[:@39579.4]
  input  [63:0] io_ins_84, // @[:@39579.4]
  input  [63:0] io_ins_85, // @[:@39579.4]
  input  [63:0] io_ins_86, // @[:@39579.4]
  input  [63:0] io_ins_87, // @[:@39579.4]
  input  [63:0] io_ins_88, // @[:@39579.4]
  input  [63:0] io_ins_89, // @[:@39579.4]
  input  [63:0] io_ins_90, // @[:@39579.4]
  input  [63:0] io_ins_91, // @[:@39579.4]
  input  [63:0] io_ins_92, // @[:@39579.4]
  input  [63:0] io_ins_93, // @[:@39579.4]
  input  [63:0] io_ins_94, // @[:@39579.4]
  input  [63:0] io_ins_95, // @[:@39579.4]
  input  [63:0] io_ins_96, // @[:@39579.4]
  input  [63:0] io_ins_97, // @[:@39579.4]
  input  [63:0] io_ins_98, // @[:@39579.4]
  input  [63:0] io_ins_99, // @[:@39579.4]
  input  [63:0] io_ins_100, // @[:@39579.4]
  input  [63:0] io_ins_101, // @[:@39579.4]
  input  [63:0] io_ins_102, // @[:@39579.4]
  input  [63:0] io_ins_103, // @[:@39579.4]
  input  [63:0] io_ins_104, // @[:@39579.4]
  input  [63:0] io_ins_105, // @[:@39579.4]
  input  [63:0] io_ins_106, // @[:@39579.4]
  input  [63:0] io_ins_107, // @[:@39579.4]
  input  [63:0] io_ins_108, // @[:@39579.4]
  input  [63:0] io_ins_109, // @[:@39579.4]
  input  [63:0] io_ins_110, // @[:@39579.4]
  input  [63:0] io_ins_111, // @[:@39579.4]
  input  [63:0] io_ins_112, // @[:@39579.4]
  input  [63:0] io_ins_113, // @[:@39579.4]
  input  [63:0] io_ins_114, // @[:@39579.4]
  input  [63:0] io_ins_115, // @[:@39579.4]
  input  [63:0] io_ins_116, // @[:@39579.4]
  input  [63:0] io_ins_117, // @[:@39579.4]
  input  [63:0] io_ins_118, // @[:@39579.4]
  input  [63:0] io_ins_119, // @[:@39579.4]
  input  [63:0] io_ins_120, // @[:@39579.4]
  input  [63:0] io_ins_121, // @[:@39579.4]
  input  [63:0] io_ins_122, // @[:@39579.4]
  input  [63:0] io_ins_123, // @[:@39579.4]
  input  [63:0] io_ins_124, // @[:@39579.4]
  input  [63:0] io_ins_125, // @[:@39579.4]
  input  [63:0] io_ins_126, // @[:@39579.4]
  input  [63:0] io_ins_127, // @[:@39579.4]
  input  [63:0] io_ins_128, // @[:@39579.4]
  input  [63:0] io_ins_129, // @[:@39579.4]
  input  [63:0] io_ins_130, // @[:@39579.4]
  input  [63:0] io_ins_131, // @[:@39579.4]
  input  [63:0] io_ins_132, // @[:@39579.4]
  input  [63:0] io_ins_133, // @[:@39579.4]
  input  [63:0] io_ins_134, // @[:@39579.4]
  input  [63:0] io_ins_135, // @[:@39579.4]
  input  [63:0] io_ins_136, // @[:@39579.4]
  input  [63:0] io_ins_137, // @[:@39579.4]
  input  [63:0] io_ins_138, // @[:@39579.4]
  input  [63:0] io_ins_139, // @[:@39579.4]
  input  [63:0] io_ins_140, // @[:@39579.4]
  input  [63:0] io_ins_141, // @[:@39579.4]
  input  [63:0] io_ins_142, // @[:@39579.4]
  input  [63:0] io_ins_143, // @[:@39579.4]
  input  [63:0] io_ins_144, // @[:@39579.4]
  input  [63:0] io_ins_145, // @[:@39579.4]
  input  [63:0] io_ins_146, // @[:@39579.4]
  input  [63:0] io_ins_147, // @[:@39579.4]
  input  [63:0] io_ins_148, // @[:@39579.4]
  input  [63:0] io_ins_149, // @[:@39579.4]
  input  [63:0] io_ins_150, // @[:@39579.4]
  input  [63:0] io_ins_151, // @[:@39579.4]
  input  [63:0] io_ins_152, // @[:@39579.4]
  input  [63:0] io_ins_153, // @[:@39579.4]
  input  [63:0] io_ins_154, // @[:@39579.4]
  input  [63:0] io_ins_155, // @[:@39579.4]
  input  [63:0] io_ins_156, // @[:@39579.4]
  input  [63:0] io_ins_157, // @[:@39579.4]
  input  [63:0] io_ins_158, // @[:@39579.4]
  input  [63:0] io_ins_159, // @[:@39579.4]
  input  [63:0] io_ins_160, // @[:@39579.4]
  input  [63:0] io_ins_161, // @[:@39579.4]
  input  [63:0] io_ins_162, // @[:@39579.4]
  input  [63:0] io_ins_163, // @[:@39579.4]
  input  [63:0] io_ins_164, // @[:@39579.4]
  input  [63:0] io_ins_165, // @[:@39579.4]
  input  [63:0] io_ins_166, // @[:@39579.4]
  input  [63:0] io_ins_167, // @[:@39579.4]
  input  [63:0] io_ins_168, // @[:@39579.4]
  input  [63:0] io_ins_169, // @[:@39579.4]
  input  [63:0] io_ins_170, // @[:@39579.4]
  input  [63:0] io_ins_171, // @[:@39579.4]
  input  [63:0] io_ins_172, // @[:@39579.4]
  input  [63:0] io_ins_173, // @[:@39579.4]
  input  [63:0] io_ins_174, // @[:@39579.4]
  input  [63:0] io_ins_175, // @[:@39579.4]
  input  [63:0] io_ins_176, // @[:@39579.4]
  input  [63:0] io_ins_177, // @[:@39579.4]
  input  [63:0] io_ins_178, // @[:@39579.4]
  input  [63:0] io_ins_179, // @[:@39579.4]
  input  [63:0] io_ins_180, // @[:@39579.4]
  input  [63:0] io_ins_181, // @[:@39579.4]
  input  [63:0] io_ins_182, // @[:@39579.4]
  input  [63:0] io_ins_183, // @[:@39579.4]
  input  [63:0] io_ins_184, // @[:@39579.4]
  input  [63:0] io_ins_185, // @[:@39579.4]
  input  [63:0] io_ins_186, // @[:@39579.4]
  input  [63:0] io_ins_187, // @[:@39579.4]
  input  [63:0] io_ins_188, // @[:@39579.4]
  input  [63:0] io_ins_189, // @[:@39579.4]
  input  [63:0] io_ins_190, // @[:@39579.4]
  input  [63:0] io_ins_191, // @[:@39579.4]
  input  [63:0] io_ins_192, // @[:@39579.4]
  input  [63:0] io_ins_193, // @[:@39579.4]
  input  [63:0] io_ins_194, // @[:@39579.4]
  input  [63:0] io_ins_195, // @[:@39579.4]
  input  [63:0] io_ins_196, // @[:@39579.4]
  input  [63:0] io_ins_197, // @[:@39579.4]
  input  [63:0] io_ins_198, // @[:@39579.4]
  input  [63:0] io_ins_199, // @[:@39579.4]
  input  [63:0] io_ins_200, // @[:@39579.4]
  input  [63:0] io_ins_201, // @[:@39579.4]
  input  [63:0] io_ins_202, // @[:@39579.4]
  input  [63:0] io_ins_203, // @[:@39579.4]
  input  [63:0] io_ins_204, // @[:@39579.4]
  input  [63:0] io_ins_205, // @[:@39579.4]
  input  [63:0] io_ins_206, // @[:@39579.4]
  input  [63:0] io_ins_207, // @[:@39579.4]
  input  [63:0] io_ins_208, // @[:@39579.4]
  input  [63:0] io_ins_209, // @[:@39579.4]
  input  [63:0] io_ins_210, // @[:@39579.4]
  input  [63:0] io_ins_211, // @[:@39579.4]
  input  [63:0] io_ins_212, // @[:@39579.4]
  input  [63:0] io_ins_213, // @[:@39579.4]
  input  [63:0] io_ins_214, // @[:@39579.4]
  input  [63:0] io_ins_215, // @[:@39579.4]
  input  [63:0] io_ins_216, // @[:@39579.4]
  input  [63:0] io_ins_217, // @[:@39579.4]
  input  [63:0] io_ins_218, // @[:@39579.4]
  input  [63:0] io_ins_219, // @[:@39579.4]
  input  [63:0] io_ins_220, // @[:@39579.4]
  input  [63:0] io_ins_221, // @[:@39579.4]
  input  [63:0] io_ins_222, // @[:@39579.4]
  input  [63:0] io_ins_223, // @[:@39579.4]
  input  [63:0] io_ins_224, // @[:@39579.4]
  input  [63:0] io_ins_225, // @[:@39579.4]
  input  [63:0] io_ins_226, // @[:@39579.4]
  input  [63:0] io_ins_227, // @[:@39579.4]
  input  [63:0] io_ins_228, // @[:@39579.4]
  input  [63:0] io_ins_229, // @[:@39579.4]
  input  [63:0] io_ins_230, // @[:@39579.4]
  input  [63:0] io_ins_231, // @[:@39579.4]
  input  [63:0] io_ins_232, // @[:@39579.4]
  input  [63:0] io_ins_233, // @[:@39579.4]
  input  [63:0] io_ins_234, // @[:@39579.4]
  input  [63:0] io_ins_235, // @[:@39579.4]
  input  [63:0] io_ins_236, // @[:@39579.4]
  input  [63:0] io_ins_237, // @[:@39579.4]
  input  [63:0] io_ins_238, // @[:@39579.4]
  input  [63:0] io_ins_239, // @[:@39579.4]
  input  [63:0] io_ins_240, // @[:@39579.4]
  input  [63:0] io_ins_241, // @[:@39579.4]
  input  [63:0] io_ins_242, // @[:@39579.4]
  input  [63:0] io_ins_243, // @[:@39579.4]
  input  [63:0] io_ins_244, // @[:@39579.4]
  input  [63:0] io_ins_245, // @[:@39579.4]
  input  [63:0] io_ins_246, // @[:@39579.4]
  input  [63:0] io_ins_247, // @[:@39579.4]
  input  [63:0] io_ins_248, // @[:@39579.4]
  input  [63:0] io_ins_249, // @[:@39579.4]
  input  [63:0] io_ins_250, // @[:@39579.4]
  input  [63:0] io_ins_251, // @[:@39579.4]
  input  [63:0] io_ins_252, // @[:@39579.4]
  input  [63:0] io_ins_253, // @[:@39579.4]
  input  [63:0] io_ins_254, // @[:@39579.4]
  input  [63:0] io_ins_255, // @[:@39579.4]
  input  [63:0] io_ins_256, // @[:@39579.4]
  input  [63:0] io_ins_257, // @[:@39579.4]
  input  [63:0] io_ins_258, // @[:@39579.4]
  input  [63:0] io_ins_259, // @[:@39579.4]
  input  [63:0] io_ins_260, // @[:@39579.4]
  input  [63:0] io_ins_261, // @[:@39579.4]
  input  [63:0] io_ins_262, // @[:@39579.4]
  input  [63:0] io_ins_263, // @[:@39579.4]
  input  [63:0] io_ins_264, // @[:@39579.4]
  input  [63:0] io_ins_265, // @[:@39579.4]
  input  [63:0] io_ins_266, // @[:@39579.4]
  input  [63:0] io_ins_267, // @[:@39579.4]
  input  [63:0] io_ins_268, // @[:@39579.4]
  input  [63:0] io_ins_269, // @[:@39579.4]
  input  [63:0] io_ins_270, // @[:@39579.4]
  input  [63:0] io_ins_271, // @[:@39579.4]
  input  [63:0] io_ins_272, // @[:@39579.4]
  input  [63:0] io_ins_273, // @[:@39579.4]
  input  [63:0] io_ins_274, // @[:@39579.4]
  input  [63:0] io_ins_275, // @[:@39579.4]
  input  [63:0] io_ins_276, // @[:@39579.4]
  input  [63:0] io_ins_277, // @[:@39579.4]
  input  [63:0] io_ins_278, // @[:@39579.4]
  input  [63:0] io_ins_279, // @[:@39579.4]
  input  [63:0] io_ins_280, // @[:@39579.4]
  input  [63:0] io_ins_281, // @[:@39579.4]
  input  [63:0] io_ins_282, // @[:@39579.4]
  input  [63:0] io_ins_283, // @[:@39579.4]
  input  [63:0] io_ins_284, // @[:@39579.4]
  input  [63:0] io_ins_285, // @[:@39579.4]
  input  [63:0] io_ins_286, // @[:@39579.4]
  input  [63:0] io_ins_287, // @[:@39579.4]
  input  [63:0] io_ins_288, // @[:@39579.4]
  input  [63:0] io_ins_289, // @[:@39579.4]
  input  [63:0] io_ins_290, // @[:@39579.4]
  input  [63:0] io_ins_291, // @[:@39579.4]
  input  [63:0] io_ins_292, // @[:@39579.4]
  input  [63:0] io_ins_293, // @[:@39579.4]
  input  [63:0] io_ins_294, // @[:@39579.4]
  input  [63:0] io_ins_295, // @[:@39579.4]
  input  [63:0] io_ins_296, // @[:@39579.4]
  input  [63:0] io_ins_297, // @[:@39579.4]
  input  [63:0] io_ins_298, // @[:@39579.4]
  input  [63:0] io_ins_299, // @[:@39579.4]
  input  [63:0] io_ins_300, // @[:@39579.4]
  input  [63:0] io_ins_301, // @[:@39579.4]
  input  [63:0] io_ins_302, // @[:@39579.4]
  input  [63:0] io_ins_303, // @[:@39579.4]
  input  [63:0] io_ins_304, // @[:@39579.4]
  input  [63:0] io_ins_305, // @[:@39579.4]
  input  [63:0] io_ins_306, // @[:@39579.4]
  input  [63:0] io_ins_307, // @[:@39579.4]
  input  [63:0] io_ins_308, // @[:@39579.4]
  input  [63:0] io_ins_309, // @[:@39579.4]
  input  [63:0] io_ins_310, // @[:@39579.4]
  input  [63:0] io_ins_311, // @[:@39579.4]
  input  [63:0] io_ins_312, // @[:@39579.4]
  input  [63:0] io_ins_313, // @[:@39579.4]
  input  [63:0] io_ins_314, // @[:@39579.4]
  input  [63:0] io_ins_315, // @[:@39579.4]
  input  [63:0] io_ins_316, // @[:@39579.4]
  input  [63:0] io_ins_317, // @[:@39579.4]
  input  [63:0] io_ins_318, // @[:@39579.4]
  input  [63:0] io_ins_319, // @[:@39579.4]
  input  [63:0] io_ins_320, // @[:@39579.4]
  input  [63:0] io_ins_321, // @[:@39579.4]
  input  [63:0] io_ins_322, // @[:@39579.4]
  input  [63:0] io_ins_323, // @[:@39579.4]
  input  [63:0] io_ins_324, // @[:@39579.4]
  input  [63:0] io_ins_325, // @[:@39579.4]
  input  [63:0] io_ins_326, // @[:@39579.4]
  input  [63:0] io_ins_327, // @[:@39579.4]
  input  [63:0] io_ins_328, // @[:@39579.4]
  input  [63:0] io_ins_329, // @[:@39579.4]
  input  [63:0] io_ins_330, // @[:@39579.4]
  input  [63:0] io_ins_331, // @[:@39579.4]
  input  [63:0] io_ins_332, // @[:@39579.4]
  input  [63:0] io_ins_333, // @[:@39579.4]
  input  [63:0] io_ins_334, // @[:@39579.4]
  input  [63:0] io_ins_335, // @[:@39579.4]
  input  [63:0] io_ins_336, // @[:@39579.4]
  input  [63:0] io_ins_337, // @[:@39579.4]
  input  [63:0] io_ins_338, // @[:@39579.4]
  input  [63:0] io_ins_339, // @[:@39579.4]
  input  [63:0] io_ins_340, // @[:@39579.4]
  input  [63:0] io_ins_341, // @[:@39579.4]
  input  [63:0] io_ins_342, // @[:@39579.4]
  input  [63:0] io_ins_343, // @[:@39579.4]
  input  [63:0] io_ins_344, // @[:@39579.4]
  input  [63:0] io_ins_345, // @[:@39579.4]
  input  [63:0] io_ins_346, // @[:@39579.4]
  input  [63:0] io_ins_347, // @[:@39579.4]
  input  [63:0] io_ins_348, // @[:@39579.4]
  input  [63:0] io_ins_349, // @[:@39579.4]
  input  [63:0] io_ins_350, // @[:@39579.4]
  input  [63:0] io_ins_351, // @[:@39579.4]
  input  [63:0] io_ins_352, // @[:@39579.4]
  input  [63:0] io_ins_353, // @[:@39579.4]
  input  [63:0] io_ins_354, // @[:@39579.4]
  input  [63:0] io_ins_355, // @[:@39579.4]
  input  [63:0] io_ins_356, // @[:@39579.4]
  input  [63:0] io_ins_357, // @[:@39579.4]
  input  [63:0] io_ins_358, // @[:@39579.4]
  input  [63:0] io_ins_359, // @[:@39579.4]
  input  [63:0] io_ins_360, // @[:@39579.4]
  input  [63:0] io_ins_361, // @[:@39579.4]
  input  [63:0] io_ins_362, // @[:@39579.4]
  input  [63:0] io_ins_363, // @[:@39579.4]
  input  [63:0] io_ins_364, // @[:@39579.4]
  input  [63:0] io_ins_365, // @[:@39579.4]
  input  [63:0] io_ins_366, // @[:@39579.4]
  input  [63:0] io_ins_367, // @[:@39579.4]
  input  [63:0] io_ins_368, // @[:@39579.4]
  input  [63:0] io_ins_369, // @[:@39579.4]
  input  [63:0] io_ins_370, // @[:@39579.4]
  input  [63:0] io_ins_371, // @[:@39579.4]
  input  [63:0] io_ins_372, // @[:@39579.4]
  input  [63:0] io_ins_373, // @[:@39579.4]
  input  [63:0] io_ins_374, // @[:@39579.4]
  input  [63:0] io_ins_375, // @[:@39579.4]
  input  [63:0] io_ins_376, // @[:@39579.4]
  input  [63:0] io_ins_377, // @[:@39579.4]
  input  [63:0] io_ins_378, // @[:@39579.4]
  input  [63:0] io_ins_379, // @[:@39579.4]
  input  [63:0] io_ins_380, // @[:@39579.4]
  input  [63:0] io_ins_381, // @[:@39579.4]
  input  [63:0] io_ins_382, // @[:@39579.4]
  input  [63:0] io_ins_383, // @[:@39579.4]
  input  [63:0] io_ins_384, // @[:@39579.4]
  input  [63:0] io_ins_385, // @[:@39579.4]
  input  [63:0] io_ins_386, // @[:@39579.4]
  input  [63:0] io_ins_387, // @[:@39579.4]
  input  [63:0] io_ins_388, // @[:@39579.4]
  input  [63:0] io_ins_389, // @[:@39579.4]
  input  [63:0] io_ins_390, // @[:@39579.4]
  input  [63:0] io_ins_391, // @[:@39579.4]
  input  [63:0] io_ins_392, // @[:@39579.4]
  input  [63:0] io_ins_393, // @[:@39579.4]
  input  [63:0] io_ins_394, // @[:@39579.4]
  input  [63:0] io_ins_395, // @[:@39579.4]
  input  [63:0] io_ins_396, // @[:@39579.4]
  input  [63:0] io_ins_397, // @[:@39579.4]
  input  [63:0] io_ins_398, // @[:@39579.4]
  input  [63:0] io_ins_399, // @[:@39579.4]
  input  [63:0] io_ins_400, // @[:@39579.4]
  input  [63:0] io_ins_401, // @[:@39579.4]
  input  [63:0] io_ins_402, // @[:@39579.4]
  input  [63:0] io_ins_403, // @[:@39579.4]
  input  [63:0] io_ins_404, // @[:@39579.4]
  input  [63:0] io_ins_405, // @[:@39579.4]
  input  [63:0] io_ins_406, // @[:@39579.4]
  input  [63:0] io_ins_407, // @[:@39579.4]
  input  [63:0] io_ins_408, // @[:@39579.4]
  input  [63:0] io_ins_409, // @[:@39579.4]
  input  [63:0] io_ins_410, // @[:@39579.4]
  input  [63:0] io_ins_411, // @[:@39579.4]
  input  [63:0] io_ins_412, // @[:@39579.4]
  input  [63:0] io_ins_413, // @[:@39579.4]
  input  [63:0] io_ins_414, // @[:@39579.4]
  input  [63:0] io_ins_415, // @[:@39579.4]
  input  [63:0] io_ins_416, // @[:@39579.4]
  input  [63:0] io_ins_417, // @[:@39579.4]
  input  [63:0] io_ins_418, // @[:@39579.4]
  input  [63:0] io_ins_419, // @[:@39579.4]
  input  [63:0] io_ins_420, // @[:@39579.4]
  input  [63:0] io_ins_421, // @[:@39579.4]
  input  [63:0] io_ins_422, // @[:@39579.4]
  input  [63:0] io_ins_423, // @[:@39579.4]
  input  [63:0] io_ins_424, // @[:@39579.4]
  input  [63:0] io_ins_425, // @[:@39579.4]
  input  [63:0] io_ins_426, // @[:@39579.4]
  input  [63:0] io_ins_427, // @[:@39579.4]
  input  [63:0] io_ins_428, // @[:@39579.4]
  input  [63:0] io_ins_429, // @[:@39579.4]
  input  [63:0] io_ins_430, // @[:@39579.4]
  input  [63:0] io_ins_431, // @[:@39579.4]
  input  [63:0] io_ins_432, // @[:@39579.4]
  input  [63:0] io_ins_433, // @[:@39579.4]
  input  [63:0] io_ins_434, // @[:@39579.4]
  input  [63:0] io_ins_435, // @[:@39579.4]
  input  [63:0] io_ins_436, // @[:@39579.4]
  input  [63:0] io_ins_437, // @[:@39579.4]
  input  [63:0] io_ins_438, // @[:@39579.4]
  input  [63:0] io_ins_439, // @[:@39579.4]
  input  [63:0] io_ins_440, // @[:@39579.4]
  input  [63:0] io_ins_441, // @[:@39579.4]
  input  [63:0] io_ins_442, // @[:@39579.4]
  input  [63:0] io_ins_443, // @[:@39579.4]
  input  [63:0] io_ins_444, // @[:@39579.4]
  input  [63:0] io_ins_445, // @[:@39579.4]
  input  [63:0] io_ins_446, // @[:@39579.4]
  input  [63:0] io_ins_447, // @[:@39579.4]
  input  [63:0] io_ins_448, // @[:@39579.4]
  input  [63:0] io_ins_449, // @[:@39579.4]
  input  [63:0] io_ins_450, // @[:@39579.4]
  input  [63:0] io_ins_451, // @[:@39579.4]
  input  [63:0] io_ins_452, // @[:@39579.4]
  input  [63:0] io_ins_453, // @[:@39579.4]
  input  [63:0] io_ins_454, // @[:@39579.4]
  input  [63:0] io_ins_455, // @[:@39579.4]
  input  [63:0] io_ins_456, // @[:@39579.4]
  input  [63:0] io_ins_457, // @[:@39579.4]
  input  [63:0] io_ins_458, // @[:@39579.4]
  input  [63:0] io_ins_459, // @[:@39579.4]
  input  [63:0] io_ins_460, // @[:@39579.4]
  input  [63:0] io_ins_461, // @[:@39579.4]
  input  [63:0] io_ins_462, // @[:@39579.4]
  input  [63:0] io_ins_463, // @[:@39579.4]
  input  [63:0] io_ins_464, // @[:@39579.4]
  input  [63:0] io_ins_465, // @[:@39579.4]
  input  [63:0] io_ins_466, // @[:@39579.4]
  input  [63:0] io_ins_467, // @[:@39579.4]
  input  [63:0] io_ins_468, // @[:@39579.4]
  input  [63:0] io_ins_469, // @[:@39579.4]
  input  [63:0] io_ins_470, // @[:@39579.4]
  input  [63:0] io_ins_471, // @[:@39579.4]
  input  [63:0] io_ins_472, // @[:@39579.4]
  input  [63:0] io_ins_473, // @[:@39579.4]
  input  [63:0] io_ins_474, // @[:@39579.4]
  input  [63:0] io_ins_475, // @[:@39579.4]
  input  [63:0] io_ins_476, // @[:@39579.4]
  input  [63:0] io_ins_477, // @[:@39579.4]
  input  [63:0] io_ins_478, // @[:@39579.4]
  input  [63:0] io_ins_479, // @[:@39579.4]
  input  [63:0] io_ins_480, // @[:@39579.4]
  input  [63:0] io_ins_481, // @[:@39579.4]
  input  [63:0] io_ins_482, // @[:@39579.4]
  input  [63:0] io_ins_483, // @[:@39579.4]
  input  [63:0] io_ins_484, // @[:@39579.4]
  input  [63:0] io_ins_485, // @[:@39579.4]
  input  [63:0] io_ins_486, // @[:@39579.4]
  input  [63:0] io_ins_487, // @[:@39579.4]
  input  [63:0] io_ins_488, // @[:@39579.4]
  input  [63:0] io_ins_489, // @[:@39579.4]
  input  [63:0] io_ins_490, // @[:@39579.4]
  input  [63:0] io_ins_491, // @[:@39579.4]
  input  [63:0] io_ins_492, // @[:@39579.4]
  input  [63:0] io_ins_493, // @[:@39579.4]
  input  [63:0] io_ins_494, // @[:@39579.4]
  input  [63:0] io_ins_495, // @[:@39579.4]
  input  [63:0] io_ins_496, // @[:@39579.4]
  input  [63:0] io_ins_497, // @[:@39579.4]
  input  [63:0] io_ins_498, // @[:@39579.4]
  input  [63:0] io_ins_499, // @[:@39579.4]
  input  [63:0] io_ins_500, // @[:@39579.4]
  input  [63:0] io_ins_501, // @[:@39579.4]
  input  [63:0] io_ins_502, // @[:@39579.4]
  input  [63:0] io_ins_503, // @[:@39579.4]
  input  [63:0] io_ins_504, // @[:@39579.4]
  input  [63:0] io_ins_505, // @[:@39579.4]
  input  [63:0] io_ins_506, // @[:@39579.4]
  input  [63:0] io_ins_507, // @[:@39579.4]
  input  [63:0] io_ins_508, // @[:@39579.4]
  input  [63:0] io_ins_509, // @[:@39579.4]
  input  [63:0] io_ins_510, // @[:@39579.4]
  input  [63:0] io_ins_511, // @[:@39579.4]
  input  [63:0] io_ins_512, // @[:@39579.4]
  input  [63:0] io_ins_513, // @[:@39579.4]
  input  [63:0] io_ins_514, // @[:@39579.4]
  input  [63:0] io_ins_515, // @[:@39579.4]
  input  [63:0] io_ins_516, // @[:@39579.4]
  input  [63:0] io_ins_517, // @[:@39579.4]
  input  [63:0] io_ins_518, // @[:@39579.4]
  input  [63:0] io_ins_519, // @[:@39579.4]
  input  [63:0] io_ins_520, // @[:@39579.4]
  input  [63:0] io_ins_521, // @[:@39579.4]
  input  [63:0] io_ins_522, // @[:@39579.4]
  input  [63:0] io_ins_523, // @[:@39579.4]
  input  [63:0] io_ins_524, // @[:@39579.4]
  input  [63:0] io_ins_525, // @[:@39579.4]
  input  [63:0] io_ins_526, // @[:@39579.4]
  input  [63:0] io_ins_527, // @[:@39579.4]
  input  [63:0] io_ins_528, // @[:@39579.4]
  input  [63:0] io_ins_529, // @[:@39579.4]
  input  [63:0] io_ins_530, // @[:@39579.4]
  input  [63:0] io_ins_531, // @[:@39579.4]
  input  [63:0] io_ins_532, // @[:@39579.4]
  input  [63:0] io_ins_533, // @[:@39579.4]
  input  [9:0]  io_sel, // @[:@39579.4]
  output [63:0] io_out // @[:@39579.4]
);
  wire [63:0] _GEN_1; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_2; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_3; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_4; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_5; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_6; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_7; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_8; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_9; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_10; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_11; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_12; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_13; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_14; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_15; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_16; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_17; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_18; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_19; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_20; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_21; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_22; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_23; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_24; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_25; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_26; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_27; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_28; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_29; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_30; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_31; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_32; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_33; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_34; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_35; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_36; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_37; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_38; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_39; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_40; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_41; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_42; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_43; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_44; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_45; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_46; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_47; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_48; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_49; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_50; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_51; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_52; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_53; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_54; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_55; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_56; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_57; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_58; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_59; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_60; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_61; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_62; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_63; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_64; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_65; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_66; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_67; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_68; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_69; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_70; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_71; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_72; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_73; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_74; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_75; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_76; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_77; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_78; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_79; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_80; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_81; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_82; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_83; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_84; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_85; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_86; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_87; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_88; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_89; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_90; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_91; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_92; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_93; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_94; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_95; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_96; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_97; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_98; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_99; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_100; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_101; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_102; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_103; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_104; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_105; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_106; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_107; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_108; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_109; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_110; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_111; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_112; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_113; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_114; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_115; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_116; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_117; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_118; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_119; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_120; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_121; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_122; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_123; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_124; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_125; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_126; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_127; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_128; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_129; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_130; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_131; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_132; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_133; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_134; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_135; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_136; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_137; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_138; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_139; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_140; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_141; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_142; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_143; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_144; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_145; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_146; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_147; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_148; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_149; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_150; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_151; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_152; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_153; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_154; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_155; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_156; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_157; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_158; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_159; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_160; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_161; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_162; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_163; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_164; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_165; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_166; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_167; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_168; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_169; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_170; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_171; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_172; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_173; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_174; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_175; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_176; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_177; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_178; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_179; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_180; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_181; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_182; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_183; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_184; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_185; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_186; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_187; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_188; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_189; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_190; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_191; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_192; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_193; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_194; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_195; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_196; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_197; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_198; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_199; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_200; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_201; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_202; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_203; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_204; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_205; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_206; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_207; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_208; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_209; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_210; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_211; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_212; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_213; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_214; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_215; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_216; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_217; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_218; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_219; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_220; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_221; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_222; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_223; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_224; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_225; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_226; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_227; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_228; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_229; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_230; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_231; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_232; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_233; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_234; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_235; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_236; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_237; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_238; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_239; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_240; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_241; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_242; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_243; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_244; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_245; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_246; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_247; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_248; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_249; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_250; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_251; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_252; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_253; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_254; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_255; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_256; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_257; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_258; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_259; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_260; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_261; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_262; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_263; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_264; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_265; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_266; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_267; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_268; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_269; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_270; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_271; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_272; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_273; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_274; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_275; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_276; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_277; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_278; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_279; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_280; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_281; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_282; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_283; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_284; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_285; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_286; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_287; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_288; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_289; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_290; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_291; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_292; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_293; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_294; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_295; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_296; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_297; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_298; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_299; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_300; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_301; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_302; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_303; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_304; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_305; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_306; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_307; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_308; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_309; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_310; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_311; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_312; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_313; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_314; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_315; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_316; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_317; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_318; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_319; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_320; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_321; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_322; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_323; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_324; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_325; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_326; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_327; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_328; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_329; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_330; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_331; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_332; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_333; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_334; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_335; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_336; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_337; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_338; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_339; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_340; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_341; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_342; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_343; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_344; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_345; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_346; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_347; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_348; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_349; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_350; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_351; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_352; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_353; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_354; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_355; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_356; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_357; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_358; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_359; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_360; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_361; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_362; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_363; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_364; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_365; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_366; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_367; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_368; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_369; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_370; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_371; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_372; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_373; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_374; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_375; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_376; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_377; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_378; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_379; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_380; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_381; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_382; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_383; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_384; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_385; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_386; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_387; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_388; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_389; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_390; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_391; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_392; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_393; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_394; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_395; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_396; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_397; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_398; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_399; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_400; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_401; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_402; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_403; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_404; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_405; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_406; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_407; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_408; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_409; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_410; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_411; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_412; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_413; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_414; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_415; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_416; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_417; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_418; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_419; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_420; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_421; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_422; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_423; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_424; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_425; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_426; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_427; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_428; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_429; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_430; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_431; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_432; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_433; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_434; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_435; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_436; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_437; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_438; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_439; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_440; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_441; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_442; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_443; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_444; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_445; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_446; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_447; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_448; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_449; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_450; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_451; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_452; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_453; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_454; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_455; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_456; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_457; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_458; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_459; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_460; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_461; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_462; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_463; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_464; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_465; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_466; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_467; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_468; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_469; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_470; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_471; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_472; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_473; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_474; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_475; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_476; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_477; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_478; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_479; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_480; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_481; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_482; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_483; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_484; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_485; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_486; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_487; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_488; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_489; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_490; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_491; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_492; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_493; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_494; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_495; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_496; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_497; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_498; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_499; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_500; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_501; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_502; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_503; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_504; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_505; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_506; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_507; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_508; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_509; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_510; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_511; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_512; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_513; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_514; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_515; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_516; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_517; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_518; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_519; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_520; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_521; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_522; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_523; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_524; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_525; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_526; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_527; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_528; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_529; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_530; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_531; // @[MuxN.scala 16:10:@39581.4]
  wire [63:0] _GEN_532; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_1 = 10'h1 == io_sel ? io_ins_1 : io_ins_0; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_2 = 10'h2 == io_sel ? io_ins_2 : _GEN_1; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_3 = 10'h3 == io_sel ? io_ins_3 : _GEN_2; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_4 = 10'h4 == io_sel ? io_ins_4 : _GEN_3; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_5 = 10'h5 == io_sel ? io_ins_5 : _GEN_4; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_6 = 10'h6 == io_sel ? io_ins_6 : _GEN_5; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_7 = 10'h7 == io_sel ? io_ins_7 : _GEN_6; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_8 = 10'h8 == io_sel ? io_ins_8 : _GEN_7; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_9 = 10'h9 == io_sel ? io_ins_9 : _GEN_8; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_10 = 10'ha == io_sel ? io_ins_10 : _GEN_9; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_11 = 10'hb == io_sel ? io_ins_11 : _GEN_10; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_12 = 10'hc == io_sel ? io_ins_12 : _GEN_11; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_13 = 10'hd == io_sel ? io_ins_13 : _GEN_12; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_14 = 10'he == io_sel ? io_ins_14 : _GEN_13; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_15 = 10'hf == io_sel ? io_ins_15 : _GEN_14; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_16 = 10'h10 == io_sel ? io_ins_16 : _GEN_15; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_17 = 10'h11 == io_sel ? io_ins_17 : _GEN_16; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_18 = 10'h12 == io_sel ? io_ins_18 : _GEN_17; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_19 = 10'h13 == io_sel ? io_ins_19 : _GEN_18; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_20 = 10'h14 == io_sel ? io_ins_20 : _GEN_19; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_21 = 10'h15 == io_sel ? io_ins_21 : _GEN_20; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_22 = 10'h16 == io_sel ? io_ins_22 : _GEN_21; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_23 = 10'h17 == io_sel ? io_ins_23 : _GEN_22; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_24 = 10'h18 == io_sel ? io_ins_24 : _GEN_23; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_25 = 10'h19 == io_sel ? io_ins_25 : _GEN_24; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_26 = 10'h1a == io_sel ? io_ins_26 : _GEN_25; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_27 = 10'h1b == io_sel ? io_ins_27 : _GEN_26; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_28 = 10'h1c == io_sel ? io_ins_28 : _GEN_27; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_29 = 10'h1d == io_sel ? io_ins_29 : _GEN_28; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_30 = 10'h1e == io_sel ? io_ins_30 : _GEN_29; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_31 = 10'h1f == io_sel ? io_ins_31 : _GEN_30; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_32 = 10'h20 == io_sel ? io_ins_32 : _GEN_31; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_33 = 10'h21 == io_sel ? io_ins_33 : _GEN_32; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_34 = 10'h22 == io_sel ? io_ins_34 : _GEN_33; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_35 = 10'h23 == io_sel ? io_ins_35 : _GEN_34; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_36 = 10'h24 == io_sel ? io_ins_36 : _GEN_35; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_37 = 10'h25 == io_sel ? io_ins_37 : _GEN_36; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_38 = 10'h26 == io_sel ? io_ins_38 : _GEN_37; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_39 = 10'h27 == io_sel ? io_ins_39 : _GEN_38; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_40 = 10'h28 == io_sel ? io_ins_40 : _GEN_39; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_41 = 10'h29 == io_sel ? io_ins_41 : _GEN_40; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_42 = 10'h2a == io_sel ? io_ins_42 : _GEN_41; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_43 = 10'h2b == io_sel ? io_ins_43 : _GEN_42; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_44 = 10'h2c == io_sel ? io_ins_44 : _GEN_43; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_45 = 10'h2d == io_sel ? io_ins_45 : _GEN_44; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_46 = 10'h2e == io_sel ? io_ins_46 : _GEN_45; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_47 = 10'h2f == io_sel ? io_ins_47 : _GEN_46; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_48 = 10'h30 == io_sel ? io_ins_48 : _GEN_47; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_49 = 10'h31 == io_sel ? io_ins_49 : _GEN_48; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_50 = 10'h32 == io_sel ? io_ins_50 : _GEN_49; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_51 = 10'h33 == io_sel ? io_ins_51 : _GEN_50; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_52 = 10'h34 == io_sel ? io_ins_52 : _GEN_51; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_53 = 10'h35 == io_sel ? io_ins_53 : _GEN_52; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_54 = 10'h36 == io_sel ? io_ins_54 : _GEN_53; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_55 = 10'h37 == io_sel ? io_ins_55 : _GEN_54; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_56 = 10'h38 == io_sel ? io_ins_56 : _GEN_55; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_57 = 10'h39 == io_sel ? io_ins_57 : _GEN_56; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_58 = 10'h3a == io_sel ? io_ins_58 : _GEN_57; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_59 = 10'h3b == io_sel ? io_ins_59 : _GEN_58; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_60 = 10'h3c == io_sel ? io_ins_60 : _GEN_59; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_61 = 10'h3d == io_sel ? io_ins_61 : _GEN_60; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_62 = 10'h3e == io_sel ? io_ins_62 : _GEN_61; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_63 = 10'h3f == io_sel ? io_ins_63 : _GEN_62; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_64 = 10'h40 == io_sel ? io_ins_64 : _GEN_63; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_65 = 10'h41 == io_sel ? io_ins_65 : _GEN_64; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_66 = 10'h42 == io_sel ? io_ins_66 : _GEN_65; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_67 = 10'h43 == io_sel ? io_ins_67 : _GEN_66; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_68 = 10'h44 == io_sel ? io_ins_68 : _GEN_67; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_69 = 10'h45 == io_sel ? io_ins_69 : _GEN_68; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_70 = 10'h46 == io_sel ? io_ins_70 : _GEN_69; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_71 = 10'h47 == io_sel ? io_ins_71 : _GEN_70; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_72 = 10'h48 == io_sel ? io_ins_72 : _GEN_71; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_73 = 10'h49 == io_sel ? io_ins_73 : _GEN_72; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_74 = 10'h4a == io_sel ? io_ins_74 : _GEN_73; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_75 = 10'h4b == io_sel ? io_ins_75 : _GEN_74; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_76 = 10'h4c == io_sel ? io_ins_76 : _GEN_75; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_77 = 10'h4d == io_sel ? io_ins_77 : _GEN_76; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_78 = 10'h4e == io_sel ? io_ins_78 : _GEN_77; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_79 = 10'h4f == io_sel ? io_ins_79 : _GEN_78; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_80 = 10'h50 == io_sel ? io_ins_80 : _GEN_79; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_81 = 10'h51 == io_sel ? io_ins_81 : _GEN_80; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_82 = 10'h52 == io_sel ? io_ins_82 : _GEN_81; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_83 = 10'h53 == io_sel ? io_ins_83 : _GEN_82; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_84 = 10'h54 == io_sel ? io_ins_84 : _GEN_83; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_85 = 10'h55 == io_sel ? io_ins_85 : _GEN_84; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_86 = 10'h56 == io_sel ? io_ins_86 : _GEN_85; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_87 = 10'h57 == io_sel ? io_ins_87 : _GEN_86; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_88 = 10'h58 == io_sel ? io_ins_88 : _GEN_87; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_89 = 10'h59 == io_sel ? io_ins_89 : _GEN_88; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_90 = 10'h5a == io_sel ? io_ins_90 : _GEN_89; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_91 = 10'h5b == io_sel ? io_ins_91 : _GEN_90; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_92 = 10'h5c == io_sel ? io_ins_92 : _GEN_91; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_93 = 10'h5d == io_sel ? io_ins_93 : _GEN_92; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_94 = 10'h5e == io_sel ? io_ins_94 : _GEN_93; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_95 = 10'h5f == io_sel ? io_ins_95 : _GEN_94; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_96 = 10'h60 == io_sel ? io_ins_96 : _GEN_95; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_97 = 10'h61 == io_sel ? io_ins_97 : _GEN_96; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_98 = 10'h62 == io_sel ? io_ins_98 : _GEN_97; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_99 = 10'h63 == io_sel ? io_ins_99 : _GEN_98; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_100 = 10'h64 == io_sel ? io_ins_100 : _GEN_99; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_101 = 10'h65 == io_sel ? io_ins_101 : _GEN_100; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_102 = 10'h66 == io_sel ? io_ins_102 : _GEN_101; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_103 = 10'h67 == io_sel ? io_ins_103 : _GEN_102; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_104 = 10'h68 == io_sel ? io_ins_104 : _GEN_103; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_105 = 10'h69 == io_sel ? io_ins_105 : _GEN_104; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_106 = 10'h6a == io_sel ? io_ins_106 : _GEN_105; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_107 = 10'h6b == io_sel ? io_ins_107 : _GEN_106; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_108 = 10'h6c == io_sel ? io_ins_108 : _GEN_107; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_109 = 10'h6d == io_sel ? io_ins_109 : _GEN_108; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_110 = 10'h6e == io_sel ? io_ins_110 : _GEN_109; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_111 = 10'h6f == io_sel ? io_ins_111 : _GEN_110; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_112 = 10'h70 == io_sel ? io_ins_112 : _GEN_111; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_113 = 10'h71 == io_sel ? io_ins_113 : _GEN_112; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_114 = 10'h72 == io_sel ? io_ins_114 : _GEN_113; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_115 = 10'h73 == io_sel ? io_ins_115 : _GEN_114; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_116 = 10'h74 == io_sel ? io_ins_116 : _GEN_115; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_117 = 10'h75 == io_sel ? io_ins_117 : _GEN_116; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_118 = 10'h76 == io_sel ? io_ins_118 : _GEN_117; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_119 = 10'h77 == io_sel ? io_ins_119 : _GEN_118; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_120 = 10'h78 == io_sel ? io_ins_120 : _GEN_119; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_121 = 10'h79 == io_sel ? io_ins_121 : _GEN_120; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_122 = 10'h7a == io_sel ? io_ins_122 : _GEN_121; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_123 = 10'h7b == io_sel ? io_ins_123 : _GEN_122; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_124 = 10'h7c == io_sel ? io_ins_124 : _GEN_123; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_125 = 10'h7d == io_sel ? io_ins_125 : _GEN_124; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_126 = 10'h7e == io_sel ? io_ins_126 : _GEN_125; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_127 = 10'h7f == io_sel ? io_ins_127 : _GEN_126; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_128 = 10'h80 == io_sel ? io_ins_128 : _GEN_127; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_129 = 10'h81 == io_sel ? io_ins_129 : _GEN_128; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_130 = 10'h82 == io_sel ? io_ins_130 : _GEN_129; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_131 = 10'h83 == io_sel ? io_ins_131 : _GEN_130; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_132 = 10'h84 == io_sel ? io_ins_132 : _GEN_131; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_133 = 10'h85 == io_sel ? io_ins_133 : _GEN_132; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_134 = 10'h86 == io_sel ? io_ins_134 : _GEN_133; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_135 = 10'h87 == io_sel ? io_ins_135 : _GEN_134; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_136 = 10'h88 == io_sel ? io_ins_136 : _GEN_135; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_137 = 10'h89 == io_sel ? io_ins_137 : _GEN_136; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_138 = 10'h8a == io_sel ? io_ins_138 : _GEN_137; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_139 = 10'h8b == io_sel ? io_ins_139 : _GEN_138; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_140 = 10'h8c == io_sel ? io_ins_140 : _GEN_139; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_141 = 10'h8d == io_sel ? io_ins_141 : _GEN_140; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_142 = 10'h8e == io_sel ? io_ins_142 : _GEN_141; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_143 = 10'h8f == io_sel ? io_ins_143 : _GEN_142; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_144 = 10'h90 == io_sel ? io_ins_144 : _GEN_143; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_145 = 10'h91 == io_sel ? io_ins_145 : _GEN_144; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_146 = 10'h92 == io_sel ? io_ins_146 : _GEN_145; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_147 = 10'h93 == io_sel ? io_ins_147 : _GEN_146; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_148 = 10'h94 == io_sel ? io_ins_148 : _GEN_147; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_149 = 10'h95 == io_sel ? io_ins_149 : _GEN_148; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_150 = 10'h96 == io_sel ? io_ins_150 : _GEN_149; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_151 = 10'h97 == io_sel ? io_ins_151 : _GEN_150; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_152 = 10'h98 == io_sel ? io_ins_152 : _GEN_151; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_153 = 10'h99 == io_sel ? io_ins_153 : _GEN_152; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_154 = 10'h9a == io_sel ? io_ins_154 : _GEN_153; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_155 = 10'h9b == io_sel ? io_ins_155 : _GEN_154; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_156 = 10'h9c == io_sel ? io_ins_156 : _GEN_155; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_157 = 10'h9d == io_sel ? io_ins_157 : _GEN_156; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_158 = 10'h9e == io_sel ? io_ins_158 : _GEN_157; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_159 = 10'h9f == io_sel ? io_ins_159 : _GEN_158; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_160 = 10'ha0 == io_sel ? io_ins_160 : _GEN_159; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_161 = 10'ha1 == io_sel ? io_ins_161 : _GEN_160; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_162 = 10'ha2 == io_sel ? io_ins_162 : _GEN_161; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_163 = 10'ha3 == io_sel ? io_ins_163 : _GEN_162; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_164 = 10'ha4 == io_sel ? io_ins_164 : _GEN_163; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_165 = 10'ha5 == io_sel ? io_ins_165 : _GEN_164; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_166 = 10'ha6 == io_sel ? io_ins_166 : _GEN_165; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_167 = 10'ha7 == io_sel ? io_ins_167 : _GEN_166; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_168 = 10'ha8 == io_sel ? io_ins_168 : _GEN_167; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_169 = 10'ha9 == io_sel ? io_ins_169 : _GEN_168; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_170 = 10'haa == io_sel ? io_ins_170 : _GEN_169; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_171 = 10'hab == io_sel ? io_ins_171 : _GEN_170; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_172 = 10'hac == io_sel ? io_ins_172 : _GEN_171; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_173 = 10'had == io_sel ? io_ins_173 : _GEN_172; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_174 = 10'hae == io_sel ? io_ins_174 : _GEN_173; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_175 = 10'haf == io_sel ? io_ins_175 : _GEN_174; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_176 = 10'hb0 == io_sel ? io_ins_176 : _GEN_175; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_177 = 10'hb1 == io_sel ? io_ins_177 : _GEN_176; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_178 = 10'hb2 == io_sel ? io_ins_178 : _GEN_177; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_179 = 10'hb3 == io_sel ? io_ins_179 : _GEN_178; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_180 = 10'hb4 == io_sel ? io_ins_180 : _GEN_179; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_181 = 10'hb5 == io_sel ? io_ins_181 : _GEN_180; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_182 = 10'hb6 == io_sel ? io_ins_182 : _GEN_181; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_183 = 10'hb7 == io_sel ? io_ins_183 : _GEN_182; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_184 = 10'hb8 == io_sel ? io_ins_184 : _GEN_183; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_185 = 10'hb9 == io_sel ? io_ins_185 : _GEN_184; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_186 = 10'hba == io_sel ? io_ins_186 : _GEN_185; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_187 = 10'hbb == io_sel ? io_ins_187 : _GEN_186; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_188 = 10'hbc == io_sel ? io_ins_188 : _GEN_187; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_189 = 10'hbd == io_sel ? io_ins_189 : _GEN_188; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_190 = 10'hbe == io_sel ? io_ins_190 : _GEN_189; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_191 = 10'hbf == io_sel ? io_ins_191 : _GEN_190; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_192 = 10'hc0 == io_sel ? io_ins_192 : _GEN_191; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_193 = 10'hc1 == io_sel ? io_ins_193 : _GEN_192; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_194 = 10'hc2 == io_sel ? io_ins_194 : _GEN_193; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_195 = 10'hc3 == io_sel ? io_ins_195 : _GEN_194; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_196 = 10'hc4 == io_sel ? io_ins_196 : _GEN_195; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_197 = 10'hc5 == io_sel ? io_ins_197 : _GEN_196; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_198 = 10'hc6 == io_sel ? io_ins_198 : _GEN_197; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_199 = 10'hc7 == io_sel ? io_ins_199 : _GEN_198; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_200 = 10'hc8 == io_sel ? io_ins_200 : _GEN_199; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_201 = 10'hc9 == io_sel ? io_ins_201 : _GEN_200; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_202 = 10'hca == io_sel ? io_ins_202 : _GEN_201; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_203 = 10'hcb == io_sel ? io_ins_203 : _GEN_202; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_204 = 10'hcc == io_sel ? io_ins_204 : _GEN_203; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_205 = 10'hcd == io_sel ? io_ins_205 : _GEN_204; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_206 = 10'hce == io_sel ? io_ins_206 : _GEN_205; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_207 = 10'hcf == io_sel ? io_ins_207 : _GEN_206; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_208 = 10'hd0 == io_sel ? io_ins_208 : _GEN_207; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_209 = 10'hd1 == io_sel ? io_ins_209 : _GEN_208; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_210 = 10'hd2 == io_sel ? io_ins_210 : _GEN_209; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_211 = 10'hd3 == io_sel ? io_ins_211 : _GEN_210; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_212 = 10'hd4 == io_sel ? io_ins_212 : _GEN_211; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_213 = 10'hd5 == io_sel ? io_ins_213 : _GEN_212; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_214 = 10'hd6 == io_sel ? io_ins_214 : _GEN_213; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_215 = 10'hd7 == io_sel ? io_ins_215 : _GEN_214; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_216 = 10'hd8 == io_sel ? io_ins_216 : _GEN_215; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_217 = 10'hd9 == io_sel ? io_ins_217 : _GEN_216; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_218 = 10'hda == io_sel ? io_ins_218 : _GEN_217; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_219 = 10'hdb == io_sel ? io_ins_219 : _GEN_218; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_220 = 10'hdc == io_sel ? io_ins_220 : _GEN_219; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_221 = 10'hdd == io_sel ? io_ins_221 : _GEN_220; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_222 = 10'hde == io_sel ? io_ins_222 : _GEN_221; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_223 = 10'hdf == io_sel ? io_ins_223 : _GEN_222; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_224 = 10'he0 == io_sel ? io_ins_224 : _GEN_223; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_225 = 10'he1 == io_sel ? io_ins_225 : _GEN_224; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_226 = 10'he2 == io_sel ? io_ins_226 : _GEN_225; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_227 = 10'he3 == io_sel ? io_ins_227 : _GEN_226; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_228 = 10'he4 == io_sel ? io_ins_228 : _GEN_227; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_229 = 10'he5 == io_sel ? io_ins_229 : _GEN_228; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_230 = 10'he6 == io_sel ? io_ins_230 : _GEN_229; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_231 = 10'he7 == io_sel ? io_ins_231 : _GEN_230; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_232 = 10'he8 == io_sel ? io_ins_232 : _GEN_231; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_233 = 10'he9 == io_sel ? io_ins_233 : _GEN_232; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_234 = 10'hea == io_sel ? io_ins_234 : _GEN_233; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_235 = 10'heb == io_sel ? io_ins_235 : _GEN_234; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_236 = 10'hec == io_sel ? io_ins_236 : _GEN_235; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_237 = 10'hed == io_sel ? io_ins_237 : _GEN_236; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_238 = 10'hee == io_sel ? io_ins_238 : _GEN_237; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_239 = 10'hef == io_sel ? io_ins_239 : _GEN_238; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_240 = 10'hf0 == io_sel ? io_ins_240 : _GEN_239; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_241 = 10'hf1 == io_sel ? io_ins_241 : _GEN_240; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_242 = 10'hf2 == io_sel ? io_ins_242 : _GEN_241; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_243 = 10'hf3 == io_sel ? io_ins_243 : _GEN_242; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_244 = 10'hf4 == io_sel ? io_ins_244 : _GEN_243; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_245 = 10'hf5 == io_sel ? io_ins_245 : _GEN_244; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_246 = 10'hf6 == io_sel ? io_ins_246 : _GEN_245; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_247 = 10'hf7 == io_sel ? io_ins_247 : _GEN_246; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_248 = 10'hf8 == io_sel ? io_ins_248 : _GEN_247; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_249 = 10'hf9 == io_sel ? io_ins_249 : _GEN_248; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_250 = 10'hfa == io_sel ? io_ins_250 : _GEN_249; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_251 = 10'hfb == io_sel ? io_ins_251 : _GEN_250; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_252 = 10'hfc == io_sel ? io_ins_252 : _GEN_251; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_253 = 10'hfd == io_sel ? io_ins_253 : _GEN_252; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_254 = 10'hfe == io_sel ? io_ins_254 : _GEN_253; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_255 = 10'hff == io_sel ? io_ins_255 : _GEN_254; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_256 = 10'h100 == io_sel ? io_ins_256 : _GEN_255; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_257 = 10'h101 == io_sel ? io_ins_257 : _GEN_256; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_258 = 10'h102 == io_sel ? io_ins_258 : _GEN_257; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_259 = 10'h103 == io_sel ? io_ins_259 : _GEN_258; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_260 = 10'h104 == io_sel ? io_ins_260 : _GEN_259; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_261 = 10'h105 == io_sel ? io_ins_261 : _GEN_260; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_262 = 10'h106 == io_sel ? io_ins_262 : _GEN_261; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_263 = 10'h107 == io_sel ? io_ins_263 : _GEN_262; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_264 = 10'h108 == io_sel ? io_ins_264 : _GEN_263; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_265 = 10'h109 == io_sel ? io_ins_265 : _GEN_264; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_266 = 10'h10a == io_sel ? io_ins_266 : _GEN_265; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_267 = 10'h10b == io_sel ? io_ins_267 : _GEN_266; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_268 = 10'h10c == io_sel ? io_ins_268 : _GEN_267; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_269 = 10'h10d == io_sel ? io_ins_269 : _GEN_268; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_270 = 10'h10e == io_sel ? io_ins_270 : _GEN_269; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_271 = 10'h10f == io_sel ? io_ins_271 : _GEN_270; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_272 = 10'h110 == io_sel ? io_ins_272 : _GEN_271; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_273 = 10'h111 == io_sel ? io_ins_273 : _GEN_272; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_274 = 10'h112 == io_sel ? io_ins_274 : _GEN_273; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_275 = 10'h113 == io_sel ? io_ins_275 : _GEN_274; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_276 = 10'h114 == io_sel ? io_ins_276 : _GEN_275; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_277 = 10'h115 == io_sel ? io_ins_277 : _GEN_276; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_278 = 10'h116 == io_sel ? io_ins_278 : _GEN_277; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_279 = 10'h117 == io_sel ? io_ins_279 : _GEN_278; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_280 = 10'h118 == io_sel ? io_ins_280 : _GEN_279; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_281 = 10'h119 == io_sel ? io_ins_281 : _GEN_280; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_282 = 10'h11a == io_sel ? io_ins_282 : _GEN_281; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_283 = 10'h11b == io_sel ? io_ins_283 : _GEN_282; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_284 = 10'h11c == io_sel ? io_ins_284 : _GEN_283; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_285 = 10'h11d == io_sel ? io_ins_285 : _GEN_284; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_286 = 10'h11e == io_sel ? io_ins_286 : _GEN_285; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_287 = 10'h11f == io_sel ? io_ins_287 : _GEN_286; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_288 = 10'h120 == io_sel ? io_ins_288 : _GEN_287; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_289 = 10'h121 == io_sel ? io_ins_289 : _GEN_288; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_290 = 10'h122 == io_sel ? io_ins_290 : _GEN_289; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_291 = 10'h123 == io_sel ? io_ins_291 : _GEN_290; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_292 = 10'h124 == io_sel ? io_ins_292 : _GEN_291; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_293 = 10'h125 == io_sel ? io_ins_293 : _GEN_292; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_294 = 10'h126 == io_sel ? io_ins_294 : _GEN_293; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_295 = 10'h127 == io_sel ? io_ins_295 : _GEN_294; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_296 = 10'h128 == io_sel ? io_ins_296 : _GEN_295; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_297 = 10'h129 == io_sel ? io_ins_297 : _GEN_296; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_298 = 10'h12a == io_sel ? io_ins_298 : _GEN_297; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_299 = 10'h12b == io_sel ? io_ins_299 : _GEN_298; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_300 = 10'h12c == io_sel ? io_ins_300 : _GEN_299; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_301 = 10'h12d == io_sel ? io_ins_301 : _GEN_300; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_302 = 10'h12e == io_sel ? io_ins_302 : _GEN_301; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_303 = 10'h12f == io_sel ? io_ins_303 : _GEN_302; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_304 = 10'h130 == io_sel ? io_ins_304 : _GEN_303; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_305 = 10'h131 == io_sel ? io_ins_305 : _GEN_304; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_306 = 10'h132 == io_sel ? io_ins_306 : _GEN_305; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_307 = 10'h133 == io_sel ? io_ins_307 : _GEN_306; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_308 = 10'h134 == io_sel ? io_ins_308 : _GEN_307; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_309 = 10'h135 == io_sel ? io_ins_309 : _GEN_308; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_310 = 10'h136 == io_sel ? io_ins_310 : _GEN_309; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_311 = 10'h137 == io_sel ? io_ins_311 : _GEN_310; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_312 = 10'h138 == io_sel ? io_ins_312 : _GEN_311; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_313 = 10'h139 == io_sel ? io_ins_313 : _GEN_312; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_314 = 10'h13a == io_sel ? io_ins_314 : _GEN_313; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_315 = 10'h13b == io_sel ? io_ins_315 : _GEN_314; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_316 = 10'h13c == io_sel ? io_ins_316 : _GEN_315; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_317 = 10'h13d == io_sel ? io_ins_317 : _GEN_316; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_318 = 10'h13e == io_sel ? io_ins_318 : _GEN_317; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_319 = 10'h13f == io_sel ? io_ins_319 : _GEN_318; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_320 = 10'h140 == io_sel ? io_ins_320 : _GEN_319; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_321 = 10'h141 == io_sel ? io_ins_321 : _GEN_320; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_322 = 10'h142 == io_sel ? io_ins_322 : _GEN_321; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_323 = 10'h143 == io_sel ? io_ins_323 : _GEN_322; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_324 = 10'h144 == io_sel ? io_ins_324 : _GEN_323; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_325 = 10'h145 == io_sel ? io_ins_325 : _GEN_324; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_326 = 10'h146 == io_sel ? io_ins_326 : _GEN_325; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_327 = 10'h147 == io_sel ? io_ins_327 : _GEN_326; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_328 = 10'h148 == io_sel ? io_ins_328 : _GEN_327; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_329 = 10'h149 == io_sel ? io_ins_329 : _GEN_328; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_330 = 10'h14a == io_sel ? io_ins_330 : _GEN_329; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_331 = 10'h14b == io_sel ? io_ins_331 : _GEN_330; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_332 = 10'h14c == io_sel ? io_ins_332 : _GEN_331; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_333 = 10'h14d == io_sel ? io_ins_333 : _GEN_332; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_334 = 10'h14e == io_sel ? io_ins_334 : _GEN_333; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_335 = 10'h14f == io_sel ? io_ins_335 : _GEN_334; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_336 = 10'h150 == io_sel ? io_ins_336 : _GEN_335; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_337 = 10'h151 == io_sel ? io_ins_337 : _GEN_336; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_338 = 10'h152 == io_sel ? io_ins_338 : _GEN_337; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_339 = 10'h153 == io_sel ? io_ins_339 : _GEN_338; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_340 = 10'h154 == io_sel ? io_ins_340 : _GEN_339; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_341 = 10'h155 == io_sel ? io_ins_341 : _GEN_340; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_342 = 10'h156 == io_sel ? io_ins_342 : _GEN_341; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_343 = 10'h157 == io_sel ? io_ins_343 : _GEN_342; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_344 = 10'h158 == io_sel ? io_ins_344 : _GEN_343; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_345 = 10'h159 == io_sel ? io_ins_345 : _GEN_344; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_346 = 10'h15a == io_sel ? io_ins_346 : _GEN_345; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_347 = 10'h15b == io_sel ? io_ins_347 : _GEN_346; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_348 = 10'h15c == io_sel ? io_ins_348 : _GEN_347; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_349 = 10'h15d == io_sel ? io_ins_349 : _GEN_348; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_350 = 10'h15e == io_sel ? io_ins_350 : _GEN_349; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_351 = 10'h15f == io_sel ? io_ins_351 : _GEN_350; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_352 = 10'h160 == io_sel ? io_ins_352 : _GEN_351; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_353 = 10'h161 == io_sel ? io_ins_353 : _GEN_352; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_354 = 10'h162 == io_sel ? io_ins_354 : _GEN_353; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_355 = 10'h163 == io_sel ? io_ins_355 : _GEN_354; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_356 = 10'h164 == io_sel ? io_ins_356 : _GEN_355; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_357 = 10'h165 == io_sel ? io_ins_357 : _GEN_356; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_358 = 10'h166 == io_sel ? io_ins_358 : _GEN_357; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_359 = 10'h167 == io_sel ? io_ins_359 : _GEN_358; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_360 = 10'h168 == io_sel ? io_ins_360 : _GEN_359; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_361 = 10'h169 == io_sel ? io_ins_361 : _GEN_360; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_362 = 10'h16a == io_sel ? io_ins_362 : _GEN_361; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_363 = 10'h16b == io_sel ? io_ins_363 : _GEN_362; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_364 = 10'h16c == io_sel ? io_ins_364 : _GEN_363; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_365 = 10'h16d == io_sel ? io_ins_365 : _GEN_364; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_366 = 10'h16e == io_sel ? io_ins_366 : _GEN_365; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_367 = 10'h16f == io_sel ? io_ins_367 : _GEN_366; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_368 = 10'h170 == io_sel ? io_ins_368 : _GEN_367; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_369 = 10'h171 == io_sel ? io_ins_369 : _GEN_368; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_370 = 10'h172 == io_sel ? io_ins_370 : _GEN_369; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_371 = 10'h173 == io_sel ? io_ins_371 : _GEN_370; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_372 = 10'h174 == io_sel ? io_ins_372 : _GEN_371; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_373 = 10'h175 == io_sel ? io_ins_373 : _GEN_372; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_374 = 10'h176 == io_sel ? io_ins_374 : _GEN_373; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_375 = 10'h177 == io_sel ? io_ins_375 : _GEN_374; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_376 = 10'h178 == io_sel ? io_ins_376 : _GEN_375; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_377 = 10'h179 == io_sel ? io_ins_377 : _GEN_376; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_378 = 10'h17a == io_sel ? io_ins_378 : _GEN_377; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_379 = 10'h17b == io_sel ? io_ins_379 : _GEN_378; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_380 = 10'h17c == io_sel ? io_ins_380 : _GEN_379; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_381 = 10'h17d == io_sel ? io_ins_381 : _GEN_380; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_382 = 10'h17e == io_sel ? io_ins_382 : _GEN_381; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_383 = 10'h17f == io_sel ? io_ins_383 : _GEN_382; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_384 = 10'h180 == io_sel ? io_ins_384 : _GEN_383; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_385 = 10'h181 == io_sel ? io_ins_385 : _GEN_384; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_386 = 10'h182 == io_sel ? io_ins_386 : _GEN_385; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_387 = 10'h183 == io_sel ? io_ins_387 : _GEN_386; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_388 = 10'h184 == io_sel ? io_ins_388 : _GEN_387; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_389 = 10'h185 == io_sel ? io_ins_389 : _GEN_388; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_390 = 10'h186 == io_sel ? io_ins_390 : _GEN_389; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_391 = 10'h187 == io_sel ? io_ins_391 : _GEN_390; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_392 = 10'h188 == io_sel ? io_ins_392 : _GEN_391; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_393 = 10'h189 == io_sel ? io_ins_393 : _GEN_392; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_394 = 10'h18a == io_sel ? io_ins_394 : _GEN_393; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_395 = 10'h18b == io_sel ? io_ins_395 : _GEN_394; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_396 = 10'h18c == io_sel ? io_ins_396 : _GEN_395; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_397 = 10'h18d == io_sel ? io_ins_397 : _GEN_396; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_398 = 10'h18e == io_sel ? io_ins_398 : _GEN_397; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_399 = 10'h18f == io_sel ? io_ins_399 : _GEN_398; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_400 = 10'h190 == io_sel ? io_ins_400 : _GEN_399; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_401 = 10'h191 == io_sel ? io_ins_401 : _GEN_400; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_402 = 10'h192 == io_sel ? io_ins_402 : _GEN_401; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_403 = 10'h193 == io_sel ? io_ins_403 : _GEN_402; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_404 = 10'h194 == io_sel ? io_ins_404 : _GEN_403; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_405 = 10'h195 == io_sel ? io_ins_405 : _GEN_404; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_406 = 10'h196 == io_sel ? io_ins_406 : _GEN_405; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_407 = 10'h197 == io_sel ? io_ins_407 : _GEN_406; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_408 = 10'h198 == io_sel ? io_ins_408 : _GEN_407; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_409 = 10'h199 == io_sel ? io_ins_409 : _GEN_408; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_410 = 10'h19a == io_sel ? io_ins_410 : _GEN_409; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_411 = 10'h19b == io_sel ? io_ins_411 : _GEN_410; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_412 = 10'h19c == io_sel ? io_ins_412 : _GEN_411; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_413 = 10'h19d == io_sel ? io_ins_413 : _GEN_412; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_414 = 10'h19e == io_sel ? io_ins_414 : _GEN_413; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_415 = 10'h19f == io_sel ? io_ins_415 : _GEN_414; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_416 = 10'h1a0 == io_sel ? io_ins_416 : _GEN_415; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_417 = 10'h1a1 == io_sel ? io_ins_417 : _GEN_416; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_418 = 10'h1a2 == io_sel ? io_ins_418 : _GEN_417; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_419 = 10'h1a3 == io_sel ? io_ins_419 : _GEN_418; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_420 = 10'h1a4 == io_sel ? io_ins_420 : _GEN_419; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_421 = 10'h1a5 == io_sel ? io_ins_421 : _GEN_420; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_422 = 10'h1a6 == io_sel ? io_ins_422 : _GEN_421; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_423 = 10'h1a7 == io_sel ? io_ins_423 : _GEN_422; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_424 = 10'h1a8 == io_sel ? io_ins_424 : _GEN_423; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_425 = 10'h1a9 == io_sel ? io_ins_425 : _GEN_424; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_426 = 10'h1aa == io_sel ? io_ins_426 : _GEN_425; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_427 = 10'h1ab == io_sel ? io_ins_427 : _GEN_426; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_428 = 10'h1ac == io_sel ? io_ins_428 : _GEN_427; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_429 = 10'h1ad == io_sel ? io_ins_429 : _GEN_428; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_430 = 10'h1ae == io_sel ? io_ins_430 : _GEN_429; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_431 = 10'h1af == io_sel ? io_ins_431 : _GEN_430; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_432 = 10'h1b0 == io_sel ? io_ins_432 : _GEN_431; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_433 = 10'h1b1 == io_sel ? io_ins_433 : _GEN_432; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_434 = 10'h1b2 == io_sel ? io_ins_434 : _GEN_433; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_435 = 10'h1b3 == io_sel ? io_ins_435 : _GEN_434; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_436 = 10'h1b4 == io_sel ? io_ins_436 : _GEN_435; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_437 = 10'h1b5 == io_sel ? io_ins_437 : _GEN_436; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_438 = 10'h1b6 == io_sel ? io_ins_438 : _GEN_437; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_439 = 10'h1b7 == io_sel ? io_ins_439 : _GEN_438; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_440 = 10'h1b8 == io_sel ? io_ins_440 : _GEN_439; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_441 = 10'h1b9 == io_sel ? io_ins_441 : _GEN_440; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_442 = 10'h1ba == io_sel ? io_ins_442 : _GEN_441; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_443 = 10'h1bb == io_sel ? io_ins_443 : _GEN_442; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_444 = 10'h1bc == io_sel ? io_ins_444 : _GEN_443; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_445 = 10'h1bd == io_sel ? io_ins_445 : _GEN_444; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_446 = 10'h1be == io_sel ? io_ins_446 : _GEN_445; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_447 = 10'h1bf == io_sel ? io_ins_447 : _GEN_446; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_448 = 10'h1c0 == io_sel ? io_ins_448 : _GEN_447; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_449 = 10'h1c1 == io_sel ? io_ins_449 : _GEN_448; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_450 = 10'h1c2 == io_sel ? io_ins_450 : _GEN_449; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_451 = 10'h1c3 == io_sel ? io_ins_451 : _GEN_450; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_452 = 10'h1c4 == io_sel ? io_ins_452 : _GEN_451; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_453 = 10'h1c5 == io_sel ? io_ins_453 : _GEN_452; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_454 = 10'h1c6 == io_sel ? io_ins_454 : _GEN_453; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_455 = 10'h1c7 == io_sel ? io_ins_455 : _GEN_454; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_456 = 10'h1c8 == io_sel ? io_ins_456 : _GEN_455; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_457 = 10'h1c9 == io_sel ? io_ins_457 : _GEN_456; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_458 = 10'h1ca == io_sel ? io_ins_458 : _GEN_457; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_459 = 10'h1cb == io_sel ? io_ins_459 : _GEN_458; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_460 = 10'h1cc == io_sel ? io_ins_460 : _GEN_459; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_461 = 10'h1cd == io_sel ? io_ins_461 : _GEN_460; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_462 = 10'h1ce == io_sel ? io_ins_462 : _GEN_461; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_463 = 10'h1cf == io_sel ? io_ins_463 : _GEN_462; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_464 = 10'h1d0 == io_sel ? io_ins_464 : _GEN_463; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_465 = 10'h1d1 == io_sel ? io_ins_465 : _GEN_464; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_466 = 10'h1d2 == io_sel ? io_ins_466 : _GEN_465; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_467 = 10'h1d3 == io_sel ? io_ins_467 : _GEN_466; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_468 = 10'h1d4 == io_sel ? io_ins_468 : _GEN_467; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_469 = 10'h1d5 == io_sel ? io_ins_469 : _GEN_468; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_470 = 10'h1d6 == io_sel ? io_ins_470 : _GEN_469; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_471 = 10'h1d7 == io_sel ? io_ins_471 : _GEN_470; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_472 = 10'h1d8 == io_sel ? io_ins_472 : _GEN_471; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_473 = 10'h1d9 == io_sel ? io_ins_473 : _GEN_472; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_474 = 10'h1da == io_sel ? io_ins_474 : _GEN_473; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_475 = 10'h1db == io_sel ? io_ins_475 : _GEN_474; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_476 = 10'h1dc == io_sel ? io_ins_476 : _GEN_475; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_477 = 10'h1dd == io_sel ? io_ins_477 : _GEN_476; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_478 = 10'h1de == io_sel ? io_ins_478 : _GEN_477; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_479 = 10'h1df == io_sel ? io_ins_479 : _GEN_478; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_480 = 10'h1e0 == io_sel ? io_ins_480 : _GEN_479; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_481 = 10'h1e1 == io_sel ? io_ins_481 : _GEN_480; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_482 = 10'h1e2 == io_sel ? io_ins_482 : _GEN_481; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_483 = 10'h1e3 == io_sel ? io_ins_483 : _GEN_482; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_484 = 10'h1e4 == io_sel ? io_ins_484 : _GEN_483; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_485 = 10'h1e5 == io_sel ? io_ins_485 : _GEN_484; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_486 = 10'h1e6 == io_sel ? io_ins_486 : _GEN_485; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_487 = 10'h1e7 == io_sel ? io_ins_487 : _GEN_486; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_488 = 10'h1e8 == io_sel ? io_ins_488 : _GEN_487; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_489 = 10'h1e9 == io_sel ? io_ins_489 : _GEN_488; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_490 = 10'h1ea == io_sel ? io_ins_490 : _GEN_489; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_491 = 10'h1eb == io_sel ? io_ins_491 : _GEN_490; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_492 = 10'h1ec == io_sel ? io_ins_492 : _GEN_491; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_493 = 10'h1ed == io_sel ? io_ins_493 : _GEN_492; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_494 = 10'h1ee == io_sel ? io_ins_494 : _GEN_493; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_495 = 10'h1ef == io_sel ? io_ins_495 : _GEN_494; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_496 = 10'h1f0 == io_sel ? io_ins_496 : _GEN_495; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_497 = 10'h1f1 == io_sel ? io_ins_497 : _GEN_496; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_498 = 10'h1f2 == io_sel ? io_ins_498 : _GEN_497; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_499 = 10'h1f3 == io_sel ? io_ins_499 : _GEN_498; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_500 = 10'h1f4 == io_sel ? io_ins_500 : _GEN_499; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_501 = 10'h1f5 == io_sel ? io_ins_501 : _GEN_500; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_502 = 10'h1f6 == io_sel ? io_ins_502 : _GEN_501; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_503 = 10'h1f7 == io_sel ? io_ins_503 : _GEN_502; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_504 = 10'h1f8 == io_sel ? io_ins_504 : _GEN_503; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_505 = 10'h1f9 == io_sel ? io_ins_505 : _GEN_504; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_506 = 10'h1fa == io_sel ? io_ins_506 : _GEN_505; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_507 = 10'h1fb == io_sel ? io_ins_507 : _GEN_506; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_508 = 10'h1fc == io_sel ? io_ins_508 : _GEN_507; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_509 = 10'h1fd == io_sel ? io_ins_509 : _GEN_508; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_510 = 10'h1fe == io_sel ? io_ins_510 : _GEN_509; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_511 = 10'h1ff == io_sel ? io_ins_511 : _GEN_510; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_512 = 10'h200 == io_sel ? io_ins_512 : _GEN_511; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_513 = 10'h201 == io_sel ? io_ins_513 : _GEN_512; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_514 = 10'h202 == io_sel ? io_ins_514 : _GEN_513; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_515 = 10'h203 == io_sel ? io_ins_515 : _GEN_514; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_516 = 10'h204 == io_sel ? io_ins_516 : _GEN_515; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_517 = 10'h205 == io_sel ? io_ins_517 : _GEN_516; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_518 = 10'h206 == io_sel ? io_ins_518 : _GEN_517; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_519 = 10'h207 == io_sel ? io_ins_519 : _GEN_518; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_520 = 10'h208 == io_sel ? io_ins_520 : _GEN_519; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_521 = 10'h209 == io_sel ? io_ins_521 : _GEN_520; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_522 = 10'h20a == io_sel ? io_ins_522 : _GEN_521; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_523 = 10'h20b == io_sel ? io_ins_523 : _GEN_522; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_524 = 10'h20c == io_sel ? io_ins_524 : _GEN_523; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_525 = 10'h20d == io_sel ? io_ins_525 : _GEN_524; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_526 = 10'h20e == io_sel ? io_ins_526 : _GEN_525; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_527 = 10'h20f == io_sel ? io_ins_527 : _GEN_526; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_528 = 10'h210 == io_sel ? io_ins_528 : _GEN_527; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_529 = 10'h211 == io_sel ? io_ins_529 : _GEN_528; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_530 = 10'h212 == io_sel ? io_ins_530 : _GEN_529; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_531 = 10'h213 == io_sel ? io_ins_531 : _GEN_530; // @[MuxN.scala 16:10:@39581.4]
  assign _GEN_532 = 10'h214 == io_sel ? io_ins_532 : _GEN_531; // @[MuxN.scala 16:10:@39581.4]
  assign io_out = 10'h215 == io_sel ? io_ins_533 : _GEN_532; // @[MuxN.scala 16:10:@39581.4]
endmodule
module RegFile( // @[:@39583.2]
  input         clock, // @[:@39584.4]
  input         reset, // @[:@39585.4]
  input  [31:0] io_raddr, // @[:@39586.4]
  input         io_wen, // @[:@39586.4]
  input  [31:0] io_waddr, // @[:@39586.4]
  input  [63:0] io_wdata, // @[:@39586.4]
  output [63:0] io_rdata, // @[:@39586.4]
  input         io_reset, // @[:@39586.4]
  output [63:0] io_argIns_0, // @[:@39586.4]
  output [63:0] io_argIns_1, // @[:@39586.4]
  output [63:0] io_argIns_2, // @[:@39586.4]
  input         io_argOuts_0_valid, // @[:@39586.4]
  input  [63:0] io_argOuts_0_bits, // @[:@39586.4]
  input         io_argOuts_1_valid, // @[:@39586.4]
  input  [63:0] io_argOuts_1_bits, // @[:@39586.4]
  input         io_argOuts_2_valid, // @[:@39586.4]
  input  [63:0] io_argOuts_2_bits, // @[:@39586.4]
  input         io_argOuts_3_valid, // @[:@39586.4]
  input  [63:0] io_argOuts_3_bits, // @[:@39586.4]
  input         io_argOuts_4_valid, // @[:@39586.4]
  input  [63:0] io_argOuts_4_bits, // @[:@39586.4]
  input         io_argOuts_5_valid, // @[:@39586.4]
  input  [63:0] io_argOuts_5_bits, // @[:@39586.4]
  input         io_argOuts_6_valid, // @[:@39586.4]
  input  [63:0] io_argOuts_6_bits, // @[:@39586.4]
  input         io_argOuts_7_valid, // @[:@39586.4]
  input  [63:0] io_argOuts_7_bits, // @[:@39586.4]
  input         io_argOuts_8_valid, // @[:@39586.4]
  input  [63:0] io_argOuts_8_bits, // @[:@39586.4]
  input         io_argOuts_9_valid, // @[:@39586.4]
  input  [63:0] io_argOuts_9_bits, // @[:@39586.4]
  input         io_argOuts_10_valid, // @[:@39586.4]
  input  [63:0] io_argOuts_10_bits, // @[:@39586.4]
  input         io_argOuts_11_valid, // @[:@39586.4]
  input  [63:0] io_argOuts_11_bits, // @[:@39586.4]
  input         io_argOuts_12_valid, // @[:@39586.4]
  input  [63:0] io_argOuts_12_bits, // @[:@39586.4]
  input         io_argOuts_13_valid, // @[:@39586.4]
  input  [63:0] io_argOuts_13_bits, // @[:@39586.4]
  input         io_argOuts_14_valid, // @[:@39586.4]
  input  [63:0] io_argOuts_14_bits, // @[:@39586.4]
  input         io_argOuts_15_valid, // @[:@39586.4]
  input  [63:0] io_argOuts_15_bits, // @[:@39586.4]
  input         io_argOuts_16_valid, // @[:@39586.4]
  input  [63:0] io_argOuts_16_bits, // @[:@39586.4]
  input         io_argOuts_17_valid, // @[:@39586.4]
  input  [63:0] io_argOuts_17_bits, // @[:@39586.4]
  input         io_argOuts_18_valid, // @[:@39586.4]
  input  [63:0] io_argOuts_18_bits, // @[:@39586.4]
  input         io_argOuts_19_valid, // @[:@39586.4]
  input  [63:0] io_argOuts_19_bits, // @[:@39586.4]
  input         io_argOuts_20_valid, // @[:@39586.4]
  input  [63:0] io_argOuts_20_bits, // @[:@39586.4]
  input         io_argOuts_21_valid, // @[:@39586.4]
  input  [63:0] io_argOuts_21_bits, // @[:@39586.4]
  input         io_argOuts_22_valid, // @[:@39586.4]
  input  [63:0] io_argOuts_22_bits, // @[:@39586.4]
  input         io_argOuts_23_valid, // @[:@39586.4]
  input  [63:0] io_argOuts_23_bits, // @[:@39586.4]
  input         io_argOuts_24_valid, // @[:@39586.4]
  input  [63:0] io_argOuts_24_bits, // @[:@39586.4]
  input         io_argOuts_25_valid, // @[:@39586.4]
  input  [63:0] io_argOuts_25_bits, // @[:@39586.4]
  input         io_argOuts_26_valid, // @[:@39586.4]
  input  [63:0] io_argOuts_26_bits, // @[:@39586.4]
  input         io_argOuts_27_valid, // @[:@39586.4]
  input  [63:0] io_argOuts_27_bits, // @[:@39586.4]
  input         io_argOuts_28_valid, // @[:@39586.4]
  input  [63:0] io_argOuts_28_bits, // @[:@39586.4]
  input         io_argOuts_29_valid, // @[:@39586.4]
  input  [63:0] io_argOuts_29_bits, // @[:@39586.4]
  input         io_argOuts_30_valid, // @[:@39586.4]
  input  [63:0] io_argOuts_30_bits, // @[:@39586.4]
  input         io_argOuts_31_valid, // @[:@39586.4]
  input  [63:0] io_argOuts_31_bits, // @[:@39586.4]
  input         io_argOuts_32_valid, // @[:@39586.4]
  input  [63:0] io_argOuts_32_bits // @[:@39586.4]
);
  wire  regs_0_clock; // @[RegFile.scala 66:20:@41720.4]
  wire  regs_0_reset; // @[RegFile.scala 66:20:@41720.4]
  wire [63:0] regs_0_io_in; // @[RegFile.scala 66:20:@41720.4]
  wire  regs_0_io_reset; // @[RegFile.scala 66:20:@41720.4]
  wire [63:0] regs_0_io_out; // @[RegFile.scala 66:20:@41720.4]
  wire  regs_0_io_enable; // @[RegFile.scala 66:20:@41720.4]
  wire  regs_1_clock; // @[RegFile.scala 66:20:@41732.4]
  wire  regs_1_reset; // @[RegFile.scala 66:20:@41732.4]
  wire [63:0] regs_1_io_in; // @[RegFile.scala 66:20:@41732.4]
  wire  regs_1_io_reset; // @[RegFile.scala 66:20:@41732.4]
  wire [63:0] regs_1_io_out; // @[RegFile.scala 66:20:@41732.4]
  wire  regs_1_io_enable; // @[RegFile.scala 66:20:@41732.4]
  wire  regs_2_clock; // @[RegFile.scala 66:20:@41751.4]
  wire  regs_2_reset; // @[RegFile.scala 66:20:@41751.4]
  wire [63:0] regs_2_io_in; // @[RegFile.scala 66:20:@41751.4]
  wire  regs_2_io_reset; // @[RegFile.scala 66:20:@41751.4]
  wire [63:0] regs_2_io_out; // @[RegFile.scala 66:20:@41751.4]
  wire  regs_2_io_enable; // @[RegFile.scala 66:20:@41751.4]
  wire  regs_3_clock; // @[RegFile.scala 66:20:@41763.4]
  wire  regs_3_reset; // @[RegFile.scala 66:20:@41763.4]
  wire [63:0] regs_3_io_in; // @[RegFile.scala 66:20:@41763.4]
  wire  regs_3_io_reset; // @[RegFile.scala 66:20:@41763.4]
  wire [63:0] regs_3_io_out; // @[RegFile.scala 66:20:@41763.4]
  wire  regs_3_io_enable; // @[RegFile.scala 66:20:@41763.4]
  wire  regs_4_clock; // @[RegFile.scala 66:20:@41777.4]
  wire  regs_4_reset; // @[RegFile.scala 66:20:@41777.4]
  wire [63:0] regs_4_io_in; // @[RegFile.scala 66:20:@41777.4]
  wire  regs_4_io_reset; // @[RegFile.scala 66:20:@41777.4]
  wire [63:0] regs_4_io_out; // @[RegFile.scala 66:20:@41777.4]
  wire  regs_4_io_enable; // @[RegFile.scala 66:20:@41777.4]
  wire  regs_5_clock; // @[RegFile.scala 66:20:@41791.4]
  wire  regs_5_reset; // @[RegFile.scala 66:20:@41791.4]
  wire [63:0] regs_5_io_in; // @[RegFile.scala 66:20:@41791.4]
  wire  regs_5_io_reset; // @[RegFile.scala 66:20:@41791.4]
  wire [63:0] regs_5_io_out; // @[RegFile.scala 66:20:@41791.4]
  wire  regs_5_io_enable; // @[RegFile.scala 66:20:@41791.4]
  wire  regs_6_clock; // @[RegFile.scala 66:20:@41805.4]
  wire  regs_6_reset; // @[RegFile.scala 66:20:@41805.4]
  wire [63:0] regs_6_io_in; // @[RegFile.scala 66:20:@41805.4]
  wire  regs_6_io_reset; // @[RegFile.scala 66:20:@41805.4]
  wire [63:0] regs_6_io_out; // @[RegFile.scala 66:20:@41805.4]
  wire  regs_6_io_enable; // @[RegFile.scala 66:20:@41805.4]
  wire  regs_7_clock; // @[RegFile.scala 66:20:@41819.4]
  wire  regs_7_reset; // @[RegFile.scala 66:20:@41819.4]
  wire [63:0] regs_7_io_in; // @[RegFile.scala 66:20:@41819.4]
  wire  regs_7_io_reset; // @[RegFile.scala 66:20:@41819.4]
  wire [63:0] regs_7_io_out; // @[RegFile.scala 66:20:@41819.4]
  wire  regs_7_io_enable; // @[RegFile.scala 66:20:@41819.4]
  wire  regs_8_clock; // @[RegFile.scala 66:20:@41833.4]
  wire  regs_8_reset; // @[RegFile.scala 66:20:@41833.4]
  wire [63:0] regs_8_io_in; // @[RegFile.scala 66:20:@41833.4]
  wire  regs_8_io_reset; // @[RegFile.scala 66:20:@41833.4]
  wire [63:0] regs_8_io_out; // @[RegFile.scala 66:20:@41833.4]
  wire  regs_8_io_enable; // @[RegFile.scala 66:20:@41833.4]
  wire  regs_9_clock; // @[RegFile.scala 66:20:@41847.4]
  wire  regs_9_reset; // @[RegFile.scala 66:20:@41847.4]
  wire [63:0] regs_9_io_in; // @[RegFile.scala 66:20:@41847.4]
  wire  regs_9_io_reset; // @[RegFile.scala 66:20:@41847.4]
  wire [63:0] regs_9_io_out; // @[RegFile.scala 66:20:@41847.4]
  wire  regs_9_io_enable; // @[RegFile.scala 66:20:@41847.4]
  wire  regs_10_clock; // @[RegFile.scala 66:20:@41861.4]
  wire  regs_10_reset; // @[RegFile.scala 66:20:@41861.4]
  wire [63:0] regs_10_io_in; // @[RegFile.scala 66:20:@41861.4]
  wire  regs_10_io_reset; // @[RegFile.scala 66:20:@41861.4]
  wire [63:0] regs_10_io_out; // @[RegFile.scala 66:20:@41861.4]
  wire  regs_10_io_enable; // @[RegFile.scala 66:20:@41861.4]
  wire  regs_11_clock; // @[RegFile.scala 66:20:@41875.4]
  wire  regs_11_reset; // @[RegFile.scala 66:20:@41875.4]
  wire [63:0] regs_11_io_in; // @[RegFile.scala 66:20:@41875.4]
  wire  regs_11_io_reset; // @[RegFile.scala 66:20:@41875.4]
  wire [63:0] regs_11_io_out; // @[RegFile.scala 66:20:@41875.4]
  wire  regs_11_io_enable; // @[RegFile.scala 66:20:@41875.4]
  wire  regs_12_clock; // @[RegFile.scala 66:20:@41889.4]
  wire  regs_12_reset; // @[RegFile.scala 66:20:@41889.4]
  wire [63:0] regs_12_io_in; // @[RegFile.scala 66:20:@41889.4]
  wire  regs_12_io_reset; // @[RegFile.scala 66:20:@41889.4]
  wire [63:0] regs_12_io_out; // @[RegFile.scala 66:20:@41889.4]
  wire  regs_12_io_enable; // @[RegFile.scala 66:20:@41889.4]
  wire  regs_13_clock; // @[RegFile.scala 66:20:@41903.4]
  wire  regs_13_reset; // @[RegFile.scala 66:20:@41903.4]
  wire [63:0] regs_13_io_in; // @[RegFile.scala 66:20:@41903.4]
  wire  regs_13_io_reset; // @[RegFile.scala 66:20:@41903.4]
  wire [63:0] regs_13_io_out; // @[RegFile.scala 66:20:@41903.4]
  wire  regs_13_io_enable; // @[RegFile.scala 66:20:@41903.4]
  wire  regs_14_clock; // @[RegFile.scala 66:20:@41917.4]
  wire  regs_14_reset; // @[RegFile.scala 66:20:@41917.4]
  wire [63:0] regs_14_io_in; // @[RegFile.scala 66:20:@41917.4]
  wire  regs_14_io_reset; // @[RegFile.scala 66:20:@41917.4]
  wire [63:0] regs_14_io_out; // @[RegFile.scala 66:20:@41917.4]
  wire  regs_14_io_enable; // @[RegFile.scala 66:20:@41917.4]
  wire  regs_15_clock; // @[RegFile.scala 66:20:@41931.4]
  wire  regs_15_reset; // @[RegFile.scala 66:20:@41931.4]
  wire [63:0] regs_15_io_in; // @[RegFile.scala 66:20:@41931.4]
  wire  regs_15_io_reset; // @[RegFile.scala 66:20:@41931.4]
  wire [63:0] regs_15_io_out; // @[RegFile.scala 66:20:@41931.4]
  wire  regs_15_io_enable; // @[RegFile.scala 66:20:@41931.4]
  wire  regs_16_clock; // @[RegFile.scala 66:20:@41945.4]
  wire  regs_16_reset; // @[RegFile.scala 66:20:@41945.4]
  wire [63:0] regs_16_io_in; // @[RegFile.scala 66:20:@41945.4]
  wire  regs_16_io_reset; // @[RegFile.scala 66:20:@41945.4]
  wire [63:0] regs_16_io_out; // @[RegFile.scala 66:20:@41945.4]
  wire  regs_16_io_enable; // @[RegFile.scala 66:20:@41945.4]
  wire  regs_17_clock; // @[RegFile.scala 66:20:@41959.4]
  wire  regs_17_reset; // @[RegFile.scala 66:20:@41959.4]
  wire [63:0] regs_17_io_in; // @[RegFile.scala 66:20:@41959.4]
  wire  regs_17_io_reset; // @[RegFile.scala 66:20:@41959.4]
  wire [63:0] regs_17_io_out; // @[RegFile.scala 66:20:@41959.4]
  wire  regs_17_io_enable; // @[RegFile.scala 66:20:@41959.4]
  wire  regs_18_clock; // @[RegFile.scala 66:20:@41973.4]
  wire  regs_18_reset; // @[RegFile.scala 66:20:@41973.4]
  wire [63:0] regs_18_io_in; // @[RegFile.scala 66:20:@41973.4]
  wire  regs_18_io_reset; // @[RegFile.scala 66:20:@41973.4]
  wire [63:0] regs_18_io_out; // @[RegFile.scala 66:20:@41973.4]
  wire  regs_18_io_enable; // @[RegFile.scala 66:20:@41973.4]
  wire  regs_19_clock; // @[RegFile.scala 66:20:@41987.4]
  wire  regs_19_reset; // @[RegFile.scala 66:20:@41987.4]
  wire [63:0] regs_19_io_in; // @[RegFile.scala 66:20:@41987.4]
  wire  regs_19_io_reset; // @[RegFile.scala 66:20:@41987.4]
  wire [63:0] regs_19_io_out; // @[RegFile.scala 66:20:@41987.4]
  wire  regs_19_io_enable; // @[RegFile.scala 66:20:@41987.4]
  wire  regs_20_clock; // @[RegFile.scala 66:20:@42001.4]
  wire  regs_20_reset; // @[RegFile.scala 66:20:@42001.4]
  wire [63:0] regs_20_io_in; // @[RegFile.scala 66:20:@42001.4]
  wire  regs_20_io_reset; // @[RegFile.scala 66:20:@42001.4]
  wire [63:0] regs_20_io_out; // @[RegFile.scala 66:20:@42001.4]
  wire  regs_20_io_enable; // @[RegFile.scala 66:20:@42001.4]
  wire  regs_21_clock; // @[RegFile.scala 66:20:@42015.4]
  wire  regs_21_reset; // @[RegFile.scala 66:20:@42015.4]
  wire [63:0] regs_21_io_in; // @[RegFile.scala 66:20:@42015.4]
  wire  regs_21_io_reset; // @[RegFile.scala 66:20:@42015.4]
  wire [63:0] regs_21_io_out; // @[RegFile.scala 66:20:@42015.4]
  wire  regs_21_io_enable; // @[RegFile.scala 66:20:@42015.4]
  wire  regs_22_clock; // @[RegFile.scala 66:20:@42029.4]
  wire  regs_22_reset; // @[RegFile.scala 66:20:@42029.4]
  wire [63:0] regs_22_io_in; // @[RegFile.scala 66:20:@42029.4]
  wire  regs_22_io_reset; // @[RegFile.scala 66:20:@42029.4]
  wire [63:0] regs_22_io_out; // @[RegFile.scala 66:20:@42029.4]
  wire  regs_22_io_enable; // @[RegFile.scala 66:20:@42029.4]
  wire  regs_23_clock; // @[RegFile.scala 66:20:@42043.4]
  wire  regs_23_reset; // @[RegFile.scala 66:20:@42043.4]
  wire [63:0] regs_23_io_in; // @[RegFile.scala 66:20:@42043.4]
  wire  regs_23_io_reset; // @[RegFile.scala 66:20:@42043.4]
  wire [63:0] regs_23_io_out; // @[RegFile.scala 66:20:@42043.4]
  wire  regs_23_io_enable; // @[RegFile.scala 66:20:@42043.4]
  wire  regs_24_clock; // @[RegFile.scala 66:20:@42057.4]
  wire  regs_24_reset; // @[RegFile.scala 66:20:@42057.4]
  wire [63:0] regs_24_io_in; // @[RegFile.scala 66:20:@42057.4]
  wire  regs_24_io_reset; // @[RegFile.scala 66:20:@42057.4]
  wire [63:0] regs_24_io_out; // @[RegFile.scala 66:20:@42057.4]
  wire  regs_24_io_enable; // @[RegFile.scala 66:20:@42057.4]
  wire  regs_25_clock; // @[RegFile.scala 66:20:@42071.4]
  wire  regs_25_reset; // @[RegFile.scala 66:20:@42071.4]
  wire [63:0] regs_25_io_in; // @[RegFile.scala 66:20:@42071.4]
  wire  regs_25_io_reset; // @[RegFile.scala 66:20:@42071.4]
  wire [63:0] regs_25_io_out; // @[RegFile.scala 66:20:@42071.4]
  wire  regs_25_io_enable; // @[RegFile.scala 66:20:@42071.4]
  wire  regs_26_clock; // @[RegFile.scala 66:20:@42085.4]
  wire  regs_26_reset; // @[RegFile.scala 66:20:@42085.4]
  wire [63:0] regs_26_io_in; // @[RegFile.scala 66:20:@42085.4]
  wire  regs_26_io_reset; // @[RegFile.scala 66:20:@42085.4]
  wire [63:0] regs_26_io_out; // @[RegFile.scala 66:20:@42085.4]
  wire  regs_26_io_enable; // @[RegFile.scala 66:20:@42085.4]
  wire  regs_27_clock; // @[RegFile.scala 66:20:@42099.4]
  wire  regs_27_reset; // @[RegFile.scala 66:20:@42099.4]
  wire [63:0] regs_27_io_in; // @[RegFile.scala 66:20:@42099.4]
  wire  regs_27_io_reset; // @[RegFile.scala 66:20:@42099.4]
  wire [63:0] regs_27_io_out; // @[RegFile.scala 66:20:@42099.4]
  wire  regs_27_io_enable; // @[RegFile.scala 66:20:@42099.4]
  wire  regs_28_clock; // @[RegFile.scala 66:20:@42113.4]
  wire  regs_28_reset; // @[RegFile.scala 66:20:@42113.4]
  wire [63:0] regs_28_io_in; // @[RegFile.scala 66:20:@42113.4]
  wire  regs_28_io_reset; // @[RegFile.scala 66:20:@42113.4]
  wire [63:0] regs_28_io_out; // @[RegFile.scala 66:20:@42113.4]
  wire  regs_28_io_enable; // @[RegFile.scala 66:20:@42113.4]
  wire  regs_29_clock; // @[RegFile.scala 66:20:@42127.4]
  wire  regs_29_reset; // @[RegFile.scala 66:20:@42127.4]
  wire [63:0] regs_29_io_in; // @[RegFile.scala 66:20:@42127.4]
  wire  regs_29_io_reset; // @[RegFile.scala 66:20:@42127.4]
  wire [63:0] regs_29_io_out; // @[RegFile.scala 66:20:@42127.4]
  wire  regs_29_io_enable; // @[RegFile.scala 66:20:@42127.4]
  wire  regs_30_clock; // @[RegFile.scala 66:20:@42141.4]
  wire  regs_30_reset; // @[RegFile.scala 66:20:@42141.4]
  wire [63:0] regs_30_io_in; // @[RegFile.scala 66:20:@42141.4]
  wire  regs_30_io_reset; // @[RegFile.scala 66:20:@42141.4]
  wire [63:0] regs_30_io_out; // @[RegFile.scala 66:20:@42141.4]
  wire  regs_30_io_enable; // @[RegFile.scala 66:20:@42141.4]
  wire  regs_31_clock; // @[RegFile.scala 66:20:@42155.4]
  wire  regs_31_reset; // @[RegFile.scala 66:20:@42155.4]
  wire [63:0] regs_31_io_in; // @[RegFile.scala 66:20:@42155.4]
  wire  regs_31_io_reset; // @[RegFile.scala 66:20:@42155.4]
  wire [63:0] regs_31_io_out; // @[RegFile.scala 66:20:@42155.4]
  wire  regs_31_io_enable; // @[RegFile.scala 66:20:@42155.4]
  wire  regs_32_clock; // @[RegFile.scala 66:20:@42169.4]
  wire  regs_32_reset; // @[RegFile.scala 66:20:@42169.4]
  wire [63:0] regs_32_io_in; // @[RegFile.scala 66:20:@42169.4]
  wire  regs_32_io_reset; // @[RegFile.scala 66:20:@42169.4]
  wire [63:0] regs_32_io_out; // @[RegFile.scala 66:20:@42169.4]
  wire  regs_32_io_enable; // @[RegFile.scala 66:20:@42169.4]
  wire  regs_33_clock; // @[RegFile.scala 66:20:@42183.4]
  wire  regs_33_reset; // @[RegFile.scala 66:20:@42183.4]
  wire [63:0] regs_33_io_in; // @[RegFile.scala 66:20:@42183.4]
  wire  regs_33_io_reset; // @[RegFile.scala 66:20:@42183.4]
  wire [63:0] regs_33_io_out; // @[RegFile.scala 66:20:@42183.4]
  wire  regs_33_io_enable; // @[RegFile.scala 66:20:@42183.4]
  wire  regs_34_clock; // @[RegFile.scala 66:20:@42197.4]
  wire  regs_34_reset; // @[RegFile.scala 66:20:@42197.4]
  wire [63:0] regs_34_io_in; // @[RegFile.scala 66:20:@42197.4]
  wire  regs_34_io_reset; // @[RegFile.scala 66:20:@42197.4]
  wire [63:0] regs_34_io_out; // @[RegFile.scala 66:20:@42197.4]
  wire  regs_34_io_enable; // @[RegFile.scala 66:20:@42197.4]
  wire  regs_35_clock; // @[RegFile.scala 66:20:@42211.4]
  wire  regs_35_reset; // @[RegFile.scala 66:20:@42211.4]
  wire [63:0] regs_35_io_in; // @[RegFile.scala 66:20:@42211.4]
  wire  regs_35_io_reset; // @[RegFile.scala 66:20:@42211.4]
  wire [63:0] regs_35_io_out; // @[RegFile.scala 66:20:@42211.4]
  wire  regs_35_io_enable; // @[RegFile.scala 66:20:@42211.4]
  wire  regs_36_clock; // @[RegFile.scala 66:20:@42225.4]
  wire  regs_36_reset; // @[RegFile.scala 66:20:@42225.4]
  wire [63:0] regs_36_io_in; // @[RegFile.scala 66:20:@42225.4]
  wire  regs_36_io_reset; // @[RegFile.scala 66:20:@42225.4]
  wire [63:0] regs_36_io_out; // @[RegFile.scala 66:20:@42225.4]
  wire  regs_36_io_enable; // @[RegFile.scala 66:20:@42225.4]
  wire  regs_37_clock; // @[RegFile.scala 66:20:@42239.4]
  wire  regs_37_reset; // @[RegFile.scala 66:20:@42239.4]
  wire [63:0] regs_37_io_in; // @[RegFile.scala 66:20:@42239.4]
  wire  regs_37_io_reset; // @[RegFile.scala 66:20:@42239.4]
  wire [63:0] regs_37_io_out; // @[RegFile.scala 66:20:@42239.4]
  wire  regs_37_io_enable; // @[RegFile.scala 66:20:@42239.4]
  wire  regs_38_clock; // @[RegFile.scala 66:20:@42253.4]
  wire  regs_38_reset; // @[RegFile.scala 66:20:@42253.4]
  wire [63:0] regs_38_io_in; // @[RegFile.scala 66:20:@42253.4]
  wire  regs_38_io_reset; // @[RegFile.scala 66:20:@42253.4]
  wire [63:0] regs_38_io_out; // @[RegFile.scala 66:20:@42253.4]
  wire  regs_38_io_enable; // @[RegFile.scala 66:20:@42253.4]
  wire  regs_39_clock; // @[RegFile.scala 66:20:@42267.4]
  wire  regs_39_reset; // @[RegFile.scala 66:20:@42267.4]
  wire [63:0] regs_39_io_in; // @[RegFile.scala 66:20:@42267.4]
  wire  regs_39_io_reset; // @[RegFile.scala 66:20:@42267.4]
  wire [63:0] regs_39_io_out; // @[RegFile.scala 66:20:@42267.4]
  wire  regs_39_io_enable; // @[RegFile.scala 66:20:@42267.4]
  wire  regs_40_clock; // @[RegFile.scala 66:20:@42281.4]
  wire  regs_40_reset; // @[RegFile.scala 66:20:@42281.4]
  wire [63:0] regs_40_io_in; // @[RegFile.scala 66:20:@42281.4]
  wire  regs_40_io_reset; // @[RegFile.scala 66:20:@42281.4]
  wire [63:0] regs_40_io_out; // @[RegFile.scala 66:20:@42281.4]
  wire  regs_40_io_enable; // @[RegFile.scala 66:20:@42281.4]
  wire  regs_41_clock; // @[RegFile.scala 66:20:@42295.4]
  wire  regs_41_reset; // @[RegFile.scala 66:20:@42295.4]
  wire [63:0] regs_41_io_in; // @[RegFile.scala 66:20:@42295.4]
  wire  regs_41_io_reset; // @[RegFile.scala 66:20:@42295.4]
  wire [63:0] regs_41_io_out; // @[RegFile.scala 66:20:@42295.4]
  wire  regs_41_io_enable; // @[RegFile.scala 66:20:@42295.4]
  wire  regs_42_clock; // @[RegFile.scala 66:20:@42309.4]
  wire  regs_42_reset; // @[RegFile.scala 66:20:@42309.4]
  wire [63:0] regs_42_io_in; // @[RegFile.scala 66:20:@42309.4]
  wire  regs_42_io_reset; // @[RegFile.scala 66:20:@42309.4]
  wire [63:0] regs_42_io_out; // @[RegFile.scala 66:20:@42309.4]
  wire  regs_42_io_enable; // @[RegFile.scala 66:20:@42309.4]
  wire  regs_43_clock; // @[RegFile.scala 66:20:@42323.4]
  wire  regs_43_reset; // @[RegFile.scala 66:20:@42323.4]
  wire [63:0] regs_43_io_in; // @[RegFile.scala 66:20:@42323.4]
  wire  regs_43_io_reset; // @[RegFile.scala 66:20:@42323.4]
  wire [63:0] regs_43_io_out; // @[RegFile.scala 66:20:@42323.4]
  wire  regs_43_io_enable; // @[RegFile.scala 66:20:@42323.4]
  wire  regs_44_clock; // @[RegFile.scala 66:20:@42337.4]
  wire  regs_44_reset; // @[RegFile.scala 66:20:@42337.4]
  wire [63:0] regs_44_io_in; // @[RegFile.scala 66:20:@42337.4]
  wire  regs_44_io_reset; // @[RegFile.scala 66:20:@42337.4]
  wire [63:0] regs_44_io_out; // @[RegFile.scala 66:20:@42337.4]
  wire  regs_44_io_enable; // @[RegFile.scala 66:20:@42337.4]
  wire  regs_45_clock; // @[RegFile.scala 66:20:@42351.4]
  wire  regs_45_reset; // @[RegFile.scala 66:20:@42351.4]
  wire [63:0] regs_45_io_in; // @[RegFile.scala 66:20:@42351.4]
  wire  regs_45_io_reset; // @[RegFile.scala 66:20:@42351.4]
  wire [63:0] regs_45_io_out; // @[RegFile.scala 66:20:@42351.4]
  wire  regs_45_io_enable; // @[RegFile.scala 66:20:@42351.4]
  wire  regs_46_clock; // @[RegFile.scala 66:20:@42365.4]
  wire  regs_46_reset; // @[RegFile.scala 66:20:@42365.4]
  wire [63:0] regs_46_io_in; // @[RegFile.scala 66:20:@42365.4]
  wire  regs_46_io_reset; // @[RegFile.scala 66:20:@42365.4]
  wire [63:0] regs_46_io_out; // @[RegFile.scala 66:20:@42365.4]
  wire  regs_46_io_enable; // @[RegFile.scala 66:20:@42365.4]
  wire  regs_47_clock; // @[RegFile.scala 66:20:@42379.4]
  wire  regs_47_reset; // @[RegFile.scala 66:20:@42379.4]
  wire [63:0] regs_47_io_in; // @[RegFile.scala 66:20:@42379.4]
  wire  regs_47_io_reset; // @[RegFile.scala 66:20:@42379.4]
  wire [63:0] regs_47_io_out; // @[RegFile.scala 66:20:@42379.4]
  wire  regs_47_io_enable; // @[RegFile.scala 66:20:@42379.4]
  wire  regs_48_clock; // @[RegFile.scala 66:20:@42393.4]
  wire  regs_48_reset; // @[RegFile.scala 66:20:@42393.4]
  wire [63:0] regs_48_io_in; // @[RegFile.scala 66:20:@42393.4]
  wire  regs_48_io_reset; // @[RegFile.scala 66:20:@42393.4]
  wire [63:0] regs_48_io_out; // @[RegFile.scala 66:20:@42393.4]
  wire  regs_48_io_enable; // @[RegFile.scala 66:20:@42393.4]
  wire  regs_49_clock; // @[RegFile.scala 66:20:@42407.4]
  wire  regs_49_reset; // @[RegFile.scala 66:20:@42407.4]
  wire [63:0] regs_49_io_in; // @[RegFile.scala 66:20:@42407.4]
  wire  regs_49_io_reset; // @[RegFile.scala 66:20:@42407.4]
  wire [63:0] regs_49_io_out; // @[RegFile.scala 66:20:@42407.4]
  wire  regs_49_io_enable; // @[RegFile.scala 66:20:@42407.4]
  wire  regs_50_clock; // @[RegFile.scala 66:20:@42421.4]
  wire  regs_50_reset; // @[RegFile.scala 66:20:@42421.4]
  wire [63:0] regs_50_io_in; // @[RegFile.scala 66:20:@42421.4]
  wire  regs_50_io_reset; // @[RegFile.scala 66:20:@42421.4]
  wire [63:0] regs_50_io_out; // @[RegFile.scala 66:20:@42421.4]
  wire  regs_50_io_enable; // @[RegFile.scala 66:20:@42421.4]
  wire  regs_51_clock; // @[RegFile.scala 66:20:@42435.4]
  wire  regs_51_reset; // @[RegFile.scala 66:20:@42435.4]
  wire [63:0] regs_51_io_in; // @[RegFile.scala 66:20:@42435.4]
  wire  regs_51_io_reset; // @[RegFile.scala 66:20:@42435.4]
  wire [63:0] regs_51_io_out; // @[RegFile.scala 66:20:@42435.4]
  wire  regs_51_io_enable; // @[RegFile.scala 66:20:@42435.4]
  wire  regs_52_clock; // @[RegFile.scala 66:20:@42449.4]
  wire  regs_52_reset; // @[RegFile.scala 66:20:@42449.4]
  wire [63:0] regs_52_io_in; // @[RegFile.scala 66:20:@42449.4]
  wire  regs_52_io_reset; // @[RegFile.scala 66:20:@42449.4]
  wire [63:0] regs_52_io_out; // @[RegFile.scala 66:20:@42449.4]
  wire  regs_52_io_enable; // @[RegFile.scala 66:20:@42449.4]
  wire  regs_53_clock; // @[RegFile.scala 66:20:@42463.4]
  wire  regs_53_reset; // @[RegFile.scala 66:20:@42463.4]
  wire [63:0] regs_53_io_in; // @[RegFile.scala 66:20:@42463.4]
  wire  regs_53_io_reset; // @[RegFile.scala 66:20:@42463.4]
  wire [63:0] regs_53_io_out; // @[RegFile.scala 66:20:@42463.4]
  wire  regs_53_io_enable; // @[RegFile.scala 66:20:@42463.4]
  wire  regs_54_clock; // @[RegFile.scala 66:20:@42477.4]
  wire  regs_54_reset; // @[RegFile.scala 66:20:@42477.4]
  wire [63:0] regs_54_io_in; // @[RegFile.scala 66:20:@42477.4]
  wire  regs_54_io_reset; // @[RegFile.scala 66:20:@42477.4]
  wire [63:0] regs_54_io_out; // @[RegFile.scala 66:20:@42477.4]
  wire  regs_54_io_enable; // @[RegFile.scala 66:20:@42477.4]
  wire  regs_55_clock; // @[RegFile.scala 66:20:@42491.4]
  wire  regs_55_reset; // @[RegFile.scala 66:20:@42491.4]
  wire [63:0] regs_55_io_in; // @[RegFile.scala 66:20:@42491.4]
  wire  regs_55_io_reset; // @[RegFile.scala 66:20:@42491.4]
  wire [63:0] regs_55_io_out; // @[RegFile.scala 66:20:@42491.4]
  wire  regs_55_io_enable; // @[RegFile.scala 66:20:@42491.4]
  wire  regs_56_clock; // @[RegFile.scala 66:20:@42505.4]
  wire  regs_56_reset; // @[RegFile.scala 66:20:@42505.4]
  wire [63:0] regs_56_io_in; // @[RegFile.scala 66:20:@42505.4]
  wire  regs_56_io_reset; // @[RegFile.scala 66:20:@42505.4]
  wire [63:0] regs_56_io_out; // @[RegFile.scala 66:20:@42505.4]
  wire  regs_56_io_enable; // @[RegFile.scala 66:20:@42505.4]
  wire  regs_57_clock; // @[RegFile.scala 66:20:@42519.4]
  wire  regs_57_reset; // @[RegFile.scala 66:20:@42519.4]
  wire [63:0] regs_57_io_in; // @[RegFile.scala 66:20:@42519.4]
  wire  regs_57_io_reset; // @[RegFile.scala 66:20:@42519.4]
  wire [63:0] regs_57_io_out; // @[RegFile.scala 66:20:@42519.4]
  wire  regs_57_io_enable; // @[RegFile.scala 66:20:@42519.4]
  wire  regs_58_clock; // @[RegFile.scala 66:20:@42533.4]
  wire  regs_58_reset; // @[RegFile.scala 66:20:@42533.4]
  wire [63:0] regs_58_io_in; // @[RegFile.scala 66:20:@42533.4]
  wire  regs_58_io_reset; // @[RegFile.scala 66:20:@42533.4]
  wire [63:0] regs_58_io_out; // @[RegFile.scala 66:20:@42533.4]
  wire  regs_58_io_enable; // @[RegFile.scala 66:20:@42533.4]
  wire  regs_59_clock; // @[RegFile.scala 66:20:@42547.4]
  wire  regs_59_reset; // @[RegFile.scala 66:20:@42547.4]
  wire [63:0] regs_59_io_in; // @[RegFile.scala 66:20:@42547.4]
  wire  regs_59_io_reset; // @[RegFile.scala 66:20:@42547.4]
  wire [63:0] regs_59_io_out; // @[RegFile.scala 66:20:@42547.4]
  wire  regs_59_io_enable; // @[RegFile.scala 66:20:@42547.4]
  wire  regs_60_clock; // @[RegFile.scala 66:20:@42561.4]
  wire  regs_60_reset; // @[RegFile.scala 66:20:@42561.4]
  wire [63:0] regs_60_io_in; // @[RegFile.scala 66:20:@42561.4]
  wire  regs_60_io_reset; // @[RegFile.scala 66:20:@42561.4]
  wire [63:0] regs_60_io_out; // @[RegFile.scala 66:20:@42561.4]
  wire  regs_60_io_enable; // @[RegFile.scala 66:20:@42561.4]
  wire  regs_61_clock; // @[RegFile.scala 66:20:@42575.4]
  wire  regs_61_reset; // @[RegFile.scala 66:20:@42575.4]
  wire [63:0] regs_61_io_in; // @[RegFile.scala 66:20:@42575.4]
  wire  regs_61_io_reset; // @[RegFile.scala 66:20:@42575.4]
  wire [63:0] regs_61_io_out; // @[RegFile.scala 66:20:@42575.4]
  wire  regs_61_io_enable; // @[RegFile.scala 66:20:@42575.4]
  wire  regs_62_clock; // @[RegFile.scala 66:20:@42589.4]
  wire  regs_62_reset; // @[RegFile.scala 66:20:@42589.4]
  wire [63:0] regs_62_io_in; // @[RegFile.scala 66:20:@42589.4]
  wire  regs_62_io_reset; // @[RegFile.scala 66:20:@42589.4]
  wire [63:0] regs_62_io_out; // @[RegFile.scala 66:20:@42589.4]
  wire  regs_62_io_enable; // @[RegFile.scala 66:20:@42589.4]
  wire  regs_63_clock; // @[RegFile.scala 66:20:@42603.4]
  wire  regs_63_reset; // @[RegFile.scala 66:20:@42603.4]
  wire [63:0] regs_63_io_in; // @[RegFile.scala 66:20:@42603.4]
  wire  regs_63_io_reset; // @[RegFile.scala 66:20:@42603.4]
  wire [63:0] regs_63_io_out; // @[RegFile.scala 66:20:@42603.4]
  wire  regs_63_io_enable; // @[RegFile.scala 66:20:@42603.4]
  wire  regs_64_clock; // @[RegFile.scala 66:20:@42617.4]
  wire  regs_64_reset; // @[RegFile.scala 66:20:@42617.4]
  wire [63:0] regs_64_io_in; // @[RegFile.scala 66:20:@42617.4]
  wire  regs_64_io_reset; // @[RegFile.scala 66:20:@42617.4]
  wire [63:0] regs_64_io_out; // @[RegFile.scala 66:20:@42617.4]
  wire  regs_64_io_enable; // @[RegFile.scala 66:20:@42617.4]
  wire  regs_65_clock; // @[RegFile.scala 66:20:@42631.4]
  wire  regs_65_reset; // @[RegFile.scala 66:20:@42631.4]
  wire [63:0] regs_65_io_in; // @[RegFile.scala 66:20:@42631.4]
  wire  regs_65_io_reset; // @[RegFile.scala 66:20:@42631.4]
  wire [63:0] regs_65_io_out; // @[RegFile.scala 66:20:@42631.4]
  wire  regs_65_io_enable; // @[RegFile.scala 66:20:@42631.4]
  wire  regs_66_clock; // @[RegFile.scala 66:20:@42645.4]
  wire  regs_66_reset; // @[RegFile.scala 66:20:@42645.4]
  wire [63:0] regs_66_io_in; // @[RegFile.scala 66:20:@42645.4]
  wire  regs_66_io_reset; // @[RegFile.scala 66:20:@42645.4]
  wire [63:0] regs_66_io_out; // @[RegFile.scala 66:20:@42645.4]
  wire  regs_66_io_enable; // @[RegFile.scala 66:20:@42645.4]
  wire  regs_67_clock; // @[RegFile.scala 66:20:@42659.4]
  wire  regs_67_reset; // @[RegFile.scala 66:20:@42659.4]
  wire [63:0] regs_67_io_in; // @[RegFile.scala 66:20:@42659.4]
  wire  regs_67_io_reset; // @[RegFile.scala 66:20:@42659.4]
  wire [63:0] regs_67_io_out; // @[RegFile.scala 66:20:@42659.4]
  wire  regs_67_io_enable; // @[RegFile.scala 66:20:@42659.4]
  wire  regs_68_clock; // @[RegFile.scala 66:20:@42673.4]
  wire  regs_68_reset; // @[RegFile.scala 66:20:@42673.4]
  wire [63:0] regs_68_io_in; // @[RegFile.scala 66:20:@42673.4]
  wire  regs_68_io_reset; // @[RegFile.scala 66:20:@42673.4]
  wire [63:0] regs_68_io_out; // @[RegFile.scala 66:20:@42673.4]
  wire  regs_68_io_enable; // @[RegFile.scala 66:20:@42673.4]
  wire  regs_69_clock; // @[RegFile.scala 66:20:@42687.4]
  wire  regs_69_reset; // @[RegFile.scala 66:20:@42687.4]
  wire [63:0] regs_69_io_in; // @[RegFile.scala 66:20:@42687.4]
  wire  regs_69_io_reset; // @[RegFile.scala 66:20:@42687.4]
  wire [63:0] regs_69_io_out; // @[RegFile.scala 66:20:@42687.4]
  wire  regs_69_io_enable; // @[RegFile.scala 66:20:@42687.4]
  wire  regs_70_clock; // @[RegFile.scala 66:20:@42701.4]
  wire  regs_70_reset; // @[RegFile.scala 66:20:@42701.4]
  wire [63:0] regs_70_io_in; // @[RegFile.scala 66:20:@42701.4]
  wire  regs_70_io_reset; // @[RegFile.scala 66:20:@42701.4]
  wire [63:0] regs_70_io_out; // @[RegFile.scala 66:20:@42701.4]
  wire  regs_70_io_enable; // @[RegFile.scala 66:20:@42701.4]
  wire  regs_71_clock; // @[RegFile.scala 66:20:@42715.4]
  wire  regs_71_reset; // @[RegFile.scala 66:20:@42715.4]
  wire [63:0] regs_71_io_in; // @[RegFile.scala 66:20:@42715.4]
  wire  regs_71_io_reset; // @[RegFile.scala 66:20:@42715.4]
  wire [63:0] regs_71_io_out; // @[RegFile.scala 66:20:@42715.4]
  wire  regs_71_io_enable; // @[RegFile.scala 66:20:@42715.4]
  wire  regs_72_clock; // @[RegFile.scala 66:20:@42729.4]
  wire  regs_72_reset; // @[RegFile.scala 66:20:@42729.4]
  wire [63:0] regs_72_io_in; // @[RegFile.scala 66:20:@42729.4]
  wire  regs_72_io_reset; // @[RegFile.scala 66:20:@42729.4]
  wire [63:0] regs_72_io_out; // @[RegFile.scala 66:20:@42729.4]
  wire  regs_72_io_enable; // @[RegFile.scala 66:20:@42729.4]
  wire  regs_73_clock; // @[RegFile.scala 66:20:@42743.4]
  wire  regs_73_reset; // @[RegFile.scala 66:20:@42743.4]
  wire [63:0] regs_73_io_in; // @[RegFile.scala 66:20:@42743.4]
  wire  regs_73_io_reset; // @[RegFile.scala 66:20:@42743.4]
  wire [63:0] regs_73_io_out; // @[RegFile.scala 66:20:@42743.4]
  wire  regs_73_io_enable; // @[RegFile.scala 66:20:@42743.4]
  wire  regs_74_clock; // @[RegFile.scala 66:20:@42757.4]
  wire  regs_74_reset; // @[RegFile.scala 66:20:@42757.4]
  wire [63:0] regs_74_io_in; // @[RegFile.scala 66:20:@42757.4]
  wire  regs_74_io_reset; // @[RegFile.scala 66:20:@42757.4]
  wire [63:0] regs_74_io_out; // @[RegFile.scala 66:20:@42757.4]
  wire  regs_74_io_enable; // @[RegFile.scala 66:20:@42757.4]
  wire  regs_75_clock; // @[RegFile.scala 66:20:@42771.4]
  wire  regs_75_reset; // @[RegFile.scala 66:20:@42771.4]
  wire [63:0] regs_75_io_in; // @[RegFile.scala 66:20:@42771.4]
  wire  regs_75_io_reset; // @[RegFile.scala 66:20:@42771.4]
  wire [63:0] regs_75_io_out; // @[RegFile.scala 66:20:@42771.4]
  wire  regs_75_io_enable; // @[RegFile.scala 66:20:@42771.4]
  wire  regs_76_clock; // @[RegFile.scala 66:20:@42785.4]
  wire  regs_76_reset; // @[RegFile.scala 66:20:@42785.4]
  wire [63:0] regs_76_io_in; // @[RegFile.scala 66:20:@42785.4]
  wire  regs_76_io_reset; // @[RegFile.scala 66:20:@42785.4]
  wire [63:0] regs_76_io_out; // @[RegFile.scala 66:20:@42785.4]
  wire  regs_76_io_enable; // @[RegFile.scala 66:20:@42785.4]
  wire  regs_77_clock; // @[RegFile.scala 66:20:@42799.4]
  wire  regs_77_reset; // @[RegFile.scala 66:20:@42799.4]
  wire [63:0] regs_77_io_in; // @[RegFile.scala 66:20:@42799.4]
  wire  regs_77_io_reset; // @[RegFile.scala 66:20:@42799.4]
  wire [63:0] regs_77_io_out; // @[RegFile.scala 66:20:@42799.4]
  wire  regs_77_io_enable; // @[RegFile.scala 66:20:@42799.4]
  wire  regs_78_clock; // @[RegFile.scala 66:20:@42813.4]
  wire  regs_78_reset; // @[RegFile.scala 66:20:@42813.4]
  wire [63:0] regs_78_io_in; // @[RegFile.scala 66:20:@42813.4]
  wire  regs_78_io_reset; // @[RegFile.scala 66:20:@42813.4]
  wire [63:0] regs_78_io_out; // @[RegFile.scala 66:20:@42813.4]
  wire  regs_78_io_enable; // @[RegFile.scala 66:20:@42813.4]
  wire  regs_79_clock; // @[RegFile.scala 66:20:@42827.4]
  wire  regs_79_reset; // @[RegFile.scala 66:20:@42827.4]
  wire [63:0] regs_79_io_in; // @[RegFile.scala 66:20:@42827.4]
  wire  regs_79_io_reset; // @[RegFile.scala 66:20:@42827.4]
  wire [63:0] regs_79_io_out; // @[RegFile.scala 66:20:@42827.4]
  wire  regs_79_io_enable; // @[RegFile.scala 66:20:@42827.4]
  wire  regs_80_clock; // @[RegFile.scala 66:20:@42841.4]
  wire  regs_80_reset; // @[RegFile.scala 66:20:@42841.4]
  wire [63:0] regs_80_io_in; // @[RegFile.scala 66:20:@42841.4]
  wire  regs_80_io_reset; // @[RegFile.scala 66:20:@42841.4]
  wire [63:0] regs_80_io_out; // @[RegFile.scala 66:20:@42841.4]
  wire  regs_80_io_enable; // @[RegFile.scala 66:20:@42841.4]
  wire  regs_81_clock; // @[RegFile.scala 66:20:@42855.4]
  wire  regs_81_reset; // @[RegFile.scala 66:20:@42855.4]
  wire [63:0] regs_81_io_in; // @[RegFile.scala 66:20:@42855.4]
  wire  regs_81_io_reset; // @[RegFile.scala 66:20:@42855.4]
  wire [63:0] regs_81_io_out; // @[RegFile.scala 66:20:@42855.4]
  wire  regs_81_io_enable; // @[RegFile.scala 66:20:@42855.4]
  wire  regs_82_clock; // @[RegFile.scala 66:20:@42869.4]
  wire  regs_82_reset; // @[RegFile.scala 66:20:@42869.4]
  wire [63:0] regs_82_io_in; // @[RegFile.scala 66:20:@42869.4]
  wire  regs_82_io_reset; // @[RegFile.scala 66:20:@42869.4]
  wire [63:0] regs_82_io_out; // @[RegFile.scala 66:20:@42869.4]
  wire  regs_82_io_enable; // @[RegFile.scala 66:20:@42869.4]
  wire  regs_83_clock; // @[RegFile.scala 66:20:@42883.4]
  wire  regs_83_reset; // @[RegFile.scala 66:20:@42883.4]
  wire [63:0] regs_83_io_in; // @[RegFile.scala 66:20:@42883.4]
  wire  regs_83_io_reset; // @[RegFile.scala 66:20:@42883.4]
  wire [63:0] regs_83_io_out; // @[RegFile.scala 66:20:@42883.4]
  wire  regs_83_io_enable; // @[RegFile.scala 66:20:@42883.4]
  wire  regs_84_clock; // @[RegFile.scala 66:20:@42897.4]
  wire  regs_84_reset; // @[RegFile.scala 66:20:@42897.4]
  wire [63:0] regs_84_io_in; // @[RegFile.scala 66:20:@42897.4]
  wire  regs_84_io_reset; // @[RegFile.scala 66:20:@42897.4]
  wire [63:0] regs_84_io_out; // @[RegFile.scala 66:20:@42897.4]
  wire  regs_84_io_enable; // @[RegFile.scala 66:20:@42897.4]
  wire  regs_85_clock; // @[RegFile.scala 66:20:@42911.4]
  wire  regs_85_reset; // @[RegFile.scala 66:20:@42911.4]
  wire [63:0] regs_85_io_in; // @[RegFile.scala 66:20:@42911.4]
  wire  regs_85_io_reset; // @[RegFile.scala 66:20:@42911.4]
  wire [63:0] regs_85_io_out; // @[RegFile.scala 66:20:@42911.4]
  wire  regs_85_io_enable; // @[RegFile.scala 66:20:@42911.4]
  wire  regs_86_clock; // @[RegFile.scala 66:20:@42925.4]
  wire  regs_86_reset; // @[RegFile.scala 66:20:@42925.4]
  wire [63:0] regs_86_io_in; // @[RegFile.scala 66:20:@42925.4]
  wire  regs_86_io_reset; // @[RegFile.scala 66:20:@42925.4]
  wire [63:0] regs_86_io_out; // @[RegFile.scala 66:20:@42925.4]
  wire  regs_86_io_enable; // @[RegFile.scala 66:20:@42925.4]
  wire  regs_87_clock; // @[RegFile.scala 66:20:@42939.4]
  wire  regs_87_reset; // @[RegFile.scala 66:20:@42939.4]
  wire [63:0] regs_87_io_in; // @[RegFile.scala 66:20:@42939.4]
  wire  regs_87_io_reset; // @[RegFile.scala 66:20:@42939.4]
  wire [63:0] regs_87_io_out; // @[RegFile.scala 66:20:@42939.4]
  wire  regs_87_io_enable; // @[RegFile.scala 66:20:@42939.4]
  wire  regs_88_clock; // @[RegFile.scala 66:20:@42953.4]
  wire  regs_88_reset; // @[RegFile.scala 66:20:@42953.4]
  wire [63:0] regs_88_io_in; // @[RegFile.scala 66:20:@42953.4]
  wire  regs_88_io_reset; // @[RegFile.scala 66:20:@42953.4]
  wire [63:0] regs_88_io_out; // @[RegFile.scala 66:20:@42953.4]
  wire  regs_88_io_enable; // @[RegFile.scala 66:20:@42953.4]
  wire  regs_89_clock; // @[RegFile.scala 66:20:@42967.4]
  wire  regs_89_reset; // @[RegFile.scala 66:20:@42967.4]
  wire [63:0] regs_89_io_in; // @[RegFile.scala 66:20:@42967.4]
  wire  regs_89_io_reset; // @[RegFile.scala 66:20:@42967.4]
  wire [63:0] regs_89_io_out; // @[RegFile.scala 66:20:@42967.4]
  wire  regs_89_io_enable; // @[RegFile.scala 66:20:@42967.4]
  wire  regs_90_clock; // @[RegFile.scala 66:20:@42981.4]
  wire  regs_90_reset; // @[RegFile.scala 66:20:@42981.4]
  wire [63:0] regs_90_io_in; // @[RegFile.scala 66:20:@42981.4]
  wire  regs_90_io_reset; // @[RegFile.scala 66:20:@42981.4]
  wire [63:0] regs_90_io_out; // @[RegFile.scala 66:20:@42981.4]
  wire  regs_90_io_enable; // @[RegFile.scala 66:20:@42981.4]
  wire  regs_91_clock; // @[RegFile.scala 66:20:@42995.4]
  wire  regs_91_reset; // @[RegFile.scala 66:20:@42995.4]
  wire [63:0] regs_91_io_in; // @[RegFile.scala 66:20:@42995.4]
  wire  regs_91_io_reset; // @[RegFile.scala 66:20:@42995.4]
  wire [63:0] regs_91_io_out; // @[RegFile.scala 66:20:@42995.4]
  wire  regs_91_io_enable; // @[RegFile.scala 66:20:@42995.4]
  wire  regs_92_clock; // @[RegFile.scala 66:20:@43009.4]
  wire  regs_92_reset; // @[RegFile.scala 66:20:@43009.4]
  wire [63:0] regs_92_io_in; // @[RegFile.scala 66:20:@43009.4]
  wire  regs_92_io_reset; // @[RegFile.scala 66:20:@43009.4]
  wire [63:0] regs_92_io_out; // @[RegFile.scala 66:20:@43009.4]
  wire  regs_92_io_enable; // @[RegFile.scala 66:20:@43009.4]
  wire  regs_93_clock; // @[RegFile.scala 66:20:@43023.4]
  wire  regs_93_reset; // @[RegFile.scala 66:20:@43023.4]
  wire [63:0] regs_93_io_in; // @[RegFile.scala 66:20:@43023.4]
  wire  regs_93_io_reset; // @[RegFile.scala 66:20:@43023.4]
  wire [63:0] regs_93_io_out; // @[RegFile.scala 66:20:@43023.4]
  wire  regs_93_io_enable; // @[RegFile.scala 66:20:@43023.4]
  wire  regs_94_clock; // @[RegFile.scala 66:20:@43037.4]
  wire  regs_94_reset; // @[RegFile.scala 66:20:@43037.4]
  wire [63:0] regs_94_io_in; // @[RegFile.scala 66:20:@43037.4]
  wire  regs_94_io_reset; // @[RegFile.scala 66:20:@43037.4]
  wire [63:0] regs_94_io_out; // @[RegFile.scala 66:20:@43037.4]
  wire  regs_94_io_enable; // @[RegFile.scala 66:20:@43037.4]
  wire  regs_95_clock; // @[RegFile.scala 66:20:@43051.4]
  wire  regs_95_reset; // @[RegFile.scala 66:20:@43051.4]
  wire [63:0] regs_95_io_in; // @[RegFile.scala 66:20:@43051.4]
  wire  regs_95_io_reset; // @[RegFile.scala 66:20:@43051.4]
  wire [63:0] regs_95_io_out; // @[RegFile.scala 66:20:@43051.4]
  wire  regs_95_io_enable; // @[RegFile.scala 66:20:@43051.4]
  wire  regs_96_clock; // @[RegFile.scala 66:20:@43065.4]
  wire  regs_96_reset; // @[RegFile.scala 66:20:@43065.4]
  wire [63:0] regs_96_io_in; // @[RegFile.scala 66:20:@43065.4]
  wire  regs_96_io_reset; // @[RegFile.scala 66:20:@43065.4]
  wire [63:0] regs_96_io_out; // @[RegFile.scala 66:20:@43065.4]
  wire  regs_96_io_enable; // @[RegFile.scala 66:20:@43065.4]
  wire  regs_97_clock; // @[RegFile.scala 66:20:@43079.4]
  wire  regs_97_reset; // @[RegFile.scala 66:20:@43079.4]
  wire [63:0] regs_97_io_in; // @[RegFile.scala 66:20:@43079.4]
  wire  regs_97_io_reset; // @[RegFile.scala 66:20:@43079.4]
  wire [63:0] regs_97_io_out; // @[RegFile.scala 66:20:@43079.4]
  wire  regs_97_io_enable; // @[RegFile.scala 66:20:@43079.4]
  wire  regs_98_clock; // @[RegFile.scala 66:20:@43093.4]
  wire  regs_98_reset; // @[RegFile.scala 66:20:@43093.4]
  wire [63:0] regs_98_io_in; // @[RegFile.scala 66:20:@43093.4]
  wire  regs_98_io_reset; // @[RegFile.scala 66:20:@43093.4]
  wire [63:0] regs_98_io_out; // @[RegFile.scala 66:20:@43093.4]
  wire  regs_98_io_enable; // @[RegFile.scala 66:20:@43093.4]
  wire  regs_99_clock; // @[RegFile.scala 66:20:@43107.4]
  wire  regs_99_reset; // @[RegFile.scala 66:20:@43107.4]
  wire [63:0] regs_99_io_in; // @[RegFile.scala 66:20:@43107.4]
  wire  regs_99_io_reset; // @[RegFile.scala 66:20:@43107.4]
  wire [63:0] regs_99_io_out; // @[RegFile.scala 66:20:@43107.4]
  wire  regs_99_io_enable; // @[RegFile.scala 66:20:@43107.4]
  wire  regs_100_clock; // @[RegFile.scala 66:20:@43121.4]
  wire  regs_100_reset; // @[RegFile.scala 66:20:@43121.4]
  wire [63:0] regs_100_io_in; // @[RegFile.scala 66:20:@43121.4]
  wire  regs_100_io_reset; // @[RegFile.scala 66:20:@43121.4]
  wire [63:0] regs_100_io_out; // @[RegFile.scala 66:20:@43121.4]
  wire  regs_100_io_enable; // @[RegFile.scala 66:20:@43121.4]
  wire  regs_101_clock; // @[RegFile.scala 66:20:@43135.4]
  wire  regs_101_reset; // @[RegFile.scala 66:20:@43135.4]
  wire [63:0] regs_101_io_in; // @[RegFile.scala 66:20:@43135.4]
  wire  regs_101_io_reset; // @[RegFile.scala 66:20:@43135.4]
  wire [63:0] regs_101_io_out; // @[RegFile.scala 66:20:@43135.4]
  wire  regs_101_io_enable; // @[RegFile.scala 66:20:@43135.4]
  wire  regs_102_clock; // @[RegFile.scala 66:20:@43149.4]
  wire  regs_102_reset; // @[RegFile.scala 66:20:@43149.4]
  wire [63:0] regs_102_io_in; // @[RegFile.scala 66:20:@43149.4]
  wire  regs_102_io_reset; // @[RegFile.scala 66:20:@43149.4]
  wire [63:0] regs_102_io_out; // @[RegFile.scala 66:20:@43149.4]
  wire  regs_102_io_enable; // @[RegFile.scala 66:20:@43149.4]
  wire  regs_103_clock; // @[RegFile.scala 66:20:@43163.4]
  wire  regs_103_reset; // @[RegFile.scala 66:20:@43163.4]
  wire [63:0] regs_103_io_in; // @[RegFile.scala 66:20:@43163.4]
  wire  regs_103_io_reset; // @[RegFile.scala 66:20:@43163.4]
  wire [63:0] regs_103_io_out; // @[RegFile.scala 66:20:@43163.4]
  wire  regs_103_io_enable; // @[RegFile.scala 66:20:@43163.4]
  wire  regs_104_clock; // @[RegFile.scala 66:20:@43177.4]
  wire  regs_104_reset; // @[RegFile.scala 66:20:@43177.4]
  wire [63:0] regs_104_io_in; // @[RegFile.scala 66:20:@43177.4]
  wire  regs_104_io_reset; // @[RegFile.scala 66:20:@43177.4]
  wire [63:0] regs_104_io_out; // @[RegFile.scala 66:20:@43177.4]
  wire  regs_104_io_enable; // @[RegFile.scala 66:20:@43177.4]
  wire  regs_105_clock; // @[RegFile.scala 66:20:@43191.4]
  wire  regs_105_reset; // @[RegFile.scala 66:20:@43191.4]
  wire [63:0] regs_105_io_in; // @[RegFile.scala 66:20:@43191.4]
  wire  regs_105_io_reset; // @[RegFile.scala 66:20:@43191.4]
  wire [63:0] regs_105_io_out; // @[RegFile.scala 66:20:@43191.4]
  wire  regs_105_io_enable; // @[RegFile.scala 66:20:@43191.4]
  wire  regs_106_clock; // @[RegFile.scala 66:20:@43205.4]
  wire  regs_106_reset; // @[RegFile.scala 66:20:@43205.4]
  wire [63:0] regs_106_io_in; // @[RegFile.scala 66:20:@43205.4]
  wire  regs_106_io_reset; // @[RegFile.scala 66:20:@43205.4]
  wire [63:0] regs_106_io_out; // @[RegFile.scala 66:20:@43205.4]
  wire  regs_106_io_enable; // @[RegFile.scala 66:20:@43205.4]
  wire  regs_107_clock; // @[RegFile.scala 66:20:@43219.4]
  wire  regs_107_reset; // @[RegFile.scala 66:20:@43219.4]
  wire [63:0] regs_107_io_in; // @[RegFile.scala 66:20:@43219.4]
  wire  regs_107_io_reset; // @[RegFile.scala 66:20:@43219.4]
  wire [63:0] regs_107_io_out; // @[RegFile.scala 66:20:@43219.4]
  wire  regs_107_io_enable; // @[RegFile.scala 66:20:@43219.4]
  wire  regs_108_clock; // @[RegFile.scala 66:20:@43233.4]
  wire  regs_108_reset; // @[RegFile.scala 66:20:@43233.4]
  wire [63:0] regs_108_io_in; // @[RegFile.scala 66:20:@43233.4]
  wire  regs_108_io_reset; // @[RegFile.scala 66:20:@43233.4]
  wire [63:0] regs_108_io_out; // @[RegFile.scala 66:20:@43233.4]
  wire  regs_108_io_enable; // @[RegFile.scala 66:20:@43233.4]
  wire  regs_109_clock; // @[RegFile.scala 66:20:@43247.4]
  wire  regs_109_reset; // @[RegFile.scala 66:20:@43247.4]
  wire [63:0] regs_109_io_in; // @[RegFile.scala 66:20:@43247.4]
  wire  regs_109_io_reset; // @[RegFile.scala 66:20:@43247.4]
  wire [63:0] regs_109_io_out; // @[RegFile.scala 66:20:@43247.4]
  wire  regs_109_io_enable; // @[RegFile.scala 66:20:@43247.4]
  wire  regs_110_clock; // @[RegFile.scala 66:20:@43261.4]
  wire  regs_110_reset; // @[RegFile.scala 66:20:@43261.4]
  wire [63:0] regs_110_io_in; // @[RegFile.scala 66:20:@43261.4]
  wire  regs_110_io_reset; // @[RegFile.scala 66:20:@43261.4]
  wire [63:0] regs_110_io_out; // @[RegFile.scala 66:20:@43261.4]
  wire  regs_110_io_enable; // @[RegFile.scala 66:20:@43261.4]
  wire  regs_111_clock; // @[RegFile.scala 66:20:@43275.4]
  wire  regs_111_reset; // @[RegFile.scala 66:20:@43275.4]
  wire [63:0] regs_111_io_in; // @[RegFile.scala 66:20:@43275.4]
  wire  regs_111_io_reset; // @[RegFile.scala 66:20:@43275.4]
  wire [63:0] regs_111_io_out; // @[RegFile.scala 66:20:@43275.4]
  wire  regs_111_io_enable; // @[RegFile.scala 66:20:@43275.4]
  wire  regs_112_clock; // @[RegFile.scala 66:20:@43289.4]
  wire  regs_112_reset; // @[RegFile.scala 66:20:@43289.4]
  wire [63:0] regs_112_io_in; // @[RegFile.scala 66:20:@43289.4]
  wire  regs_112_io_reset; // @[RegFile.scala 66:20:@43289.4]
  wire [63:0] regs_112_io_out; // @[RegFile.scala 66:20:@43289.4]
  wire  regs_112_io_enable; // @[RegFile.scala 66:20:@43289.4]
  wire  regs_113_clock; // @[RegFile.scala 66:20:@43303.4]
  wire  regs_113_reset; // @[RegFile.scala 66:20:@43303.4]
  wire [63:0] regs_113_io_in; // @[RegFile.scala 66:20:@43303.4]
  wire  regs_113_io_reset; // @[RegFile.scala 66:20:@43303.4]
  wire [63:0] regs_113_io_out; // @[RegFile.scala 66:20:@43303.4]
  wire  regs_113_io_enable; // @[RegFile.scala 66:20:@43303.4]
  wire  regs_114_clock; // @[RegFile.scala 66:20:@43317.4]
  wire  regs_114_reset; // @[RegFile.scala 66:20:@43317.4]
  wire [63:0] regs_114_io_in; // @[RegFile.scala 66:20:@43317.4]
  wire  regs_114_io_reset; // @[RegFile.scala 66:20:@43317.4]
  wire [63:0] regs_114_io_out; // @[RegFile.scala 66:20:@43317.4]
  wire  regs_114_io_enable; // @[RegFile.scala 66:20:@43317.4]
  wire  regs_115_clock; // @[RegFile.scala 66:20:@43331.4]
  wire  regs_115_reset; // @[RegFile.scala 66:20:@43331.4]
  wire [63:0] regs_115_io_in; // @[RegFile.scala 66:20:@43331.4]
  wire  regs_115_io_reset; // @[RegFile.scala 66:20:@43331.4]
  wire [63:0] regs_115_io_out; // @[RegFile.scala 66:20:@43331.4]
  wire  regs_115_io_enable; // @[RegFile.scala 66:20:@43331.4]
  wire  regs_116_clock; // @[RegFile.scala 66:20:@43345.4]
  wire  regs_116_reset; // @[RegFile.scala 66:20:@43345.4]
  wire [63:0] regs_116_io_in; // @[RegFile.scala 66:20:@43345.4]
  wire  regs_116_io_reset; // @[RegFile.scala 66:20:@43345.4]
  wire [63:0] regs_116_io_out; // @[RegFile.scala 66:20:@43345.4]
  wire  regs_116_io_enable; // @[RegFile.scala 66:20:@43345.4]
  wire  regs_117_clock; // @[RegFile.scala 66:20:@43359.4]
  wire  regs_117_reset; // @[RegFile.scala 66:20:@43359.4]
  wire [63:0] regs_117_io_in; // @[RegFile.scala 66:20:@43359.4]
  wire  regs_117_io_reset; // @[RegFile.scala 66:20:@43359.4]
  wire [63:0] regs_117_io_out; // @[RegFile.scala 66:20:@43359.4]
  wire  regs_117_io_enable; // @[RegFile.scala 66:20:@43359.4]
  wire  regs_118_clock; // @[RegFile.scala 66:20:@43373.4]
  wire  regs_118_reset; // @[RegFile.scala 66:20:@43373.4]
  wire [63:0] regs_118_io_in; // @[RegFile.scala 66:20:@43373.4]
  wire  regs_118_io_reset; // @[RegFile.scala 66:20:@43373.4]
  wire [63:0] regs_118_io_out; // @[RegFile.scala 66:20:@43373.4]
  wire  regs_118_io_enable; // @[RegFile.scala 66:20:@43373.4]
  wire  regs_119_clock; // @[RegFile.scala 66:20:@43387.4]
  wire  regs_119_reset; // @[RegFile.scala 66:20:@43387.4]
  wire [63:0] regs_119_io_in; // @[RegFile.scala 66:20:@43387.4]
  wire  regs_119_io_reset; // @[RegFile.scala 66:20:@43387.4]
  wire [63:0] regs_119_io_out; // @[RegFile.scala 66:20:@43387.4]
  wire  regs_119_io_enable; // @[RegFile.scala 66:20:@43387.4]
  wire  regs_120_clock; // @[RegFile.scala 66:20:@43401.4]
  wire  regs_120_reset; // @[RegFile.scala 66:20:@43401.4]
  wire [63:0] regs_120_io_in; // @[RegFile.scala 66:20:@43401.4]
  wire  regs_120_io_reset; // @[RegFile.scala 66:20:@43401.4]
  wire [63:0] regs_120_io_out; // @[RegFile.scala 66:20:@43401.4]
  wire  regs_120_io_enable; // @[RegFile.scala 66:20:@43401.4]
  wire  regs_121_clock; // @[RegFile.scala 66:20:@43415.4]
  wire  regs_121_reset; // @[RegFile.scala 66:20:@43415.4]
  wire [63:0] regs_121_io_in; // @[RegFile.scala 66:20:@43415.4]
  wire  regs_121_io_reset; // @[RegFile.scala 66:20:@43415.4]
  wire [63:0] regs_121_io_out; // @[RegFile.scala 66:20:@43415.4]
  wire  regs_121_io_enable; // @[RegFile.scala 66:20:@43415.4]
  wire  regs_122_clock; // @[RegFile.scala 66:20:@43429.4]
  wire  regs_122_reset; // @[RegFile.scala 66:20:@43429.4]
  wire [63:0] regs_122_io_in; // @[RegFile.scala 66:20:@43429.4]
  wire  regs_122_io_reset; // @[RegFile.scala 66:20:@43429.4]
  wire [63:0] regs_122_io_out; // @[RegFile.scala 66:20:@43429.4]
  wire  regs_122_io_enable; // @[RegFile.scala 66:20:@43429.4]
  wire  regs_123_clock; // @[RegFile.scala 66:20:@43443.4]
  wire  regs_123_reset; // @[RegFile.scala 66:20:@43443.4]
  wire [63:0] regs_123_io_in; // @[RegFile.scala 66:20:@43443.4]
  wire  regs_123_io_reset; // @[RegFile.scala 66:20:@43443.4]
  wire [63:0] regs_123_io_out; // @[RegFile.scala 66:20:@43443.4]
  wire  regs_123_io_enable; // @[RegFile.scala 66:20:@43443.4]
  wire  regs_124_clock; // @[RegFile.scala 66:20:@43457.4]
  wire  regs_124_reset; // @[RegFile.scala 66:20:@43457.4]
  wire [63:0] regs_124_io_in; // @[RegFile.scala 66:20:@43457.4]
  wire  regs_124_io_reset; // @[RegFile.scala 66:20:@43457.4]
  wire [63:0] regs_124_io_out; // @[RegFile.scala 66:20:@43457.4]
  wire  regs_124_io_enable; // @[RegFile.scala 66:20:@43457.4]
  wire  regs_125_clock; // @[RegFile.scala 66:20:@43471.4]
  wire  regs_125_reset; // @[RegFile.scala 66:20:@43471.4]
  wire [63:0] regs_125_io_in; // @[RegFile.scala 66:20:@43471.4]
  wire  regs_125_io_reset; // @[RegFile.scala 66:20:@43471.4]
  wire [63:0] regs_125_io_out; // @[RegFile.scala 66:20:@43471.4]
  wire  regs_125_io_enable; // @[RegFile.scala 66:20:@43471.4]
  wire  regs_126_clock; // @[RegFile.scala 66:20:@43485.4]
  wire  regs_126_reset; // @[RegFile.scala 66:20:@43485.4]
  wire [63:0] regs_126_io_in; // @[RegFile.scala 66:20:@43485.4]
  wire  regs_126_io_reset; // @[RegFile.scala 66:20:@43485.4]
  wire [63:0] regs_126_io_out; // @[RegFile.scala 66:20:@43485.4]
  wire  regs_126_io_enable; // @[RegFile.scala 66:20:@43485.4]
  wire  regs_127_clock; // @[RegFile.scala 66:20:@43499.4]
  wire  regs_127_reset; // @[RegFile.scala 66:20:@43499.4]
  wire [63:0] regs_127_io_in; // @[RegFile.scala 66:20:@43499.4]
  wire  regs_127_io_reset; // @[RegFile.scala 66:20:@43499.4]
  wire [63:0] regs_127_io_out; // @[RegFile.scala 66:20:@43499.4]
  wire  regs_127_io_enable; // @[RegFile.scala 66:20:@43499.4]
  wire  regs_128_clock; // @[RegFile.scala 66:20:@43513.4]
  wire  regs_128_reset; // @[RegFile.scala 66:20:@43513.4]
  wire [63:0] regs_128_io_in; // @[RegFile.scala 66:20:@43513.4]
  wire  regs_128_io_reset; // @[RegFile.scala 66:20:@43513.4]
  wire [63:0] regs_128_io_out; // @[RegFile.scala 66:20:@43513.4]
  wire  regs_128_io_enable; // @[RegFile.scala 66:20:@43513.4]
  wire  regs_129_clock; // @[RegFile.scala 66:20:@43527.4]
  wire  regs_129_reset; // @[RegFile.scala 66:20:@43527.4]
  wire [63:0] regs_129_io_in; // @[RegFile.scala 66:20:@43527.4]
  wire  regs_129_io_reset; // @[RegFile.scala 66:20:@43527.4]
  wire [63:0] regs_129_io_out; // @[RegFile.scala 66:20:@43527.4]
  wire  regs_129_io_enable; // @[RegFile.scala 66:20:@43527.4]
  wire  regs_130_clock; // @[RegFile.scala 66:20:@43541.4]
  wire  regs_130_reset; // @[RegFile.scala 66:20:@43541.4]
  wire [63:0] regs_130_io_in; // @[RegFile.scala 66:20:@43541.4]
  wire  regs_130_io_reset; // @[RegFile.scala 66:20:@43541.4]
  wire [63:0] regs_130_io_out; // @[RegFile.scala 66:20:@43541.4]
  wire  regs_130_io_enable; // @[RegFile.scala 66:20:@43541.4]
  wire  regs_131_clock; // @[RegFile.scala 66:20:@43555.4]
  wire  regs_131_reset; // @[RegFile.scala 66:20:@43555.4]
  wire [63:0] regs_131_io_in; // @[RegFile.scala 66:20:@43555.4]
  wire  regs_131_io_reset; // @[RegFile.scala 66:20:@43555.4]
  wire [63:0] regs_131_io_out; // @[RegFile.scala 66:20:@43555.4]
  wire  regs_131_io_enable; // @[RegFile.scala 66:20:@43555.4]
  wire  regs_132_clock; // @[RegFile.scala 66:20:@43569.4]
  wire  regs_132_reset; // @[RegFile.scala 66:20:@43569.4]
  wire [63:0] regs_132_io_in; // @[RegFile.scala 66:20:@43569.4]
  wire  regs_132_io_reset; // @[RegFile.scala 66:20:@43569.4]
  wire [63:0] regs_132_io_out; // @[RegFile.scala 66:20:@43569.4]
  wire  regs_132_io_enable; // @[RegFile.scala 66:20:@43569.4]
  wire  regs_133_clock; // @[RegFile.scala 66:20:@43583.4]
  wire  regs_133_reset; // @[RegFile.scala 66:20:@43583.4]
  wire [63:0] regs_133_io_in; // @[RegFile.scala 66:20:@43583.4]
  wire  regs_133_io_reset; // @[RegFile.scala 66:20:@43583.4]
  wire [63:0] regs_133_io_out; // @[RegFile.scala 66:20:@43583.4]
  wire  regs_133_io_enable; // @[RegFile.scala 66:20:@43583.4]
  wire  regs_134_clock; // @[RegFile.scala 66:20:@43597.4]
  wire  regs_134_reset; // @[RegFile.scala 66:20:@43597.4]
  wire [63:0] regs_134_io_in; // @[RegFile.scala 66:20:@43597.4]
  wire  regs_134_io_reset; // @[RegFile.scala 66:20:@43597.4]
  wire [63:0] regs_134_io_out; // @[RegFile.scala 66:20:@43597.4]
  wire  regs_134_io_enable; // @[RegFile.scala 66:20:@43597.4]
  wire  regs_135_clock; // @[RegFile.scala 66:20:@43611.4]
  wire  regs_135_reset; // @[RegFile.scala 66:20:@43611.4]
  wire [63:0] regs_135_io_in; // @[RegFile.scala 66:20:@43611.4]
  wire  regs_135_io_reset; // @[RegFile.scala 66:20:@43611.4]
  wire [63:0] regs_135_io_out; // @[RegFile.scala 66:20:@43611.4]
  wire  regs_135_io_enable; // @[RegFile.scala 66:20:@43611.4]
  wire  regs_136_clock; // @[RegFile.scala 66:20:@43625.4]
  wire  regs_136_reset; // @[RegFile.scala 66:20:@43625.4]
  wire [63:0] regs_136_io_in; // @[RegFile.scala 66:20:@43625.4]
  wire  regs_136_io_reset; // @[RegFile.scala 66:20:@43625.4]
  wire [63:0] regs_136_io_out; // @[RegFile.scala 66:20:@43625.4]
  wire  regs_136_io_enable; // @[RegFile.scala 66:20:@43625.4]
  wire  regs_137_clock; // @[RegFile.scala 66:20:@43639.4]
  wire  regs_137_reset; // @[RegFile.scala 66:20:@43639.4]
  wire [63:0] regs_137_io_in; // @[RegFile.scala 66:20:@43639.4]
  wire  regs_137_io_reset; // @[RegFile.scala 66:20:@43639.4]
  wire [63:0] regs_137_io_out; // @[RegFile.scala 66:20:@43639.4]
  wire  regs_137_io_enable; // @[RegFile.scala 66:20:@43639.4]
  wire  regs_138_clock; // @[RegFile.scala 66:20:@43653.4]
  wire  regs_138_reset; // @[RegFile.scala 66:20:@43653.4]
  wire [63:0] regs_138_io_in; // @[RegFile.scala 66:20:@43653.4]
  wire  regs_138_io_reset; // @[RegFile.scala 66:20:@43653.4]
  wire [63:0] regs_138_io_out; // @[RegFile.scala 66:20:@43653.4]
  wire  regs_138_io_enable; // @[RegFile.scala 66:20:@43653.4]
  wire  regs_139_clock; // @[RegFile.scala 66:20:@43667.4]
  wire  regs_139_reset; // @[RegFile.scala 66:20:@43667.4]
  wire [63:0] regs_139_io_in; // @[RegFile.scala 66:20:@43667.4]
  wire  regs_139_io_reset; // @[RegFile.scala 66:20:@43667.4]
  wire [63:0] regs_139_io_out; // @[RegFile.scala 66:20:@43667.4]
  wire  regs_139_io_enable; // @[RegFile.scala 66:20:@43667.4]
  wire  regs_140_clock; // @[RegFile.scala 66:20:@43681.4]
  wire  regs_140_reset; // @[RegFile.scala 66:20:@43681.4]
  wire [63:0] regs_140_io_in; // @[RegFile.scala 66:20:@43681.4]
  wire  regs_140_io_reset; // @[RegFile.scala 66:20:@43681.4]
  wire [63:0] regs_140_io_out; // @[RegFile.scala 66:20:@43681.4]
  wire  regs_140_io_enable; // @[RegFile.scala 66:20:@43681.4]
  wire  regs_141_clock; // @[RegFile.scala 66:20:@43695.4]
  wire  regs_141_reset; // @[RegFile.scala 66:20:@43695.4]
  wire [63:0] regs_141_io_in; // @[RegFile.scala 66:20:@43695.4]
  wire  regs_141_io_reset; // @[RegFile.scala 66:20:@43695.4]
  wire [63:0] regs_141_io_out; // @[RegFile.scala 66:20:@43695.4]
  wire  regs_141_io_enable; // @[RegFile.scala 66:20:@43695.4]
  wire  regs_142_clock; // @[RegFile.scala 66:20:@43709.4]
  wire  regs_142_reset; // @[RegFile.scala 66:20:@43709.4]
  wire [63:0] regs_142_io_in; // @[RegFile.scala 66:20:@43709.4]
  wire  regs_142_io_reset; // @[RegFile.scala 66:20:@43709.4]
  wire [63:0] regs_142_io_out; // @[RegFile.scala 66:20:@43709.4]
  wire  regs_142_io_enable; // @[RegFile.scala 66:20:@43709.4]
  wire  regs_143_clock; // @[RegFile.scala 66:20:@43723.4]
  wire  regs_143_reset; // @[RegFile.scala 66:20:@43723.4]
  wire [63:0] regs_143_io_in; // @[RegFile.scala 66:20:@43723.4]
  wire  regs_143_io_reset; // @[RegFile.scala 66:20:@43723.4]
  wire [63:0] regs_143_io_out; // @[RegFile.scala 66:20:@43723.4]
  wire  regs_143_io_enable; // @[RegFile.scala 66:20:@43723.4]
  wire  regs_144_clock; // @[RegFile.scala 66:20:@43737.4]
  wire  regs_144_reset; // @[RegFile.scala 66:20:@43737.4]
  wire [63:0] regs_144_io_in; // @[RegFile.scala 66:20:@43737.4]
  wire  regs_144_io_reset; // @[RegFile.scala 66:20:@43737.4]
  wire [63:0] regs_144_io_out; // @[RegFile.scala 66:20:@43737.4]
  wire  regs_144_io_enable; // @[RegFile.scala 66:20:@43737.4]
  wire  regs_145_clock; // @[RegFile.scala 66:20:@43751.4]
  wire  regs_145_reset; // @[RegFile.scala 66:20:@43751.4]
  wire [63:0] regs_145_io_in; // @[RegFile.scala 66:20:@43751.4]
  wire  regs_145_io_reset; // @[RegFile.scala 66:20:@43751.4]
  wire [63:0] regs_145_io_out; // @[RegFile.scala 66:20:@43751.4]
  wire  regs_145_io_enable; // @[RegFile.scala 66:20:@43751.4]
  wire  regs_146_clock; // @[RegFile.scala 66:20:@43765.4]
  wire  regs_146_reset; // @[RegFile.scala 66:20:@43765.4]
  wire [63:0] regs_146_io_in; // @[RegFile.scala 66:20:@43765.4]
  wire  regs_146_io_reset; // @[RegFile.scala 66:20:@43765.4]
  wire [63:0] regs_146_io_out; // @[RegFile.scala 66:20:@43765.4]
  wire  regs_146_io_enable; // @[RegFile.scala 66:20:@43765.4]
  wire  regs_147_clock; // @[RegFile.scala 66:20:@43779.4]
  wire  regs_147_reset; // @[RegFile.scala 66:20:@43779.4]
  wire [63:0] regs_147_io_in; // @[RegFile.scala 66:20:@43779.4]
  wire  regs_147_io_reset; // @[RegFile.scala 66:20:@43779.4]
  wire [63:0] regs_147_io_out; // @[RegFile.scala 66:20:@43779.4]
  wire  regs_147_io_enable; // @[RegFile.scala 66:20:@43779.4]
  wire  regs_148_clock; // @[RegFile.scala 66:20:@43793.4]
  wire  regs_148_reset; // @[RegFile.scala 66:20:@43793.4]
  wire [63:0] regs_148_io_in; // @[RegFile.scala 66:20:@43793.4]
  wire  regs_148_io_reset; // @[RegFile.scala 66:20:@43793.4]
  wire [63:0] regs_148_io_out; // @[RegFile.scala 66:20:@43793.4]
  wire  regs_148_io_enable; // @[RegFile.scala 66:20:@43793.4]
  wire  regs_149_clock; // @[RegFile.scala 66:20:@43807.4]
  wire  regs_149_reset; // @[RegFile.scala 66:20:@43807.4]
  wire [63:0] regs_149_io_in; // @[RegFile.scala 66:20:@43807.4]
  wire  regs_149_io_reset; // @[RegFile.scala 66:20:@43807.4]
  wire [63:0] regs_149_io_out; // @[RegFile.scala 66:20:@43807.4]
  wire  regs_149_io_enable; // @[RegFile.scala 66:20:@43807.4]
  wire  regs_150_clock; // @[RegFile.scala 66:20:@43821.4]
  wire  regs_150_reset; // @[RegFile.scala 66:20:@43821.4]
  wire [63:0] regs_150_io_in; // @[RegFile.scala 66:20:@43821.4]
  wire  regs_150_io_reset; // @[RegFile.scala 66:20:@43821.4]
  wire [63:0] regs_150_io_out; // @[RegFile.scala 66:20:@43821.4]
  wire  regs_150_io_enable; // @[RegFile.scala 66:20:@43821.4]
  wire  regs_151_clock; // @[RegFile.scala 66:20:@43835.4]
  wire  regs_151_reset; // @[RegFile.scala 66:20:@43835.4]
  wire [63:0] regs_151_io_in; // @[RegFile.scala 66:20:@43835.4]
  wire  regs_151_io_reset; // @[RegFile.scala 66:20:@43835.4]
  wire [63:0] regs_151_io_out; // @[RegFile.scala 66:20:@43835.4]
  wire  regs_151_io_enable; // @[RegFile.scala 66:20:@43835.4]
  wire  regs_152_clock; // @[RegFile.scala 66:20:@43849.4]
  wire  regs_152_reset; // @[RegFile.scala 66:20:@43849.4]
  wire [63:0] regs_152_io_in; // @[RegFile.scala 66:20:@43849.4]
  wire  regs_152_io_reset; // @[RegFile.scala 66:20:@43849.4]
  wire [63:0] regs_152_io_out; // @[RegFile.scala 66:20:@43849.4]
  wire  regs_152_io_enable; // @[RegFile.scala 66:20:@43849.4]
  wire  regs_153_clock; // @[RegFile.scala 66:20:@43863.4]
  wire  regs_153_reset; // @[RegFile.scala 66:20:@43863.4]
  wire [63:0] regs_153_io_in; // @[RegFile.scala 66:20:@43863.4]
  wire  regs_153_io_reset; // @[RegFile.scala 66:20:@43863.4]
  wire [63:0] regs_153_io_out; // @[RegFile.scala 66:20:@43863.4]
  wire  regs_153_io_enable; // @[RegFile.scala 66:20:@43863.4]
  wire  regs_154_clock; // @[RegFile.scala 66:20:@43877.4]
  wire  regs_154_reset; // @[RegFile.scala 66:20:@43877.4]
  wire [63:0] regs_154_io_in; // @[RegFile.scala 66:20:@43877.4]
  wire  regs_154_io_reset; // @[RegFile.scala 66:20:@43877.4]
  wire [63:0] regs_154_io_out; // @[RegFile.scala 66:20:@43877.4]
  wire  regs_154_io_enable; // @[RegFile.scala 66:20:@43877.4]
  wire  regs_155_clock; // @[RegFile.scala 66:20:@43891.4]
  wire  regs_155_reset; // @[RegFile.scala 66:20:@43891.4]
  wire [63:0] regs_155_io_in; // @[RegFile.scala 66:20:@43891.4]
  wire  regs_155_io_reset; // @[RegFile.scala 66:20:@43891.4]
  wire [63:0] regs_155_io_out; // @[RegFile.scala 66:20:@43891.4]
  wire  regs_155_io_enable; // @[RegFile.scala 66:20:@43891.4]
  wire  regs_156_clock; // @[RegFile.scala 66:20:@43905.4]
  wire  regs_156_reset; // @[RegFile.scala 66:20:@43905.4]
  wire [63:0] regs_156_io_in; // @[RegFile.scala 66:20:@43905.4]
  wire  regs_156_io_reset; // @[RegFile.scala 66:20:@43905.4]
  wire [63:0] regs_156_io_out; // @[RegFile.scala 66:20:@43905.4]
  wire  regs_156_io_enable; // @[RegFile.scala 66:20:@43905.4]
  wire  regs_157_clock; // @[RegFile.scala 66:20:@43919.4]
  wire  regs_157_reset; // @[RegFile.scala 66:20:@43919.4]
  wire [63:0] regs_157_io_in; // @[RegFile.scala 66:20:@43919.4]
  wire  regs_157_io_reset; // @[RegFile.scala 66:20:@43919.4]
  wire [63:0] regs_157_io_out; // @[RegFile.scala 66:20:@43919.4]
  wire  regs_157_io_enable; // @[RegFile.scala 66:20:@43919.4]
  wire  regs_158_clock; // @[RegFile.scala 66:20:@43933.4]
  wire  regs_158_reset; // @[RegFile.scala 66:20:@43933.4]
  wire [63:0] regs_158_io_in; // @[RegFile.scala 66:20:@43933.4]
  wire  regs_158_io_reset; // @[RegFile.scala 66:20:@43933.4]
  wire [63:0] regs_158_io_out; // @[RegFile.scala 66:20:@43933.4]
  wire  regs_158_io_enable; // @[RegFile.scala 66:20:@43933.4]
  wire  regs_159_clock; // @[RegFile.scala 66:20:@43947.4]
  wire  regs_159_reset; // @[RegFile.scala 66:20:@43947.4]
  wire [63:0] regs_159_io_in; // @[RegFile.scala 66:20:@43947.4]
  wire  regs_159_io_reset; // @[RegFile.scala 66:20:@43947.4]
  wire [63:0] regs_159_io_out; // @[RegFile.scala 66:20:@43947.4]
  wire  regs_159_io_enable; // @[RegFile.scala 66:20:@43947.4]
  wire  regs_160_clock; // @[RegFile.scala 66:20:@43961.4]
  wire  regs_160_reset; // @[RegFile.scala 66:20:@43961.4]
  wire [63:0] regs_160_io_in; // @[RegFile.scala 66:20:@43961.4]
  wire  regs_160_io_reset; // @[RegFile.scala 66:20:@43961.4]
  wire [63:0] regs_160_io_out; // @[RegFile.scala 66:20:@43961.4]
  wire  regs_160_io_enable; // @[RegFile.scala 66:20:@43961.4]
  wire  regs_161_clock; // @[RegFile.scala 66:20:@43975.4]
  wire  regs_161_reset; // @[RegFile.scala 66:20:@43975.4]
  wire [63:0] regs_161_io_in; // @[RegFile.scala 66:20:@43975.4]
  wire  regs_161_io_reset; // @[RegFile.scala 66:20:@43975.4]
  wire [63:0] regs_161_io_out; // @[RegFile.scala 66:20:@43975.4]
  wire  regs_161_io_enable; // @[RegFile.scala 66:20:@43975.4]
  wire  regs_162_clock; // @[RegFile.scala 66:20:@43989.4]
  wire  regs_162_reset; // @[RegFile.scala 66:20:@43989.4]
  wire [63:0] regs_162_io_in; // @[RegFile.scala 66:20:@43989.4]
  wire  regs_162_io_reset; // @[RegFile.scala 66:20:@43989.4]
  wire [63:0] regs_162_io_out; // @[RegFile.scala 66:20:@43989.4]
  wire  regs_162_io_enable; // @[RegFile.scala 66:20:@43989.4]
  wire  regs_163_clock; // @[RegFile.scala 66:20:@44003.4]
  wire  regs_163_reset; // @[RegFile.scala 66:20:@44003.4]
  wire [63:0] regs_163_io_in; // @[RegFile.scala 66:20:@44003.4]
  wire  regs_163_io_reset; // @[RegFile.scala 66:20:@44003.4]
  wire [63:0] regs_163_io_out; // @[RegFile.scala 66:20:@44003.4]
  wire  regs_163_io_enable; // @[RegFile.scala 66:20:@44003.4]
  wire  regs_164_clock; // @[RegFile.scala 66:20:@44017.4]
  wire  regs_164_reset; // @[RegFile.scala 66:20:@44017.4]
  wire [63:0] regs_164_io_in; // @[RegFile.scala 66:20:@44017.4]
  wire  regs_164_io_reset; // @[RegFile.scala 66:20:@44017.4]
  wire [63:0] regs_164_io_out; // @[RegFile.scala 66:20:@44017.4]
  wire  regs_164_io_enable; // @[RegFile.scala 66:20:@44017.4]
  wire  regs_165_clock; // @[RegFile.scala 66:20:@44031.4]
  wire  regs_165_reset; // @[RegFile.scala 66:20:@44031.4]
  wire [63:0] regs_165_io_in; // @[RegFile.scala 66:20:@44031.4]
  wire  regs_165_io_reset; // @[RegFile.scala 66:20:@44031.4]
  wire [63:0] regs_165_io_out; // @[RegFile.scala 66:20:@44031.4]
  wire  regs_165_io_enable; // @[RegFile.scala 66:20:@44031.4]
  wire  regs_166_clock; // @[RegFile.scala 66:20:@44045.4]
  wire  regs_166_reset; // @[RegFile.scala 66:20:@44045.4]
  wire [63:0] regs_166_io_in; // @[RegFile.scala 66:20:@44045.4]
  wire  regs_166_io_reset; // @[RegFile.scala 66:20:@44045.4]
  wire [63:0] regs_166_io_out; // @[RegFile.scala 66:20:@44045.4]
  wire  regs_166_io_enable; // @[RegFile.scala 66:20:@44045.4]
  wire  regs_167_clock; // @[RegFile.scala 66:20:@44059.4]
  wire  regs_167_reset; // @[RegFile.scala 66:20:@44059.4]
  wire [63:0] regs_167_io_in; // @[RegFile.scala 66:20:@44059.4]
  wire  regs_167_io_reset; // @[RegFile.scala 66:20:@44059.4]
  wire [63:0] regs_167_io_out; // @[RegFile.scala 66:20:@44059.4]
  wire  regs_167_io_enable; // @[RegFile.scala 66:20:@44059.4]
  wire  regs_168_clock; // @[RegFile.scala 66:20:@44073.4]
  wire  regs_168_reset; // @[RegFile.scala 66:20:@44073.4]
  wire [63:0] regs_168_io_in; // @[RegFile.scala 66:20:@44073.4]
  wire  regs_168_io_reset; // @[RegFile.scala 66:20:@44073.4]
  wire [63:0] regs_168_io_out; // @[RegFile.scala 66:20:@44073.4]
  wire  regs_168_io_enable; // @[RegFile.scala 66:20:@44073.4]
  wire  regs_169_clock; // @[RegFile.scala 66:20:@44087.4]
  wire  regs_169_reset; // @[RegFile.scala 66:20:@44087.4]
  wire [63:0] regs_169_io_in; // @[RegFile.scala 66:20:@44087.4]
  wire  regs_169_io_reset; // @[RegFile.scala 66:20:@44087.4]
  wire [63:0] regs_169_io_out; // @[RegFile.scala 66:20:@44087.4]
  wire  regs_169_io_enable; // @[RegFile.scala 66:20:@44087.4]
  wire  regs_170_clock; // @[RegFile.scala 66:20:@44101.4]
  wire  regs_170_reset; // @[RegFile.scala 66:20:@44101.4]
  wire [63:0] regs_170_io_in; // @[RegFile.scala 66:20:@44101.4]
  wire  regs_170_io_reset; // @[RegFile.scala 66:20:@44101.4]
  wire [63:0] regs_170_io_out; // @[RegFile.scala 66:20:@44101.4]
  wire  regs_170_io_enable; // @[RegFile.scala 66:20:@44101.4]
  wire  regs_171_clock; // @[RegFile.scala 66:20:@44115.4]
  wire  regs_171_reset; // @[RegFile.scala 66:20:@44115.4]
  wire [63:0] regs_171_io_in; // @[RegFile.scala 66:20:@44115.4]
  wire  regs_171_io_reset; // @[RegFile.scala 66:20:@44115.4]
  wire [63:0] regs_171_io_out; // @[RegFile.scala 66:20:@44115.4]
  wire  regs_171_io_enable; // @[RegFile.scala 66:20:@44115.4]
  wire  regs_172_clock; // @[RegFile.scala 66:20:@44129.4]
  wire  regs_172_reset; // @[RegFile.scala 66:20:@44129.4]
  wire [63:0] regs_172_io_in; // @[RegFile.scala 66:20:@44129.4]
  wire  regs_172_io_reset; // @[RegFile.scala 66:20:@44129.4]
  wire [63:0] regs_172_io_out; // @[RegFile.scala 66:20:@44129.4]
  wire  regs_172_io_enable; // @[RegFile.scala 66:20:@44129.4]
  wire  regs_173_clock; // @[RegFile.scala 66:20:@44143.4]
  wire  regs_173_reset; // @[RegFile.scala 66:20:@44143.4]
  wire [63:0] regs_173_io_in; // @[RegFile.scala 66:20:@44143.4]
  wire  regs_173_io_reset; // @[RegFile.scala 66:20:@44143.4]
  wire [63:0] regs_173_io_out; // @[RegFile.scala 66:20:@44143.4]
  wire  regs_173_io_enable; // @[RegFile.scala 66:20:@44143.4]
  wire  regs_174_clock; // @[RegFile.scala 66:20:@44157.4]
  wire  regs_174_reset; // @[RegFile.scala 66:20:@44157.4]
  wire [63:0] regs_174_io_in; // @[RegFile.scala 66:20:@44157.4]
  wire  regs_174_io_reset; // @[RegFile.scala 66:20:@44157.4]
  wire [63:0] regs_174_io_out; // @[RegFile.scala 66:20:@44157.4]
  wire  regs_174_io_enable; // @[RegFile.scala 66:20:@44157.4]
  wire  regs_175_clock; // @[RegFile.scala 66:20:@44171.4]
  wire  regs_175_reset; // @[RegFile.scala 66:20:@44171.4]
  wire [63:0] regs_175_io_in; // @[RegFile.scala 66:20:@44171.4]
  wire  regs_175_io_reset; // @[RegFile.scala 66:20:@44171.4]
  wire [63:0] regs_175_io_out; // @[RegFile.scala 66:20:@44171.4]
  wire  regs_175_io_enable; // @[RegFile.scala 66:20:@44171.4]
  wire  regs_176_clock; // @[RegFile.scala 66:20:@44185.4]
  wire  regs_176_reset; // @[RegFile.scala 66:20:@44185.4]
  wire [63:0] regs_176_io_in; // @[RegFile.scala 66:20:@44185.4]
  wire  regs_176_io_reset; // @[RegFile.scala 66:20:@44185.4]
  wire [63:0] regs_176_io_out; // @[RegFile.scala 66:20:@44185.4]
  wire  regs_176_io_enable; // @[RegFile.scala 66:20:@44185.4]
  wire  regs_177_clock; // @[RegFile.scala 66:20:@44199.4]
  wire  regs_177_reset; // @[RegFile.scala 66:20:@44199.4]
  wire [63:0] regs_177_io_in; // @[RegFile.scala 66:20:@44199.4]
  wire  regs_177_io_reset; // @[RegFile.scala 66:20:@44199.4]
  wire [63:0] regs_177_io_out; // @[RegFile.scala 66:20:@44199.4]
  wire  regs_177_io_enable; // @[RegFile.scala 66:20:@44199.4]
  wire  regs_178_clock; // @[RegFile.scala 66:20:@44213.4]
  wire  regs_178_reset; // @[RegFile.scala 66:20:@44213.4]
  wire [63:0] regs_178_io_in; // @[RegFile.scala 66:20:@44213.4]
  wire  regs_178_io_reset; // @[RegFile.scala 66:20:@44213.4]
  wire [63:0] regs_178_io_out; // @[RegFile.scala 66:20:@44213.4]
  wire  regs_178_io_enable; // @[RegFile.scala 66:20:@44213.4]
  wire  regs_179_clock; // @[RegFile.scala 66:20:@44227.4]
  wire  regs_179_reset; // @[RegFile.scala 66:20:@44227.4]
  wire [63:0] regs_179_io_in; // @[RegFile.scala 66:20:@44227.4]
  wire  regs_179_io_reset; // @[RegFile.scala 66:20:@44227.4]
  wire [63:0] regs_179_io_out; // @[RegFile.scala 66:20:@44227.4]
  wire  regs_179_io_enable; // @[RegFile.scala 66:20:@44227.4]
  wire  regs_180_clock; // @[RegFile.scala 66:20:@44241.4]
  wire  regs_180_reset; // @[RegFile.scala 66:20:@44241.4]
  wire [63:0] regs_180_io_in; // @[RegFile.scala 66:20:@44241.4]
  wire  regs_180_io_reset; // @[RegFile.scala 66:20:@44241.4]
  wire [63:0] regs_180_io_out; // @[RegFile.scala 66:20:@44241.4]
  wire  regs_180_io_enable; // @[RegFile.scala 66:20:@44241.4]
  wire  regs_181_clock; // @[RegFile.scala 66:20:@44255.4]
  wire  regs_181_reset; // @[RegFile.scala 66:20:@44255.4]
  wire [63:0] regs_181_io_in; // @[RegFile.scala 66:20:@44255.4]
  wire  regs_181_io_reset; // @[RegFile.scala 66:20:@44255.4]
  wire [63:0] regs_181_io_out; // @[RegFile.scala 66:20:@44255.4]
  wire  regs_181_io_enable; // @[RegFile.scala 66:20:@44255.4]
  wire  regs_182_clock; // @[RegFile.scala 66:20:@44269.4]
  wire  regs_182_reset; // @[RegFile.scala 66:20:@44269.4]
  wire [63:0] regs_182_io_in; // @[RegFile.scala 66:20:@44269.4]
  wire  regs_182_io_reset; // @[RegFile.scala 66:20:@44269.4]
  wire [63:0] regs_182_io_out; // @[RegFile.scala 66:20:@44269.4]
  wire  regs_182_io_enable; // @[RegFile.scala 66:20:@44269.4]
  wire  regs_183_clock; // @[RegFile.scala 66:20:@44283.4]
  wire  regs_183_reset; // @[RegFile.scala 66:20:@44283.4]
  wire [63:0] regs_183_io_in; // @[RegFile.scala 66:20:@44283.4]
  wire  regs_183_io_reset; // @[RegFile.scala 66:20:@44283.4]
  wire [63:0] regs_183_io_out; // @[RegFile.scala 66:20:@44283.4]
  wire  regs_183_io_enable; // @[RegFile.scala 66:20:@44283.4]
  wire  regs_184_clock; // @[RegFile.scala 66:20:@44297.4]
  wire  regs_184_reset; // @[RegFile.scala 66:20:@44297.4]
  wire [63:0] regs_184_io_in; // @[RegFile.scala 66:20:@44297.4]
  wire  regs_184_io_reset; // @[RegFile.scala 66:20:@44297.4]
  wire [63:0] regs_184_io_out; // @[RegFile.scala 66:20:@44297.4]
  wire  regs_184_io_enable; // @[RegFile.scala 66:20:@44297.4]
  wire  regs_185_clock; // @[RegFile.scala 66:20:@44311.4]
  wire  regs_185_reset; // @[RegFile.scala 66:20:@44311.4]
  wire [63:0] regs_185_io_in; // @[RegFile.scala 66:20:@44311.4]
  wire  regs_185_io_reset; // @[RegFile.scala 66:20:@44311.4]
  wire [63:0] regs_185_io_out; // @[RegFile.scala 66:20:@44311.4]
  wire  regs_185_io_enable; // @[RegFile.scala 66:20:@44311.4]
  wire  regs_186_clock; // @[RegFile.scala 66:20:@44325.4]
  wire  regs_186_reset; // @[RegFile.scala 66:20:@44325.4]
  wire [63:0] regs_186_io_in; // @[RegFile.scala 66:20:@44325.4]
  wire  regs_186_io_reset; // @[RegFile.scala 66:20:@44325.4]
  wire [63:0] regs_186_io_out; // @[RegFile.scala 66:20:@44325.4]
  wire  regs_186_io_enable; // @[RegFile.scala 66:20:@44325.4]
  wire  regs_187_clock; // @[RegFile.scala 66:20:@44339.4]
  wire  regs_187_reset; // @[RegFile.scala 66:20:@44339.4]
  wire [63:0] regs_187_io_in; // @[RegFile.scala 66:20:@44339.4]
  wire  regs_187_io_reset; // @[RegFile.scala 66:20:@44339.4]
  wire [63:0] regs_187_io_out; // @[RegFile.scala 66:20:@44339.4]
  wire  regs_187_io_enable; // @[RegFile.scala 66:20:@44339.4]
  wire  regs_188_clock; // @[RegFile.scala 66:20:@44353.4]
  wire  regs_188_reset; // @[RegFile.scala 66:20:@44353.4]
  wire [63:0] regs_188_io_in; // @[RegFile.scala 66:20:@44353.4]
  wire  regs_188_io_reset; // @[RegFile.scala 66:20:@44353.4]
  wire [63:0] regs_188_io_out; // @[RegFile.scala 66:20:@44353.4]
  wire  regs_188_io_enable; // @[RegFile.scala 66:20:@44353.4]
  wire  regs_189_clock; // @[RegFile.scala 66:20:@44367.4]
  wire  regs_189_reset; // @[RegFile.scala 66:20:@44367.4]
  wire [63:0] regs_189_io_in; // @[RegFile.scala 66:20:@44367.4]
  wire  regs_189_io_reset; // @[RegFile.scala 66:20:@44367.4]
  wire [63:0] regs_189_io_out; // @[RegFile.scala 66:20:@44367.4]
  wire  regs_189_io_enable; // @[RegFile.scala 66:20:@44367.4]
  wire  regs_190_clock; // @[RegFile.scala 66:20:@44381.4]
  wire  regs_190_reset; // @[RegFile.scala 66:20:@44381.4]
  wire [63:0] regs_190_io_in; // @[RegFile.scala 66:20:@44381.4]
  wire  regs_190_io_reset; // @[RegFile.scala 66:20:@44381.4]
  wire [63:0] regs_190_io_out; // @[RegFile.scala 66:20:@44381.4]
  wire  regs_190_io_enable; // @[RegFile.scala 66:20:@44381.4]
  wire  regs_191_clock; // @[RegFile.scala 66:20:@44395.4]
  wire  regs_191_reset; // @[RegFile.scala 66:20:@44395.4]
  wire [63:0] regs_191_io_in; // @[RegFile.scala 66:20:@44395.4]
  wire  regs_191_io_reset; // @[RegFile.scala 66:20:@44395.4]
  wire [63:0] regs_191_io_out; // @[RegFile.scala 66:20:@44395.4]
  wire  regs_191_io_enable; // @[RegFile.scala 66:20:@44395.4]
  wire  regs_192_clock; // @[RegFile.scala 66:20:@44409.4]
  wire  regs_192_reset; // @[RegFile.scala 66:20:@44409.4]
  wire [63:0] regs_192_io_in; // @[RegFile.scala 66:20:@44409.4]
  wire  regs_192_io_reset; // @[RegFile.scala 66:20:@44409.4]
  wire [63:0] regs_192_io_out; // @[RegFile.scala 66:20:@44409.4]
  wire  regs_192_io_enable; // @[RegFile.scala 66:20:@44409.4]
  wire  regs_193_clock; // @[RegFile.scala 66:20:@44423.4]
  wire  regs_193_reset; // @[RegFile.scala 66:20:@44423.4]
  wire [63:0] regs_193_io_in; // @[RegFile.scala 66:20:@44423.4]
  wire  regs_193_io_reset; // @[RegFile.scala 66:20:@44423.4]
  wire [63:0] regs_193_io_out; // @[RegFile.scala 66:20:@44423.4]
  wire  regs_193_io_enable; // @[RegFile.scala 66:20:@44423.4]
  wire  regs_194_clock; // @[RegFile.scala 66:20:@44437.4]
  wire  regs_194_reset; // @[RegFile.scala 66:20:@44437.4]
  wire [63:0] regs_194_io_in; // @[RegFile.scala 66:20:@44437.4]
  wire  regs_194_io_reset; // @[RegFile.scala 66:20:@44437.4]
  wire [63:0] regs_194_io_out; // @[RegFile.scala 66:20:@44437.4]
  wire  regs_194_io_enable; // @[RegFile.scala 66:20:@44437.4]
  wire  regs_195_clock; // @[RegFile.scala 66:20:@44451.4]
  wire  regs_195_reset; // @[RegFile.scala 66:20:@44451.4]
  wire [63:0] regs_195_io_in; // @[RegFile.scala 66:20:@44451.4]
  wire  regs_195_io_reset; // @[RegFile.scala 66:20:@44451.4]
  wire [63:0] regs_195_io_out; // @[RegFile.scala 66:20:@44451.4]
  wire  regs_195_io_enable; // @[RegFile.scala 66:20:@44451.4]
  wire  regs_196_clock; // @[RegFile.scala 66:20:@44465.4]
  wire  regs_196_reset; // @[RegFile.scala 66:20:@44465.4]
  wire [63:0] regs_196_io_in; // @[RegFile.scala 66:20:@44465.4]
  wire  regs_196_io_reset; // @[RegFile.scala 66:20:@44465.4]
  wire [63:0] regs_196_io_out; // @[RegFile.scala 66:20:@44465.4]
  wire  regs_196_io_enable; // @[RegFile.scala 66:20:@44465.4]
  wire  regs_197_clock; // @[RegFile.scala 66:20:@44479.4]
  wire  regs_197_reset; // @[RegFile.scala 66:20:@44479.4]
  wire [63:0] regs_197_io_in; // @[RegFile.scala 66:20:@44479.4]
  wire  regs_197_io_reset; // @[RegFile.scala 66:20:@44479.4]
  wire [63:0] regs_197_io_out; // @[RegFile.scala 66:20:@44479.4]
  wire  regs_197_io_enable; // @[RegFile.scala 66:20:@44479.4]
  wire  regs_198_clock; // @[RegFile.scala 66:20:@44493.4]
  wire  regs_198_reset; // @[RegFile.scala 66:20:@44493.4]
  wire [63:0] regs_198_io_in; // @[RegFile.scala 66:20:@44493.4]
  wire  regs_198_io_reset; // @[RegFile.scala 66:20:@44493.4]
  wire [63:0] regs_198_io_out; // @[RegFile.scala 66:20:@44493.4]
  wire  regs_198_io_enable; // @[RegFile.scala 66:20:@44493.4]
  wire  regs_199_clock; // @[RegFile.scala 66:20:@44507.4]
  wire  regs_199_reset; // @[RegFile.scala 66:20:@44507.4]
  wire [63:0] regs_199_io_in; // @[RegFile.scala 66:20:@44507.4]
  wire  regs_199_io_reset; // @[RegFile.scala 66:20:@44507.4]
  wire [63:0] regs_199_io_out; // @[RegFile.scala 66:20:@44507.4]
  wire  regs_199_io_enable; // @[RegFile.scala 66:20:@44507.4]
  wire  regs_200_clock; // @[RegFile.scala 66:20:@44521.4]
  wire  regs_200_reset; // @[RegFile.scala 66:20:@44521.4]
  wire [63:0] regs_200_io_in; // @[RegFile.scala 66:20:@44521.4]
  wire  regs_200_io_reset; // @[RegFile.scala 66:20:@44521.4]
  wire [63:0] regs_200_io_out; // @[RegFile.scala 66:20:@44521.4]
  wire  regs_200_io_enable; // @[RegFile.scala 66:20:@44521.4]
  wire  regs_201_clock; // @[RegFile.scala 66:20:@44535.4]
  wire  regs_201_reset; // @[RegFile.scala 66:20:@44535.4]
  wire [63:0] regs_201_io_in; // @[RegFile.scala 66:20:@44535.4]
  wire  regs_201_io_reset; // @[RegFile.scala 66:20:@44535.4]
  wire [63:0] regs_201_io_out; // @[RegFile.scala 66:20:@44535.4]
  wire  regs_201_io_enable; // @[RegFile.scala 66:20:@44535.4]
  wire  regs_202_clock; // @[RegFile.scala 66:20:@44549.4]
  wire  regs_202_reset; // @[RegFile.scala 66:20:@44549.4]
  wire [63:0] regs_202_io_in; // @[RegFile.scala 66:20:@44549.4]
  wire  regs_202_io_reset; // @[RegFile.scala 66:20:@44549.4]
  wire [63:0] regs_202_io_out; // @[RegFile.scala 66:20:@44549.4]
  wire  regs_202_io_enable; // @[RegFile.scala 66:20:@44549.4]
  wire  regs_203_clock; // @[RegFile.scala 66:20:@44563.4]
  wire  regs_203_reset; // @[RegFile.scala 66:20:@44563.4]
  wire [63:0] regs_203_io_in; // @[RegFile.scala 66:20:@44563.4]
  wire  regs_203_io_reset; // @[RegFile.scala 66:20:@44563.4]
  wire [63:0] regs_203_io_out; // @[RegFile.scala 66:20:@44563.4]
  wire  regs_203_io_enable; // @[RegFile.scala 66:20:@44563.4]
  wire  regs_204_clock; // @[RegFile.scala 66:20:@44577.4]
  wire  regs_204_reset; // @[RegFile.scala 66:20:@44577.4]
  wire [63:0] regs_204_io_in; // @[RegFile.scala 66:20:@44577.4]
  wire  regs_204_io_reset; // @[RegFile.scala 66:20:@44577.4]
  wire [63:0] regs_204_io_out; // @[RegFile.scala 66:20:@44577.4]
  wire  regs_204_io_enable; // @[RegFile.scala 66:20:@44577.4]
  wire  regs_205_clock; // @[RegFile.scala 66:20:@44591.4]
  wire  regs_205_reset; // @[RegFile.scala 66:20:@44591.4]
  wire [63:0] regs_205_io_in; // @[RegFile.scala 66:20:@44591.4]
  wire  regs_205_io_reset; // @[RegFile.scala 66:20:@44591.4]
  wire [63:0] regs_205_io_out; // @[RegFile.scala 66:20:@44591.4]
  wire  regs_205_io_enable; // @[RegFile.scala 66:20:@44591.4]
  wire  regs_206_clock; // @[RegFile.scala 66:20:@44605.4]
  wire  regs_206_reset; // @[RegFile.scala 66:20:@44605.4]
  wire [63:0] regs_206_io_in; // @[RegFile.scala 66:20:@44605.4]
  wire  regs_206_io_reset; // @[RegFile.scala 66:20:@44605.4]
  wire [63:0] regs_206_io_out; // @[RegFile.scala 66:20:@44605.4]
  wire  regs_206_io_enable; // @[RegFile.scala 66:20:@44605.4]
  wire  regs_207_clock; // @[RegFile.scala 66:20:@44619.4]
  wire  regs_207_reset; // @[RegFile.scala 66:20:@44619.4]
  wire [63:0] regs_207_io_in; // @[RegFile.scala 66:20:@44619.4]
  wire  regs_207_io_reset; // @[RegFile.scala 66:20:@44619.4]
  wire [63:0] regs_207_io_out; // @[RegFile.scala 66:20:@44619.4]
  wire  regs_207_io_enable; // @[RegFile.scala 66:20:@44619.4]
  wire  regs_208_clock; // @[RegFile.scala 66:20:@44633.4]
  wire  regs_208_reset; // @[RegFile.scala 66:20:@44633.4]
  wire [63:0] regs_208_io_in; // @[RegFile.scala 66:20:@44633.4]
  wire  regs_208_io_reset; // @[RegFile.scala 66:20:@44633.4]
  wire [63:0] regs_208_io_out; // @[RegFile.scala 66:20:@44633.4]
  wire  regs_208_io_enable; // @[RegFile.scala 66:20:@44633.4]
  wire  regs_209_clock; // @[RegFile.scala 66:20:@44647.4]
  wire  regs_209_reset; // @[RegFile.scala 66:20:@44647.4]
  wire [63:0] regs_209_io_in; // @[RegFile.scala 66:20:@44647.4]
  wire  regs_209_io_reset; // @[RegFile.scala 66:20:@44647.4]
  wire [63:0] regs_209_io_out; // @[RegFile.scala 66:20:@44647.4]
  wire  regs_209_io_enable; // @[RegFile.scala 66:20:@44647.4]
  wire  regs_210_clock; // @[RegFile.scala 66:20:@44661.4]
  wire  regs_210_reset; // @[RegFile.scala 66:20:@44661.4]
  wire [63:0] regs_210_io_in; // @[RegFile.scala 66:20:@44661.4]
  wire  regs_210_io_reset; // @[RegFile.scala 66:20:@44661.4]
  wire [63:0] regs_210_io_out; // @[RegFile.scala 66:20:@44661.4]
  wire  regs_210_io_enable; // @[RegFile.scala 66:20:@44661.4]
  wire  regs_211_clock; // @[RegFile.scala 66:20:@44675.4]
  wire  regs_211_reset; // @[RegFile.scala 66:20:@44675.4]
  wire [63:0] regs_211_io_in; // @[RegFile.scala 66:20:@44675.4]
  wire  regs_211_io_reset; // @[RegFile.scala 66:20:@44675.4]
  wire [63:0] regs_211_io_out; // @[RegFile.scala 66:20:@44675.4]
  wire  regs_211_io_enable; // @[RegFile.scala 66:20:@44675.4]
  wire  regs_212_clock; // @[RegFile.scala 66:20:@44689.4]
  wire  regs_212_reset; // @[RegFile.scala 66:20:@44689.4]
  wire [63:0] regs_212_io_in; // @[RegFile.scala 66:20:@44689.4]
  wire  regs_212_io_reset; // @[RegFile.scala 66:20:@44689.4]
  wire [63:0] regs_212_io_out; // @[RegFile.scala 66:20:@44689.4]
  wire  regs_212_io_enable; // @[RegFile.scala 66:20:@44689.4]
  wire  regs_213_clock; // @[RegFile.scala 66:20:@44703.4]
  wire  regs_213_reset; // @[RegFile.scala 66:20:@44703.4]
  wire [63:0] regs_213_io_in; // @[RegFile.scala 66:20:@44703.4]
  wire  regs_213_io_reset; // @[RegFile.scala 66:20:@44703.4]
  wire [63:0] regs_213_io_out; // @[RegFile.scala 66:20:@44703.4]
  wire  regs_213_io_enable; // @[RegFile.scala 66:20:@44703.4]
  wire  regs_214_clock; // @[RegFile.scala 66:20:@44717.4]
  wire  regs_214_reset; // @[RegFile.scala 66:20:@44717.4]
  wire [63:0] regs_214_io_in; // @[RegFile.scala 66:20:@44717.4]
  wire  regs_214_io_reset; // @[RegFile.scala 66:20:@44717.4]
  wire [63:0] regs_214_io_out; // @[RegFile.scala 66:20:@44717.4]
  wire  regs_214_io_enable; // @[RegFile.scala 66:20:@44717.4]
  wire  regs_215_clock; // @[RegFile.scala 66:20:@44731.4]
  wire  regs_215_reset; // @[RegFile.scala 66:20:@44731.4]
  wire [63:0] regs_215_io_in; // @[RegFile.scala 66:20:@44731.4]
  wire  regs_215_io_reset; // @[RegFile.scala 66:20:@44731.4]
  wire [63:0] regs_215_io_out; // @[RegFile.scala 66:20:@44731.4]
  wire  regs_215_io_enable; // @[RegFile.scala 66:20:@44731.4]
  wire  regs_216_clock; // @[RegFile.scala 66:20:@44745.4]
  wire  regs_216_reset; // @[RegFile.scala 66:20:@44745.4]
  wire [63:0] regs_216_io_in; // @[RegFile.scala 66:20:@44745.4]
  wire  regs_216_io_reset; // @[RegFile.scala 66:20:@44745.4]
  wire [63:0] regs_216_io_out; // @[RegFile.scala 66:20:@44745.4]
  wire  regs_216_io_enable; // @[RegFile.scala 66:20:@44745.4]
  wire  regs_217_clock; // @[RegFile.scala 66:20:@44759.4]
  wire  regs_217_reset; // @[RegFile.scala 66:20:@44759.4]
  wire [63:0] regs_217_io_in; // @[RegFile.scala 66:20:@44759.4]
  wire  regs_217_io_reset; // @[RegFile.scala 66:20:@44759.4]
  wire [63:0] regs_217_io_out; // @[RegFile.scala 66:20:@44759.4]
  wire  regs_217_io_enable; // @[RegFile.scala 66:20:@44759.4]
  wire  regs_218_clock; // @[RegFile.scala 66:20:@44773.4]
  wire  regs_218_reset; // @[RegFile.scala 66:20:@44773.4]
  wire [63:0] regs_218_io_in; // @[RegFile.scala 66:20:@44773.4]
  wire  regs_218_io_reset; // @[RegFile.scala 66:20:@44773.4]
  wire [63:0] regs_218_io_out; // @[RegFile.scala 66:20:@44773.4]
  wire  regs_218_io_enable; // @[RegFile.scala 66:20:@44773.4]
  wire  regs_219_clock; // @[RegFile.scala 66:20:@44787.4]
  wire  regs_219_reset; // @[RegFile.scala 66:20:@44787.4]
  wire [63:0] regs_219_io_in; // @[RegFile.scala 66:20:@44787.4]
  wire  regs_219_io_reset; // @[RegFile.scala 66:20:@44787.4]
  wire [63:0] regs_219_io_out; // @[RegFile.scala 66:20:@44787.4]
  wire  regs_219_io_enable; // @[RegFile.scala 66:20:@44787.4]
  wire  regs_220_clock; // @[RegFile.scala 66:20:@44801.4]
  wire  regs_220_reset; // @[RegFile.scala 66:20:@44801.4]
  wire [63:0] regs_220_io_in; // @[RegFile.scala 66:20:@44801.4]
  wire  regs_220_io_reset; // @[RegFile.scala 66:20:@44801.4]
  wire [63:0] regs_220_io_out; // @[RegFile.scala 66:20:@44801.4]
  wire  regs_220_io_enable; // @[RegFile.scala 66:20:@44801.4]
  wire  regs_221_clock; // @[RegFile.scala 66:20:@44815.4]
  wire  regs_221_reset; // @[RegFile.scala 66:20:@44815.4]
  wire [63:0] regs_221_io_in; // @[RegFile.scala 66:20:@44815.4]
  wire  regs_221_io_reset; // @[RegFile.scala 66:20:@44815.4]
  wire [63:0] regs_221_io_out; // @[RegFile.scala 66:20:@44815.4]
  wire  regs_221_io_enable; // @[RegFile.scala 66:20:@44815.4]
  wire  regs_222_clock; // @[RegFile.scala 66:20:@44829.4]
  wire  regs_222_reset; // @[RegFile.scala 66:20:@44829.4]
  wire [63:0] regs_222_io_in; // @[RegFile.scala 66:20:@44829.4]
  wire  regs_222_io_reset; // @[RegFile.scala 66:20:@44829.4]
  wire [63:0] regs_222_io_out; // @[RegFile.scala 66:20:@44829.4]
  wire  regs_222_io_enable; // @[RegFile.scala 66:20:@44829.4]
  wire  regs_223_clock; // @[RegFile.scala 66:20:@44843.4]
  wire  regs_223_reset; // @[RegFile.scala 66:20:@44843.4]
  wire [63:0] regs_223_io_in; // @[RegFile.scala 66:20:@44843.4]
  wire  regs_223_io_reset; // @[RegFile.scala 66:20:@44843.4]
  wire [63:0] regs_223_io_out; // @[RegFile.scala 66:20:@44843.4]
  wire  regs_223_io_enable; // @[RegFile.scala 66:20:@44843.4]
  wire  regs_224_clock; // @[RegFile.scala 66:20:@44857.4]
  wire  regs_224_reset; // @[RegFile.scala 66:20:@44857.4]
  wire [63:0] regs_224_io_in; // @[RegFile.scala 66:20:@44857.4]
  wire  regs_224_io_reset; // @[RegFile.scala 66:20:@44857.4]
  wire [63:0] regs_224_io_out; // @[RegFile.scala 66:20:@44857.4]
  wire  regs_224_io_enable; // @[RegFile.scala 66:20:@44857.4]
  wire  regs_225_clock; // @[RegFile.scala 66:20:@44871.4]
  wire  regs_225_reset; // @[RegFile.scala 66:20:@44871.4]
  wire [63:0] regs_225_io_in; // @[RegFile.scala 66:20:@44871.4]
  wire  regs_225_io_reset; // @[RegFile.scala 66:20:@44871.4]
  wire [63:0] regs_225_io_out; // @[RegFile.scala 66:20:@44871.4]
  wire  regs_225_io_enable; // @[RegFile.scala 66:20:@44871.4]
  wire  regs_226_clock; // @[RegFile.scala 66:20:@44885.4]
  wire  regs_226_reset; // @[RegFile.scala 66:20:@44885.4]
  wire [63:0] regs_226_io_in; // @[RegFile.scala 66:20:@44885.4]
  wire  regs_226_io_reset; // @[RegFile.scala 66:20:@44885.4]
  wire [63:0] regs_226_io_out; // @[RegFile.scala 66:20:@44885.4]
  wire  regs_226_io_enable; // @[RegFile.scala 66:20:@44885.4]
  wire  regs_227_clock; // @[RegFile.scala 66:20:@44899.4]
  wire  regs_227_reset; // @[RegFile.scala 66:20:@44899.4]
  wire [63:0] regs_227_io_in; // @[RegFile.scala 66:20:@44899.4]
  wire  regs_227_io_reset; // @[RegFile.scala 66:20:@44899.4]
  wire [63:0] regs_227_io_out; // @[RegFile.scala 66:20:@44899.4]
  wire  regs_227_io_enable; // @[RegFile.scala 66:20:@44899.4]
  wire  regs_228_clock; // @[RegFile.scala 66:20:@44913.4]
  wire  regs_228_reset; // @[RegFile.scala 66:20:@44913.4]
  wire [63:0] regs_228_io_in; // @[RegFile.scala 66:20:@44913.4]
  wire  regs_228_io_reset; // @[RegFile.scala 66:20:@44913.4]
  wire [63:0] regs_228_io_out; // @[RegFile.scala 66:20:@44913.4]
  wire  regs_228_io_enable; // @[RegFile.scala 66:20:@44913.4]
  wire  regs_229_clock; // @[RegFile.scala 66:20:@44927.4]
  wire  regs_229_reset; // @[RegFile.scala 66:20:@44927.4]
  wire [63:0] regs_229_io_in; // @[RegFile.scala 66:20:@44927.4]
  wire  regs_229_io_reset; // @[RegFile.scala 66:20:@44927.4]
  wire [63:0] regs_229_io_out; // @[RegFile.scala 66:20:@44927.4]
  wire  regs_229_io_enable; // @[RegFile.scala 66:20:@44927.4]
  wire  regs_230_clock; // @[RegFile.scala 66:20:@44941.4]
  wire  regs_230_reset; // @[RegFile.scala 66:20:@44941.4]
  wire [63:0] regs_230_io_in; // @[RegFile.scala 66:20:@44941.4]
  wire  regs_230_io_reset; // @[RegFile.scala 66:20:@44941.4]
  wire [63:0] regs_230_io_out; // @[RegFile.scala 66:20:@44941.4]
  wire  regs_230_io_enable; // @[RegFile.scala 66:20:@44941.4]
  wire  regs_231_clock; // @[RegFile.scala 66:20:@44955.4]
  wire  regs_231_reset; // @[RegFile.scala 66:20:@44955.4]
  wire [63:0] regs_231_io_in; // @[RegFile.scala 66:20:@44955.4]
  wire  regs_231_io_reset; // @[RegFile.scala 66:20:@44955.4]
  wire [63:0] regs_231_io_out; // @[RegFile.scala 66:20:@44955.4]
  wire  regs_231_io_enable; // @[RegFile.scala 66:20:@44955.4]
  wire  regs_232_clock; // @[RegFile.scala 66:20:@44969.4]
  wire  regs_232_reset; // @[RegFile.scala 66:20:@44969.4]
  wire [63:0] regs_232_io_in; // @[RegFile.scala 66:20:@44969.4]
  wire  regs_232_io_reset; // @[RegFile.scala 66:20:@44969.4]
  wire [63:0] regs_232_io_out; // @[RegFile.scala 66:20:@44969.4]
  wire  regs_232_io_enable; // @[RegFile.scala 66:20:@44969.4]
  wire  regs_233_clock; // @[RegFile.scala 66:20:@44983.4]
  wire  regs_233_reset; // @[RegFile.scala 66:20:@44983.4]
  wire [63:0] regs_233_io_in; // @[RegFile.scala 66:20:@44983.4]
  wire  regs_233_io_reset; // @[RegFile.scala 66:20:@44983.4]
  wire [63:0] regs_233_io_out; // @[RegFile.scala 66:20:@44983.4]
  wire  regs_233_io_enable; // @[RegFile.scala 66:20:@44983.4]
  wire  regs_234_clock; // @[RegFile.scala 66:20:@44997.4]
  wire  regs_234_reset; // @[RegFile.scala 66:20:@44997.4]
  wire [63:0] regs_234_io_in; // @[RegFile.scala 66:20:@44997.4]
  wire  regs_234_io_reset; // @[RegFile.scala 66:20:@44997.4]
  wire [63:0] regs_234_io_out; // @[RegFile.scala 66:20:@44997.4]
  wire  regs_234_io_enable; // @[RegFile.scala 66:20:@44997.4]
  wire  regs_235_clock; // @[RegFile.scala 66:20:@45011.4]
  wire  regs_235_reset; // @[RegFile.scala 66:20:@45011.4]
  wire [63:0] regs_235_io_in; // @[RegFile.scala 66:20:@45011.4]
  wire  regs_235_io_reset; // @[RegFile.scala 66:20:@45011.4]
  wire [63:0] regs_235_io_out; // @[RegFile.scala 66:20:@45011.4]
  wire  regs_235_io_enable; // @[RegFile.scala 66:20:@45011.4]
  wire  regs_236_clock; // @[RegFile.scala 66:20:@45025.4]
  wire  regs_236_reset; // @[RegFile.scala 66:20:@45025.4]
  wire [63:0] regs_236_io_in; // @[RegFile.scala 66:20:@45025.4]
  wire  regs_236_io_reset; // @[RegFile.scala 66:20:@45025.4]
  wire [63:0] regs_236_io_out; // @[RegFile.scala 66:20:@45025.4]
  wire  regs_236_io_enable; // @[RegFile.scala 66:20:@45025.4]
  wire  regs_237_clock; // @[RegFile.scala 66:20:@45039.4]
  wire  regs_237_reset; // @[RegFile.scala 66:20:@45039.4]
  wire [63:0] regs_237_io_in; // @[RegFile.scala 66:20:@45039.4]
  wire  regs_237_io_reset; // @[RegFile.scala 66:20:@45039.4]
  wire [63:0] regs_237_io_out; // @[RegFile.scala 66:20:@45039.4]
  wire  regs_237_io_enable; // @[RegFile.scala 66:20:@45039.4]
  wire  regs_238_clock; // @[RegFile.scala 66:20:@45053.4]
  wire  regs_238_reset; // @[RegFile.scala 66:20:@45053.4]
  wire [63:0] regs_238_io_in; // @[RegFile.scala 66:20:@45053.4]
  wire  regs_238_io_reset; // @[RegFile.scala 66:20:@45053.4]
  wire [63:0] regs_238_io_out; // @[RegFile.scala 66:20:@45053.4]
  wire  regs_238_io_enable; // @[RegFile.scala 66:20:@45053.4]
  wire  regs_239_clock; // @[RegFile.scala 66:20:@45067.4]
  wire  regs_239_reset; // @[RegFile.scala 66:20:@45067.4]
  wire [63:0] regs_239_io_in; // @[RegFile.scala 66:20:@45067.4]
  wire  regs_239_io_reset; // @[RegFile.scala 66:20:@45067.4]
  wire [63:0] regs_239_io_out; // @[RegFile.scala 66:20:@45067.4]
  wire  regs_239_io_enable; // @[RegFile.scala 66:20:@45067.4]
  wire  regs_240_clock; // @[RegFile.scala 66:20:@45081.4]
  wire  regs_240_reset; // @[RegFile.scala 66:20:@45081.4]
  wire [63:0] regs_240_io_in; // @[RegFile.scala 66:20:@45081.4]
  wire  regs_240_io_reset; // @[RegFile.scala 66:20:@45081.4]
  wire [63:0] regs_240_io_out; // @[RegFile.scala 66:20:@45081.4]
  wire  regs_240_io_enable; // @[RegFile.scala 66:20:@45081.4]
  wire  regs_241_clock; // @[RegFile.scala 66:20:@45095.4]
  wire  regs_241_reset; // @[RegFile.scala 66:20:@45095.4]
  wire [63:0] regs_241_io_in; // @[RegFile.scala 66:20:@45095.4]
  wire  regs_241_io_reset; // @[RegFile.scala 66:20:@45095.4]
  wire [63:0] regs_241_io_out; // @[RegFile.scala 66:20:@45095.4]
  wire  regs_241_io_enable; // @[RegFile.scala 66:20:@45095.4]
  wire  regs_242_clock; // @[RegFile.scala 66:20:@45109.4]
  wire  regs_242_reset; // @[RegFile.scala 66:20:@45109.4]
  wire [63:0] regs_242_io_in; // @[RegFile.scala 66:20:@45109.4]
  wire  regs_242_io_reset; // @[RegFile.scala 66:20:@45109.4]
  wire [63:0] regs_242_io_out; // @[RegFile.scala 66:20:@45109.4]
  wire  regs_242_io_enable; // @[RegFile.scala 66:20:@45109.4]
  wire  regs_243_clock; // @[RegFile.scala 66:20:@45123.4]
  wire  regs_243_reset; // @[RegFile.scala 66:20:@45123.4]
  wire [63:0] regs_243_io_in; // @[RegFile.scala 66:20:@45123.4]
  wire  regs_243_io_reset; // @[RegFile.scala 66:20:@45123.4]
  wire [63:0] regs_243_io_out; // @[RegFile.scala 66:20:@45123.4]
  wire  regs_243_io_enable; // @[RegFile.scala 66:20:@45123.4]
  wire  regs_244_clock; // @[RegFile.scala 66:20:@45137.4]
  wire  regs_244_reset; // @[RegFile.scala 66:20:@45137.4]
  wire [63:0] regs_244_io_in; // @[RegFile.scala 66:20:@45137.4]
  wire  regs_244_io_reset; // @[RegFile.scala 66:20:@45137.4]
  wire [63:0] regs_244_io_out; // @[RegFile.scala 66:20:@45137.4]
  wire  regs_244_io_enable; // @[RegFile.scala 66:20:@45137.4]
  wire  regs_245_clock; // @[RegFile.scala 66:20:@45151.4]
  wire  regs_245_reset; // @[RegFile.scala 66:20:@45151.4]
  wire [63:0] regs_245_io_in; // @[RegFile.scala 66:20:@45151.4]
  wire  regs_245_io_reset; // @[RegFile.scala 66:20:@45151.4]
  wire [63:0] regs_245_io_out; // @[RegFile.scala 66:20:@45151.4]
  wire  regs_245_io_enable; // @[RegFile.scala 66:20:@45151.4]
  wire  regs_246_clock; // @[RegFile.scala 66:20:@45165.4]
  wire  regs_246_reset; // @[RegFile.scala 66:20:@45165.4]
  wire [63:0] regs_246_io_in; // @[RegFile.scala 66:20:@45165.4]
  wire  regs_246_io_reset; // @[RegFile.scala 66:20:@45165.4]
  wire [63:0] regs_246_io_out; // @[RegFile.scala 66:20:@45165.4]
  wire  regs_246_io_enable; // @[RegFile.scala 66:20:@45165.4]
  wire  regs_247_clock; // @[RegFile.scala 66:20:@45179.4]
  wire  regs_247_reset; // @[RegFile.scala 66:20:@45179.4]
  wire [63:0] regs_247_io_in; // @[RegFile.scala 66:20:@45179.4]
  wire  regs_247_io_reset; // @[RegFile.scala 66:20:@45179.4]
  wire [63:0] regs_247_io_out; // @[RegFile.scala 66:20:@45179.4]
  wire  regs_247_io_enable; // @[RegFile.scala 66:20:@45179.4]
  wire  regs_248_clock; // @[RegFile.scala 66:20:@45193.4]
  wire  regs_248_reset; // @[RegFile.scala 66:20:@45193.4]
  wire [63:0] regs_248_io_in; // @[RegFile.scala 66:20:@45193.4]
  wire  regs_248_io_reset; // @[RegFile.scala 66:20:@45193.4]
  wire [63:0] regs_248_io_out; // @[RegFile.scala 66:20:@45193.4]
  wire  regs_248_io_enable; // @[RegFile.scala 66:20:@45193.4]
  wire  regs_249_clock; // @[RegFile.scala 66:20:@45207.4]
  wire  regs_249_reset; // @[RegFile.scala 66:20:@45207.4]
  wire [63:0] regs_249_io_in; // @[RegFile.scala 66:20:@45207.4]
  wire  regs_249_io_reset; // @[RegFile.scala 66:20:@45207.4]
  wire [63:0] regs_249_io_out; // @[RegFile.scala 66:20:@45207.4]
  wire  regs_249_io_enable; // @[RegFile.scala 66:20:@45207.4]
  wire  regs_250_clock; // @[RegFile.scala 66:20:@45221.4]
  wire  regs_250_reset; // @[RegFile.scala 66:20:@45221.4]
  wire [63:0] regs_250_io_in; // @[RegFile.scala 66:20:@45221.4]
  wire  regs_250_io_reset; // @[RegFile.scala 66:20:@45221.4]
  wire [63:0] regs_250_io_out; // @[RegFile.scala 66:20:@45221.4]
  wire  regs_250_io_enable; // @[RegFile.scala 66:20:@45221.4]
  wire  regs_251_clock; // @[RegFile.scala 66:20:@45235.4]
  wire  regs_251_reset; // @[RegFile.scala 66:20:@45235.4]
  wire [63:0] regs_251_io_in; // @[RegFile.scala 66:20:@45235.4]
  wire  regs_251_io_reset; // @[RegFile.scala 66:20:@45235.4]
  wire [63:0] regs_251_io_out; // @[RegFile.scala 66:20:@45235.4]
  wire  regs_251_io_enable; // @[RegFile.scala 66:20:@45235.4]
  wire  regs_252_clock; // @[RegFile.scala 66:20:@45249.4]
  wire  regs_252_reset; // @[RegFile.scala 66:20:@45249.4]
  wire [63:0] regs_252_io_in; // @[RegFile.scala 66:20:@45249.4]
  wire  regs_252_io_reset; // @[RegFile.scala 66:20:@45249.4]
  wire [63:0] regs_252_io_out; // @[RegFile.scala 66:20:@45249.4]
  wire  regs_252_io_enable; // @[RegFile.scala 66:20:@45249.4]
  wire  regs_253_clock; // @[RegFile.scala 66:20:@45263.4]
  wire  regs_253_reset; // @[RegFile.scala 66:20:@45263.4]
  wire [63:0] regs_253_io_in; // @[RegFile.scala 66:20:@45263.4]
  wire  regs_253_io_reset; // @[RegFile.scala 66:20:@45263.4]
  wire [63:0] regs_253_io_out; // @[RegFile.scala 66:20:@45263.4]
  wire  regs_253_io_enable; // @[RegFile.scala 66:20:@45263.4]
  wire  regs_254_clock; // @[RegFile.scala 66:20:@45277.4]
  wire  regs_254_reset; // @[RegFile.scala 66:20:@45277.4]
  wire [63:0] regs_254_io_in; // @[RegFile.scala 66:20:@45277.4]
  wire  regs_254_io_reset; // @[RegFile.scala 66:20:@45277.4]
  wire [63:0] regs_254_io_out; // @[RegFile.scala 66:20:@45277.4]
  wire  regs_254_io_enable; // @[RegFile.scala 66:20:@45277.4]
  wire  regs_255_clock; // @[RegFile.scala 66:20:@45291.4]
  wire  regs_255_reset; // @[RegFile.scala 66:20:@45291.4]
  wire [63:0] regs_255_io_in; // @[RegFile.scala 66:20:@45291.4]
  wire  regs_255_io_reset; // @[RegFile.scala 66:20:@45291.4]
  wire [63:0] regs_255_io_out; // @[RegFile.scala 66:20:@45291.4]
  wire  regs_255_io_enable; // @[RegFile.scala 66:20:@45291.4]
  wire  regs_256_clock; // @[RegFile.scala 66:20:@45305.4]
  wire  regs_256_reset; // @[RegFile.scala 66:20:@45305.4]
  wire [63:0] regs_256_io_in; // @[RegFile.scala 66:20:@45305.4]
  wire  regs_256_io_reset; // @[RegFile.scala 66:20:@45305.4]
  wire [63:0] regs_256_io_out; // @[RegFile.scala 66:20:@45305.4]
  wire  regs_256_io_enable; // @[RegFile.scala 66:20:@45305.4]
  wire  regs_257_clock; // @[RegFile.scala 66:20:@45319.4]
  wire  regs_257_reset; // @[RegFile.scala 66:20:@45319.4]
  wire [63:0] regs_257_io_in; // @[RegFile.scala 66:20:@45319.4]
  wire  regs_257_io_reset; // @[RegFile.scala 66:20:@45319.4]
  wire [63:0] regs_257_io_out; // @[RegFile.scala 66:20:@45319.4]
  wire  regs_257_io_enable; // @[RegFile.scala 66:20:@45319.4]
  wire  regs_258_clock; // @[RegFile.scala 66:20:@45333.4]
  wire  regs_258_reset; // @[RegFile.scala 66:20:@45333.4]
  wire [63:0] regs_258_io_in; // @[RegFile.scala 66:20:@45333.4]
  wire  regs_258_io_reset; // @[RegFile.scala 66:20:@45333.4]
  wire [63:0] regs_258_io_out; // @[RegFile.scala 66:20:@45333.4]
  wire  regs_258_io_enable; // @[RegFile.scala 66:20:@45333.4]
  wire  regs_259_clock; // @[RegFile.scala 66:20:@45347.4]
  wire  regs_259_reset; // @[RegFile.scala 66:20:@45347.4]
  wire [63:0] regs_259_io_in; // @[RegFile.scala 66:20:@45347.4]
  wire  regs_259_io_reset; // @[RegFile.scala 66:20:@45347.4]
  wire [63:0] regs_259_io_out; // @[RegFile.scala 66:20:@45347.4]
  wire  regs_259_io_enable; // @[RegFile.scala 66:20:@45347.4]
  wire  regs_260_clock; // @[RegFile.scala 66:20:@45361.4]
  wire  regs_260_reset; // @[RegFile.scala 66:20:@45361.4]
  wire [63:0] regs_260_io_in; // @[RegFile.scala 66:20:@45361.4]
  wire  regs_260_io_reset; // @[RegFile.scala 66:20:@45361.4]
  wire [63:0] regs_260_io_out; // @[RegFile.scala 66:20:@45361.4]
  wire  regs_260_io_enable; // @[RegFile.scala 66:20:@45361.4]
  wire  regs_261_clock; // @[RegFile.scala 66:20:@45375.4]
  wire  regs_261_reset; // @[RegFile.scala 66:20:@45375.4]
  wire [63:0] regs_261_io_in; // @[RegFile.scala 66:20:@45375.4]
  wire  regs_261_io_reset; // @[RegFile.scala 66:20:@45375.4]
  wire [63:0] regs_261_io_out; // @[RegFile.scala 66:20:@45375.4]
  wire  regs_261_io_enable; // @[RegFile.scala 66:20:@45375.4]
  wire  regs_262_clock; // @[RegFile.scala 66:20:@45389.4]
  wire  regs_262_reset; // @[RegFile.scala 66:20:@45389.4]
  wire [63:0] regs_262_io_in; // @[RegFile.scala 66:20:@45389.4]
  wire  regs_262_io_reset; // @[RegFile.scala 66:20:@45389.4]
  wire [63:0] regs_262_io_out; // @[RegFile.scala 66:20:@45389.4]
  wire  regs_262_io_enable; // @[RegFile.scala 66:20:@45389.4]
  wire  regs_263_clock; // @[RegFile.scala 66:20:@45403.4]
  wire  regs_263_reset; // @[RegFile.scala 66:20:@45403.4]
  wire [63:0] regs_263_io_in; // @[RegFile.scala 66:20:@45403.4]
  wire  regs_263_io_reset; // @[RegFile.scala 66:20:@45403.4]
  wire [63:0] regs_263_io_out; // @[RegFile.scala 66:20:@45403.4]
  wire  regs_263_io_enable; // @[RegFile.scala 66:20:@45403.4]
  wire  regs_264_clock; // @[RegFile.scala 66:20:@45417.4]
  wire  regs_264_reset; // @[RegFile.scala 66:20:@45417.4]
  wire [63:0] regs_264_io_in; // @[RegFile.scala 66:20:@45417.4]
  wire  regs_264_io_reset; // @[RegFile.scala 66:20:@45417.4]
  wire [63:0] regs_264_io_out; // @[RegFile.scala 66:20:@45417.4]
  wire  regs_264_io_enable; // @[RegFile.scala 66:20:@45417.4]
  wire  regs_265_clock; // @[RegFile.scala 66:20:@45431.4]
  wire  regs_265_reset; // @[RegFile.scala 66:20:@45431.4]
  wire [63:0] regs_265_io_in; // @[RegFile.scala 66:20:@45431.4]
  wire  regs_265_io_reset; // @[RegFile.scala 66:20:@45431.4]
  wire [63:0] regs_265_io_out; // @[RegFile.scala 66:20:@45431.4]
  wire  regs_265_io_enable; // @[RegFile.scala 66:20:@45431.4]
  wire  regs_266_clock; // @[RegFile.scala 66:20:@45445.4]
  wire  regs_266_reset; // @[RegFile.scala 66:20:@45445.4]
  wire [63:0] regs_266_io_in; // @[RegFile.scala 66:20:@45445.4]
  wire  regs_266_io_reset; // @[RegFile.scala 66:20:@45445.4]
  wire [63:0] regs_266_io_out; // @[RegFile.scala 66:20:@45445.4]
  wire  regs_266_io_enable; // @[RegFile.scala 66:20:@45445.4]
  wire  regs_267_clock; // @[RegFile.scala 66:20:@45459.4]
  wire  regs_267_reset; // @[RegFile.scala 66:20:@45459.4]
  wire [63:0] regs_267_io_in; // @[RegFile.scala 66:20:@45459.4]
  wire  regs_267_io_reset; // @[RegFile.scala 66:20:@45459.4]
  wire [63:0] regs_267_io_out; // @[RegFile.scala 66:20:@45459.4]
  wire  regs_267_io_enable; // @[RegFile.scala 66:20:@45459.4]
  wire  regs_268_clock; // @[RegFile.scala 66:20:@45473.4]
  wire  regs_268_reset; // @[RegFile.scala 66:20:@45473.4]
  wire [63:0] regs_268_io_in; // @[RegFile.scala 66:20:@45473.4]
  wire  regs_268_io_reset; // @[RegFile.scala 66:20:@45473.4]
  wire [63:0] regs_268_io_out; // @[RegFile.scala 66:20:@45473.4]
  wire  regs_268_io_enable; // @[RegFile.scala 66:20:@45473.4]
  wire  regs_269_clock; // @[RegFile.scala 66:20:@45487.4]
  wire  regs_269_reset; // @[RegFile.scala 66:20:@45487.4]
  wire [63:0] regs_269_io_in; // @[RegFile.scala 66:20:@45487.4]
  wire  regs_269_io_reset; // @[RegFile.scala 66:20:@45487.4]
  wire [63:0] regs_269_io_out; // @[RegFile.scala 66:20:@45487.4]
  wire  regs_269_io_enable; // @[RegFile.scala 66:20:@45487.4]
  wire  regs_270_clock; // @[RegFile.scala 66:20:@45501.4]
  wire  regs_270_reset; // @[RegFile.scala 66:20:@45501.4]
  wire [63:0] regs_270_io_in; // @[RegFile.scala 66:20:@45501.4]
  wire  regs_270_io_reset; // @[RegFile.scala 66:20:@45501.4]
  wire [63:0] regs_270_io_out; // @[RegFile.scala 66:20:@45501.4]
  wire  regs_270_io_enable; // @[RegFile.scala 66:20:@45501.4]
  wire  regs_271_clock; // @[RegFile.scala 66:20:@45515.4]
  wire  regs_271_reset; // @[RegFile.scala 66:20:@45515.4]
  wire [63:0] regs_271_io_in; // @[RegFile.scala 66:20:@45515.4]
  wire  regs_271_io_reset; // @[RegFile.scala 66:20:@45515.4]
  wire [63:0] regs_271_io_out; // @[RegFile.scala 66:20:@45515.4]
  wire  regs_271_io_enable; // @[RegFile.scala 66:20:@45515.4]
  wire  regs_272_clock; // @[RegFile.scala 66:20:@45529.4]
  wire  regs_272_reset; // @[RegFile.scala 66:20:@45529.4]
  wire [63:0] regs_272_io_in; // @[RegFile.scala 66:20:@45529.4]
  wire  regs_272_io_reset; // @[RegFile.scala 66:20:@45529.4]
  wire [63:0] regs_272_io_out; // @[RegFile.scala 66:20:@45529.4]
  wire  regs_272_io_enable; // @[RegFile.scala 66:20:@45529.4]
  wire  regs_273_clock; // @[RegFile.scala 66:20:@45543.4]
  wire  regs_273_reset; // @[RegFile.scala 66:20:@45543.4]
  wire [63:0] regs_273_io_in; // @[RegFile.scala 66:20:@45543.4]
  wire  regs_273_io_reset; // @[RegFile.scala 66:20:@45543.4]
  wire [63:0] regs_273_io_out; // @[RegFile.scala 66:20:@45543.4]
  wire  regs_273_io_enable; // @[RegFile.scala 66:20:@45543.4]
  wire  regs_274_clock; // @[RegFile.scala 66:20:@45557.4]
  wire  regs_274_reset; // @[RegFile.scala 66:20:@45557.4]
  wire [63:0] regs_274_io_in; // @[RegFile.scala 66:20:@45557.4]
  wire  regs_274_io_reset; // @[RegFile.scala 66:20:@45557.4]
  wire [63:0] regs_274_io_out; // @[RegFile.scala 66:20:@45557.4]
  wire  regs_274_io_enable; // @[RegFile.scala 66:20:@45557.4]
  wire  regs_275_clock; // @[RegFile.scala 66:20:@45571.4]
  wire  regs_275_reset; // @[RegFile.scala 66:20:@45571.4]
  wire [63:0] regs_275_io_in; // @[RegFile.scala 66:20:@45571.4]
  wire  regs_275_io_reset; // @[RegFile.scala 66:20:@45571.4]
  wire [63:0] regs_275_io_out; // @[RegFile.scala 66:20:@45571.4]
  wire  regs_275_io_enable; // @[RegFile.scala 66:20:@45571.4]
  wire  regs_276_clock; // @[RegFile.scala 66:20:@45585.4]
  wire  regs_276_reset; // @[RegFile.scala 66:20:@45585.4]
  wire [63:0] regs_276_io_in; // @[RegFile.scala 66:20:@45585.4]
  wire  regs_276_io_reset; // @[RegFile.scala 66:20:@45585.4]
  wire [63:0] regs_276_io_out; // @[RegFile.scala 66:20:@45585.4]
  wire  regs_276_io_enable; // @[RegFile.scala 66:20:@45585.4]
  wire  regs_277_clock; // @[RegFile.scala 66:20:@45599.4]
  wire  regs_277_reset; // @[RegFile.scala 66:20:@45599.4]
  wire [63:0] regs_277_io_in; // @[RegFile.scala 66:20:@45599.4]
  wire  regs_277_io_reset; // @[RegFile.scala 66:20:@45599.4]
  wire [63:0] regs_277_io_out; // @[RegFile.scala 66:20:@45599.4]
  wire  regs_277_io_enable; // @[RegFile.scala 66:20:@45599.4]
  wire  regs_278_clock; // @[RegFile.scala 66:20:@45613.4]
  wire  regs_278_reset; // @[RegFile.scala 66:20:@45613.4]
  wire [63:0] regs_278_io_in; // @[RegFile.scala 66:20:@45613.4]
  wire  regs_278_io_reset; // @[RegFile.scala 66:20:@45613.4]
  wire [63:0] regs_278_io_out; // @[RegFile.scala 66:20:@45613.4]
  wire  regs_278_io_enable; // @[RegFile.scala 66:20:@45613.4]
  wire  regs_279_clock; // @[RegFile.scala 66:20:@45627.4]
  wire  regs_279_reset; // @[RegFile.scala 66:20:@45627.4]
  wire [63:0] regs_279_io_in; // @[RegFile.scala 66:20:@45627.4]
  wire  regs_279_io_reset; // @[RegFile.scala 66:20:@45627.4]
  wire [63:0] regs_279_io_out; // @[RegFile.scala 66:20:@45627.4]
  wire  regs_279_io_enable; // @[RegFile.scala 66:20:@45627.4]
  wire  regs_280_clock; // @[RegFile.scala 66:20:@45641.4]
  wire  regs_280_reset; // @[RegFile.scala 66:20:@45641.4]
  wire [63:0] regs_280_io_in; // @[RegFile.scala 66:20:@45641.4]
  wire  regs_280_io_reset; // @[RegFile.scala 66:20:@45641.4]
  wire [63:0] regs_280_io_out; // @[RegFile.scala 66:20:@45641.4]
  wire  regs_280_io_enable; // @[RegFile.scala 66:20:@45641.4]
  wire  regs_281_clock; // @[RegFile.scala 66:20:@45655.4]
  wire  regs_281_reset; // @[RegFile.scala 66:20:@45655.4]
  wire [63:0] regs_281_io_in; // @[RegFile.scala 66:20:@45655.4]
  wire  regs_281_io_reset; // @[RegFile.scala 66:20:@45655.4]
  wire [63:0] regs_281_io_out; // @[RegFile.scala 66:20:@45655.4]
  wire  regs_281_io_enable; // @[RegFile.scala 66:20:@45655.4]
  wire  regs_282_clock; // @[RegFile.scala 66:20:@45669.4]
  wire  regs_282_reset; // @[RegFile.scala 66:20:@45669.4]
  wire [63:0] regs_282_io_in; // @[RegFile.scala 66:20:@45669.4]
  wire  regs_282_io_reset; // @[RegFile.scala 66:20:@45669.4]
  wire [63:0] regs_282_io_out; // @[RegFile.scala 66:20:@45669.4]
  wire  regs_282_io_enable; // @[RegFile.scala 66:20:@45669.4]
  wire  regs_283_clock; // @[RegFile.scala 66:20:@45683.4]
  wire  regs_283_reset; // @[RegFile.scala 66:20:@45683.4]
  wire [63:0] regs_283_io_in; // @[RegFile.scala 66:20:@45683.4]
  wire  regs_283_io_reset; // @[RegFile.scala 66:20:@45683.4]
  wire [63:0] regs_283_io_out; // @[RegFile.scala 66:20:@45683.4]
  wire  regs_283_io_enable; // @[RegFile.scala 66:20:@45683.4]
  wire  regs_284_clock; // @[RegFile.scala 66:20:@45697.4]
  wire  regs_284_reset; // @[RegFile.scala 66:20:@45697.4]
  wire [63:0] regs_284_io_in; // @[RegFile.scala 66:20:@45697.4]
  wire  regs_284_io_reset; // @[RegFile.scala 66:20:@45697.4]
  wire [63:0] regs_284_io_out; // @[RegFile.scala 66:20:@45697.4]
  wire  regs_284_io_enable; // @[RegFile.scala 66:20:@45697.4]
  wire  regs_285_clock; // @[RegFile.scala 66:20:@45711.4]
  wire  regs_285_reset; // @[RegFile.scala 66:20:@45711.4]
  wire [63:0] regs_285_io_in; // @[RegFile.scala 66:20:@45711.4]
  wire  regs_285_io_reset; // @[RegFile.scala 66:20:@45711.4]
  wire [63:0] regs_285_io_out; // @[RegFile.scala 66:20:@45711.4]
  wire  regs_285_io_enable; // @[RegFile.scala 66:20:@45711.4]
  wire  regs_286_clock; // @[RegFile.scala 66:20:@45725.4]
  wire  regs_286_reset; // @[RegFile.scala 66:20:@45725.4]
  wire [63:0] regs_286_io_in; // @[RegFile.scala 66:20:@45725.4]
  wire  regs_286_io_reset; // @[RegFile.scala 66:20:@45725.4]
  wire [63:0] regs_286_io_out; // @[RegFile.scala 66:20:@45725.4]
  wire  regs_286_io_enable; // @[RegFile.scala 66:20:@45725.4]
  wire  regs_287_clock; // @[RegFile.scala 66:20:@45739.4]
  wire  regs_287_reset; // @[RegFile.scala 66:20:@45739.4]
  wire [63:0] regs_287_io_in; // @[RegFile.scala 66:20:@45739.4]
  wire  regs_287_io_reset; // @[RegFile.scala 66:20:@45739.4]
  wire [63:0] regs_287_io_out; // @[RegFile.scala 66:20:@45739.4]
  wire  regs_287_io_enable; // @[RegFile.scala 66:20:@45739.4]
  wire  regs_288_clock; // @[RegFile.scala 66:20:@45753.4]
  wire  regs_288_reset; // @[RegFile.scala 66:20:@45753.4]
  wire [63:0] regs_288_io_in; // @[RegFile.scala 66:20:@45753.4]
  wire  regs_288_io_reset; // @[RegFile.scala 66:20:@45753.4]
  wire [63:0] regs_288_io_out; // @[RegFile.scala 66:20:@45753.4]
  wire  regs_288_io_enable; // @[RegFile.scala 66:20:@45753.4]
  wire  regs_289_clock; // @[RegFile.scala 66:20:@45767.4]
  wire  regs_289_reset; // @[RegFile.scala 66:20:@45767.4]
  wire [63:0] regs_289_io_in; // @[RegFile.scala 66:20:@45767.4]
  wire  regs_289_io_reset; // @[RegFile.scala 66:20:@45767.4]
  wire [63:0] regs_289_io_out; // @[RegFile.scala 66:20:@45767.4]
  wire  regs_289_io_enable; // @[RegFile.scala 66:20:@45767.4]
  wire  regs_290_clock; // @[RegFile.scala 66:20:@45781.4]
  wire  regs_290_reset; // @[RegFile.scala 66:20:@45781.4]
  wire [63:0] regs_290_io_in; // @[RegFile.scala 66:20:@45781.4]
  wire  regs_290_io_reset; // @[RegFile.scala 66:20:@45781.4]
  wire [63:0] regs_290_io_out; // @[RegFile.scala 66:20:@45781.4]
  wire  regs_290_io_enable; // @[RegFile.scala 66:20:@45781.4]
  wire  regs_291_clock; // @[RegFile.scala 66:20:@45795.4]
  wire  regs_291_reset; // @[RegFile.scala 66:20:@45795.4]
  wire [63:0] regs_291_io_in; // @[RegFile.scala 66:20:@45795.4]
  wire  regs_291_io_reset; // @[RegFile.scala 66:20:@45795.4]
  wire [63:0] regs_291_io_out; // @[RegFile.scala 66:20:@45795.4]
  wire  regs_291_io_enable; // @[RegFile.scala 66:20:@45795.4]
  wire  regs_292_clock; // @[RegFile.scala 66:20:@45809.4]
  wire  regs_292_reset; // @[RegFile.scala 66:20:@45809.4]
  wire [63:0] regs_292_io_in; // @[RegFile.scala 66:20:@45809.4]
  wire  regs_292_io_reset; // @[RegFile.scala 66:20:@45809.4]
  wire [63:0] regs_292_io_out; // @[RegFile.scala 66:20:@45809.4]
  wire  regs_292_io_enable; // @[RegFile.scala 66:20:@45809.4]
  wire  regs_293_clock; // @[RegFile.scala 66:20:@45823.4]
  wire  regs_293_reset; // @[RegFile.scala 66:20:@45823.4]
  wire [63:0] regs_293_io_in; // @[RegFile.scala 66:20:@45823.4]
  wire  regs_293_io_reset; // @[RegFile.scala 66:20:@45823.4]
  wire [63:0] regs_293_io_out; // @[RegFile.scala 66:20:@45823.4]
  wire  regs_293_io_enable; // @[RegFile.scala 66:20:@45823.4]
  wire  regs_294_clock; // @[RegFile.scala 66:20:@45837.4]
  wire  regs_294_reset; // @[RegFile.scala 66:20:@45837.4]
  wire [63:0] regs_294_io_in; // @[RegFile.scala 66:20:@45837.4]
  wire  regs_294_io_reset; // @[RegFile.scala 66:20:@45837.4]
  wire [63:0] regs_294_io_out; // @[RegFile.scala 66:20:@45837.4]
  wire  regs_294_io_enable; // @[RegFile.scala 66:20:@45837.4]
  wire  regs_295_clock; // @[RegFile.scala 66:20:@45851.4]
  wire  regs_295_reset; // @[RegFile.scala 66:20:@45851.4]
  wire [63:0] regs_295_io_in; // @[RegFile.scala 66:20:@45851.4]
  wire  regs_295_io_reset; // @[RegFile.scala 66:20:@45851.4]
  wire [63:0] regs_295_io_out; // @[RegFile.scala 66:20:@45851.4]
  wire  regs_295_io_enable; // @[RegFile.scala 66:20:@45851.4]
  wire  regs_296_clock; // @[RegFile.scala 66:20:@45865.4]
  wire  regs_296_reset; // @[RegFile.scala 66:20:@45865.4]
  wire [63:0] regs_296_io_in; // @[RegFile.scala 66:20:@45865.4]
  wire  regs_296_io_reset; // @[RegFile.scala 66:20:@45865.4]
  wire [63:0] regs_296_io_out; // @[RegFile.scala 66:20:@45865.4]
  wire  regs_296_io_enable; // @[RegFile.scala 66:20:@45865.4]
  wire  regs_297_clock; // @[RegFile.scala 66:20:@45879.4]
  wire  regs_297_reset; // @[RegFile.scala 66:20:@45879.4]
  wire [63:0] regs_297_io_in; // @[RegFile.scala 66:20:@45879.4]
  wire  regs_297_io_reset; // @[RegFile.scala 66:20:@45879.4]
  wire [63:0] regs_297_io_out; // @[RegFile.scala 66:20:@45879.4]
  wire  regs_297_io_enable; // @[RegFile.scala 66:20:@45879.4]
  wire  regs_298_clock; // @[RegFile.scala 66:20:@45893.4]
  wire  regs_298_reset; // @[RegFile.scala 66:20:@45893.4]
  wire [63:0] regs_298_io_in; // @[RegFile.scala 66:20:@45893.4]
  wire  regs_298_io_reset; // @[RegFile.scala 66:20:@45893.4]
  wire [63:0] regs_298_io_out; // @[RegFile.scala 66:20:@45893.4]
  wire  regs_298_io_enable; // @[RegFile.scala 66:20:@45893.4]
  wire  regs_299_clock; // @[RegFile.scala 66:20:@45907.4]
  wire  regs_299_reset; // @[RegFile.scala 66:20:@45907.4]
  wire [63:0] regs_299_io_in; // @[RegFile.scala 66:20:@45907.4]
  wire  regs_299_io_reset; // @[RegFile.scala 66:20:@45907.4]
  wire [63:0] regs_299_io_out; // @[RegFile.scala 66:20:@45907.4]
  wire  regs_299_io_enable; // @[RegFile.scala 66:20:@45907.4]
  wire  regs_300_clock; // @[RegFile.scala 66:20:@45921.4]
  wire  regs_300_reset; // @[RegFile.scala 66:20:@45921.4]
  wire [63:0] regs_300_io_in; // @[RegFile.scala 66:20:@45921.4]
  wire  regs_300_io_reset; // @[RegFile.scala 66:20:@45921.4]
  wire [63:0] regs_300_io_out; // @[RegFile.scala 66:20:@45921.4]
  wire  regs_300_io_enable; // @[RegFile.scala 66:20:@45921.4]
  wire  regs_301_clock; // @[RegFile.scala 66:20:@45935.4]
  wire  regs_301_reset; // @[RegFile.scala 66:20:@45935.4]
  wire [63:0] regs_301_io_in; // @[RegFile.scala 66:20:@45935.4]
  wire  regs_301_io_reset; // @[RegFile.scala 66:20:@45935.4]
  wire [63:0] regs_301_io_out; // @[RegFile.scala 66:20:@45935.4]
  wire  regs_301_io_enable; // @[RegFile.scala 66:20:@45935.4]
  wire  regs_302_clock; // @[RegFile.scala 66:20:@45949.4]
  wire  regs_302_reset; // @[RegFile.scala 66:20:@45949.4]
  wire [63:0] regs_302_io_in; // @[RegFile.scala 66:20:@45949.4]
  wire  regs_302_io_reset; // @[RegFile.scala 66:20:@45949.4]
  wire [63:0] regs_302_io_out; // @[RegFile.scala 66:20:@45949.4]
  wire  regs_302_io_enable; // @[RegFile.scala 66:20:@45949.4]
  wire  regs_303_clock; // @[RegFile.scala 66:20:@45963.4]
  wire  regs_303_reset; // @[RegFile.scala 66:20:@45963.4]
  wire [63:0] regs_303_io_in; // @[RegFile.scala 66:20:@45963.4]
  wire  regs_303_io_reset; // @[RegFile.scala 66:20:@45963.4]
  wire [63:0] regs_303_io_out; // @[RegFile.scala 66:20:@45963.4]
  wire  regs_303_io_enable; // @[RegFile.scala 66:20:@45963.4]
  wire  regs_304_clock; // @[RegFile.scala 66:20:@45977.4]
  wire  regs_304_reset; // @[RegFile.scala 66:20:@45977.4]
  wire [63:0] regs_304_io_in; // @[RegFile.scala 66:20:@45977.4]
  wire  regs_304_io_reset; // @[RegFile.scala 66:20:@45977.4]
  wire [63:0] regs_304_io_out; // @[RegFile.scala 66:20:@45977.4]
  wire  regs_304_io_enable; // @[RegFile.scala 66:20:@45977.4]
  wire  regs_305_clock; // @[RegFile.scala 66:20:@45991.4]
  wire  regs_305_reset; // @[RegFile.scala 66:20:@45991.4]
  wire [63:0] regs_305_io_in; // @[RegFile.scala 66:20:@45991.4]
  wire  regs_305_io_reset; // @[RegFile.scala 66:20:@45991.4]
  wire [63:0] regs_305_io_out; // @[RegFile.scala 66:20:@45991.4]
  wire  regs_305_io_enable; // @[RegFile.scala 66:20:@45991.4]
  wire  regs_306_clock; // @[RegFile.scala 66:20:@46005.4]
  wire  regs_306_reset; // @[RegFile.scala 66:20:@46005.4]
  wire [63:0] regs_306_io_in; // @[RegFile.scala 66:20:@46005.4]
  wire  regs_306_io_reset; // @[RegFile.scala 66:20:@46005.4]
  wire [63:0] regs_306_io_out; // @[RegFile.scala 66:20:@46005.4]
  wire  regs_306_io_enable; // @[RegFile.scala 66:20:@46005.4]
  wire  regs_307_clock; // @[RegFile.scala 66:20:@46019.4]
  wire  regs_307_reset; // @[RegFile.scala 66:20:@46019.4]
  wire [63:0] regs_307_io_in; // @[RegFile.scala 66:20:@46019.4]
  wire  regs_307_io_reset; // @[RegFile.scala 66:20:@46019.4]
  wire [63:0] regs_307_io_out; // @[RegFile.scala 66:20:@46019.4]
  wire  regs_307_io_enable; // @[RegFile.scala 66:20:@46019.4]
  wire  regs_308_clock; // @[RegFile.scala 66:20:@46033.4]
  wire  regs_308_reset; // @[RegFile.scala 66:20:@46033.4]
  wire [63:0] regs_308_io_in; // @[RegFile.scala 66:20:@46033.4]
  wire  regs_308_io_reset; // @[RegFile.scala 66:20:@46033.4]
  wire [63:0] regs_308_io_out; // @[RegFile.scala 66:20:@46033.4]
  wire  regs_308_io_enable; // @[RegFile.scala 66:20:@46033.4]
  wire  regs_309_clock; // @[RegFile.scala 66:20:@46047.4]
  wire  regs_309_reset; // @[RegFile.scala 66:20:@46047.4]
  wire [63:0] regs_309_io_in; // @[RegFile.scala 66:20:@46047.4]
  wire  regs_309_io_reset; // @[RegFile.scala 66:20:@46047.4]
  wire [63:0] regs_309_io_out; // @[RegFile.scala 66:20:@46047.4]
  wire  regs_309_io_enable; // @[RegFile.scala 66:20:@46047.4]
  wire  regs_310_clock; // @[RegFile.scala 66:20:@46061.4]
  wire  regs_310_reset; // @[RegFile.scala 66:20:@46061.4]
  wire [63:0] regs_310_io_in; // @[RegFile.scala 66:20:@46061.4]
  wire  regs_310_io_reset; // @[RegFile.scala 66:20:@46061.4]
  wire [63:0] regs_310_io_out; // @[RegFile.scala 66:20:@46061.4]
  wire  regs_310_io_enable; // @[RegFile.scala 66:20:@46061.4]
  wire  regs_311_clock; // @[RegFile.scala 66:20:@46075.4]
  wire  regs_311_reset; // @[RegFile.scala 66:20:@46075.4]
  wire [63:0] regs_311_io_in; // @[RegFile.scala 66:20:@46075.4]
  wire  regs_311_io_reset; // @[RegFile.scala 66:20:@46075.4]
  wire [63:0] regs_311_io_out; // @[RegFile.scala 66:20:@46075.4]
  wire  regs_311_io_enable; // @[RegFile.scala 66:20:@46075.4]
  wire  regs_312_clock; // @[RegFile.scala 66:20:@46089.4]
  wire  regs_312_reset; // @[RegFile.scala 66:20:@46089.4]
  wire [63:0] regs_312_io_in; // @[RegFile.scala 66:20:@46089.4]
  wire  regs_312_io_reset; // @[RegFile.scala 66:20:@46089.4]
  wire [63:0] regs_312_io_out; // @[RegFile.scala 66:20:@46089.4]
  wire  regs_312_io_enable; // @[RegFile.scala 66:20:@46089.4]
  wire  regs_313_clock; // @[RegFile.scala 66:20:@46103.4]
  wire  regs_313_reset; // @[RegFile.scala 66:20:@46103.4]
  wire [63:0] regs_313_io_in; // @[RegFile.scala 66:20:@46103.4]
  wire  regs_313_io_reset; // @[RegFile.scala 66:20:@46103.4]
  wire [63:0] regs_313_io_out; // @[RegFile.scala 66:20:@46103.4]
  wire  regs_313_io_enable; // @[RegFile.scala 66:20:@46103.4]
  wire  regs_314_clock; // @[RegFile.scala 66:20:@46117.4]
  wire  regs_314_reset; // @[RegFile.scala 66:20:@46117.4]
  wire [63:0] regs_314_io_in; // @[RegFile.scala 66:20:@46117.4]
  wire  regs_314_io_reset; // @[RegFile.scala 66:20:@46117.4]
  wire [63:0] regs_314_io_out; // @[RegFile.scala 66:20:@46117.4]
  wire  regs_314_io_enable; // @[RegFile.scala 66:20:@46117.4]
  wire  regs_315_clock; // @[RegFile.scala 66:20:@46131.4]
  wire  regs_315_reset; // @[RegFile.scala 66:20:@46131.4]
  wire [63:0] regs_315_io_in; // @[RegFile.scala 66:20:@46131.4]
  wire  regs_315_io_reset; // @[RegFile.scala 66:20:@46131.4]
  wire [63:0] regs_315_io_out; // @[RegFile.scala 66:20:@46131.4]
  wire  regs_315_io_enable; // @[RegFile.scala 66:20:@46131.4]
  wire  regs_316_clock; // @[RegFile.scala 66:20:@46145.4]
  wire  regs_316_reset; // @[RegFile.scala 66:20:@46145.4]
  wire [63:0] regs_316_io_in; // @[RegFile.scala 66:20:@46145.4]
  wire  regs_316_io_reset; // @[RegFile.scala 66:20:@46145.4]
  wire [63:0] regs_316_io_out; // @[RegFile.scala 66:20:@46145.4]
  wire  regs_316_io_enable; // @[RegFile.scala 66:20:@46145.4]
  wire  regs_317_clock; // @[RegFile.scala 66:20:@46159.4]
  wire  regs_317_reset; // @[RegFile.scala 66:20:@46159.4]
  wire [63:0] regs_317_io_in; // @[RegFile.scala 66:20:@46159.4]
  wire  regs_317_io_reset; // @[RegFile.scala 66:20:@46159.4]
  wire [63:0] regs_317_io_out; // @[RegFile.scala 66:20:@46159.4]
  wire  regs_317_io_enable; // @[RegFile.scala 66:20:@46159.4]
  wire  regs_318_clock; // @[RegFile.scala 66:20:@46173.4]
  wire  regs_318_reset; // @[RegFile.scala 66:20:@46173.4]
  wire [63:0] regs_318_io_in; // @[RegFile.scala 66:20:@46173.4]
  wire  regs_318_io_reset; // @[RegFile.scala 66:20:@46173.4]
  wire [63:0] regs_318_io_out; // @[RegFile.scala 66:20:@46173.4]
  wire  regs_318_io_enable; // @[RegFile.scala 66:20:@46173.4]
  wire  regs_319_clock; // @[RegFile.scala 66:20:@46187.4]
  wire  regs_319_reset; // @[RegFile.scala 66:20:@46187.4]
  wire [63:0] regs_319_io_in; // @[RegFile.scala 66:20:@46187.4]
  wire  regs_319_io_reset; // @[RegFile.scala 66:20:@46187.4]
  wire [63:0] regs_319_io_out; // @[RegFile.scala 66:20:@46187.4]
  wire  regs_319_io_enable; // @[RegFile.scala 66:20:@46187.4]
  wire  regs_320_clock; // @[RegFile.scala 66:20:@46201.4]
  wire  regs_320_reset; // @[RegFile.scala 66:20:@46201.4]
  wire [63:0] regs_320_io_in; // @[RegFile.scala 66:20:@46201.4]
  wire  regs_320_io_reset; // @[RegFile.scala 66:20:@46201.4]
  wire [63:0] regs_320_io_out; // @[RegFile.scala 66:20:@46201.4]
  wire  regs_320_io_enable; // @[RegFile.scala 66:20:@46201.4]
  wire  regs_321_clock; // @[RegFile.scala 66:20:@46215.4]
  wire  regs_321_reset; // @[RegFile.scala 66:20:@46215.4]
  wire [63:0] regs_321_io_in; // @[RegFile.scala 66:20:@46215.4]
  wire  regs_321_io_reset; // @[RegFile.scala 66:20:@46215.4]
  wire [63:0] regs_321_io_out; // @[RegFile.scala 66:20:@46215.4]
  wire  regs_321_io_enable; // @[RegFile.scala 66:20:@46215.4]
  wire  regs_322_clock; // @[RegFile.scala 66:20:@46229.4]
  wire  regs_322_reset; // @[RegFile.scala 66:20:@46229.4]
  wire [63:0] regs_322_io_in; // @[RegFile.scala 66:20:@46229.4]
  wire  regs_322_io_reset; // @[RegFile.scala 66:20:@46229.4]
  wire [63:0] regs_322_io_out; // @[RegFile.scala 66:20:@46229.4]
  wire  regs_322_io_enable; // @[RegFile.scala 66:20:@46229.4]
  wire  regs_323_clock; // @[RegFile.scala 66:20:@46243.4]
  wire  regs_323_reset; // @[RegFile.scala 66:20:@46243.4]
  wire [63:0] regs_323_io_in; // @[RegFile.scala 66:20:@46243.4]
  wire  regs_323_io_reset; // @[RegFile.scala 66:20:@46243.4]
  wire [63:0] regs_323_io_out; // @[RegFile.scala 66:20:@46243.4]
  wire  regs_323_io_enable; // @[RegFile.scala 66:20:@46243.4]
  wire  regs_324_clock; // @[RegFile.scala 66:20:@46257.4]
  wire  regs_324_reset; // @[RegFile.scala 66:20:@46257.4]
  wire [63:0] regs_324_io_in; // @[RegFile.scala 66:20:@46257.4]
  wire  regs_324_io_reset; // @[RegFile.scala 66:20:@46257.4]
  wire [63:0] regs_324_io_out; // @[RegFile.scala 66:20:@46257.4]
  wire  regs_324_io_enable; // @[RegFile.scala 66:20:@46257.4]
  wire  regs_325_clock; // @[RegFile.scala 66:20:@46271.4]
  wire  regs_325_reset; // @[RegFile.scala 66:20:@46271.4]
  wire [63:0] regs_325_io_in; // @[RegFile.scala 66:20:@46271.4]
  wire  regs_325_io_reset; // @[RegFile.scala 66:20:@46271.4]
  wire [63:0] regs_325_io_out; // @[RegFile.scala 66:20:@46271.4]
  wire  regs_325_io_enable; // @[RegFile.scala 66:20:@46271.4]
  wire  regs_326_clock; // @[RegFile.scala 66:20:@46285.4]
  wire  regs_326_reset; // @[RegFile.scala 66:20:@46285.4]
  wire [63:0] regs_326_io_in; // @[RegFile.scala 66:20:@46285.4]
  wire  regs_326_io_reset; // @[RegFile.scala 66:20:@46285.4]
  wire [63:0] regs_326_io_out; // @[RegFile.scala 66:20:@46285.4]
  wire  regs_326_io_enable; // @[RegFile.scala 66:20:@46285.4]
  wire  regs_327_clock; // @[RegFile.scala 66:20:@46299.4]
  wire  regs_327_reset; // @[RegFile.scala 66:20:@46299.4]
  wire [63:0] regs_327_io_in; // @[RegFile.scala 66:20:@46299.4]
  wire  regs_327_io_reset; // @[RegFile.scala 66:20:@46299.4]
  wire [63:0] regs_327_io_out; // @[RegFile.scala 66:20:@46299.4]
  wire  regs_327_io_enable; // @[RegFile.scala 66:20:@46299.4]
  wire  regs_328_clock; // @[RegFile.scala 66:20:@46313.4]
  wire  regs_328_reset; // @[RegFile.scala 66:20:@46313.4]
  wire [63:0] regs_328_io_in; // @[RegFile.scala 66:20:@46313.4]
  wire  regs_328_io_reset; // @[RegFile.scala 66:20:@46313.4]
  wire [63:0] regs_328_io_out; // @[RegFile.scala 66:20:@46313.4]
  wire  regs_328_io_enable; // @[RegFile.scala 66:20:@46313.4]
  wire  regs_329_clock; // @[RegFile.scala 66:20:@46327.4]
  wire  regs_329_reset; // @[RegFile.scala 66:20:@46327.4]
  wire [63:0] regs_329_io_in; // @[RegFile.scala 66:20:@46327.4]
  wire  regs_329_io_reset; // @[RegFile.scala 66:20:@46327.4]
  wire [63:0] regs_329_io_out; // @[RegFile.scala 66:20:@46327.4]
  wire  regs_329_io_enable; // @[RegFile.scala 66:20:@46327.4]
  wire  regs_330_clock; // @[RegFile.scala 66:20:@46341.4]
  wire  regs_330_reset; // @[RegFile.scala 66:20:@46341.4]
  wire [63:0] regs_330_io_in; // @[RegFile.scala 66:20:@46341.4]
  wire  regs_330_io_reset; // @[RegFile.scala 66:20:@46341.4]
  wire [63:0] regs_330_io_out; // @[RegFile.scala 66:20:@46341.4]
  wire  regs_330_io_enable; // @[RegFile.scala 66:20:@46341.4]
  wire  regs_331_clock; // @[RegFile.scala 66:20:@46355.4]
  wire  regs_331_reset; // @[RegFile.scala 66:20:@46355.4]
  wire [63:0] regs_331_io_in; // @[RegFile.scala 66:20:@46355.4]
  wire  regs_331_io_reset; // @[RegFile.scala 66:20:@46355.4]
  wire [63:0] regs_331_io_out; // @[RegFile.scala 66:20:@46355.4]
  wire  regs_331_io_enable; // @[RegFile.scala 66:20:@46355.4]
  wire  regs_332_clock; // @[RegFile.scala 66:20:@46369.4]
  wire  regs_332_reset; // @[RegFile.scala 66:20:@46369.4]
  wire [63:0] regs_332_io_in; // @[RegFile.scala 66:20:@46369.4]
  wire  regs_332_io_reset; // @[RegFile.scala 66:20:@46369.4]
  wire [63:0] regs_332_io_out; // @[RegFile.scala 66:20:@46369.4]
  wire  regs_332_io_enable; // @[RegFile.scala 66:20:@46369.4]
  wire  regs_333_clock; // @[RegFile.scala 66:20:@46383.4]
  wire  regs_333_reset; // @[RegFile.scala 66:20:@46383.4]
  wire [63:0] regs_333_io_in; // @[RegFile.scala 66:20:@46383.4]
  wire  regs_333_io_reset; // @[RegFile.scala 66:20:@46383.4]
  wire [63:0] regs_333_io_out; // @[RegFile.scala 66:20:@46383.4]
  wire  regs_333_io_enable; // @[RegFile.scala 66:20:@46383.4]
  wire  regs_334_clock; // @[RegFile.scala 66:20:@46397.4]
  wire  regs_334_reset; // @[RegFile.scala 66:20:@46397.4]
  wire [63:0] regs_334_io_in; // @[RegFile.scala 66:20:@46397.4]
  wire  regs_334_io_reset; // @[RegFile.scala 66:20:@46397.4]
  wire [63:0] regs_334_io_out; // @[RegFile.scala 66:20:@46397.4]
  wire  regs_334_io_enable; // @[RegFile.scala 66:20:@46397.4]
  wire  regs_335_clock; // @[RegFile.scala 66:20:@46411.4]
  wire  regs_335_reset; // @[RegFile.scala 66:20:@46411.4]
  wire [63:0] regs_335_io_in; // @[RegFile.scala 66:20:@46411.4]
  wire  regs_335_io_reset; // @[RegFile.scala 66:20:@46411.4]
  wire [63:0] regs_335_io_out; // @[RegFile.scala 66:20:@46411.4]
  wire  regs_335_io_enable; // @[RegFile.scala 66:20:@46411.4]
  wire  regs_336_clock; // @[RegFile.scala 66:20:@46425.4]
  wire  regs_336_reset; // @[RegFile.scala 66:20:@46425.4]
  wire [63:0] regs_336_io_in; // @[RegFile.scala 66:20:@46425.4]
  wire  regs_336_io_reset; // @[RegFile.scala 66:20:@46425.4]
  wire [63:0] regs_336_io_out; // @[RegFile.scala 66:20:@46425.4]
  wire  regs_336_io_enable; // @[RegFile.scala 66:20:@46425.4]
  wire  regs_337_clock; // @[RegFile.scala 66:20:@46439.4]
  wire  regs_337_reset; // @[RegFile.scala 66:20:@46439.4]
  wire [63:0] regs_337_io_in; // @[RegFile.scala 66:20:@46439.4]
  wire  regs_337_io_reset; // @[RegFile.scala 66:20:@46439.4]
  wire [63:0] regs_337_io_out; // @[RegFile.scala 66:20:@46439.4]
  wire  regs_337_io_enable; // @[RegFile.scala 66:20:@46439.4]
  wire  regs_338_clock; // @[RegFile.scala 66:20:@46453.4]
  wire  regs_338_reset; // @[RegFile.scala 66:20:@46453.4]
  wire [63:0] regs_338_io_in; // @[RegFile.scala 66:20:@46453.4]
  wire  regs_338_io_reset; // @[RegFile.scala 66:20:@46453.4]
  wire [63:0] regs_338_io_out; // @[RegFile.scala 66:20:@46453.4]
  wire  regs_338_io_enable; // @[RegFile.scala 66:20:@46453.4]
  wire  regs_339_clock; // @[RegFile.scala 66:20:@46467.4]
  wire  regs_339_reset; // @[RegFile.scala 66:20:@46467.4]
  wire [63:0] regs_339_io_in; // @[RegFile.scala 66:20:@46467.4]
  wire  regs_339_io_reset; // @[RegFile.scala 66:20:@46467.4]
  wire [63:0] regs_339_io_out; // @[RegFile.scala 66:20:@46467.4]
  wire  regs_339_io_enable; // @[RegFile.scala 66:20:@46467.4]
  wire  regs_340_clock; // @[RegFile.scala 66:20:@46481.4]
  wire  regs_340_reset; // @[RegFile.scala 66:20:@46481.4]
  wire [63:0] regs_340_io_in; // @[RegFile.scala 66:20:@46481.4]
  wire  regs_340_io_reset; // @[RegFile.scala 66:20:@46481.4]
  wire [63:0] regs_340_io_out; // @[RegFile.scala 66:20:@46481.4]
  wire  regs_340_io_enable; // @[RegFile.scala 66:20:@46481.4]
  wire  regs_341_clock; // @[RegFile.scala 66:20:@46495.4]
  wire  regs_341_reset; // @[RegFile.scala 66:20:@46495.4]
  wire [63:0] regs_341_io_in; // @[RegFile.scala 66:20:@46495.4]
  wire  regs_341_io_reset; // @[RegFile.scala 66:20:@46495.4]
  wire [63:0] regs_341_io_out; // @[RegFile.scala 66:20:@46495.4]
  wire  regs_341_io_enable; // @[RegFile.scala 66:20:@46495.4]
  wire  regs_342_clock; // @[RegFile.scala 66:20:@46509.4]
  wire  regs_342_reset; // @[RegFile.scala 66:20:@46509.4]
  wire [63:0] regs_342_io_in; // @[RegFile.scala 66:20:@46509.4]
  wire  regs_342_io_reset; // @[RegFile.scala 66:20:@46509.4]
  wire [63:0] regs_342_io_out; // @[RegFile.scala 66:20:@46509.4]
  wire  regs_342_io_enable; // @[RegFile.scala 66:20:@46509.4]
  wire  regs_343_clock; // @[RegFile.scala 66:20:@46523.4]
  wire  regs_343_reset; // @[RegFile.scala 66:20:@46523.4]
  wire [63:0] regs_343_io_in; // @[RegFile.scala 66:20:@46523.4]
  wire  regs_343_io_reset; // @[RegFile.scala 66:20:@46523.4]
  wire [63:0] regs_343_io_out; // @[RegFile.scala 66:20:@46523.4]
  wire  regs_343_io_enable; // @[RegFile.scala 66:20:@46523.4]
  wire  regs_344_clock; // @[RegFile.scala 66:20:@46537.4]
  wire  regs_344_reset; // @[RegFile.scala 66:20:@46537.4]
  wire [63:0] regs_344_io_in; // @[RegFile.scala 66:20:@46537.4]
  wire  regs_344_io_reset; // @[RegFile.scala 66:20:@46537.4]
  wire [63:0] regs_344_io_out; // @[RegFile.scala 66:20:@46537.4]
  wire  regs_344_io_enable; // @[RegFile.scala 66:20:@46537.4]
  wire  regs_345_clock; // @[RegFile.scala 66:20:@46551.4]
  wire  regs_345_reset; // @[RegFile.scala 66:20:@46551.4]
  wire [63:0] regs_345_io_in; // @[RegFile.scala 66:20:@46551.4]
  wire  regs_345_io_reset; // @[RegFile.scala 66:20:@46551.4]
  wire [63:0] regs_345_io_out; // @[RegFile.scala 66:20:@46551.4]
  wire  regs_345_io_enable; // @[RegFile.scala 66:20:@46551.4]
  wire  regs_346_clock; // @[RegFile.scala 66:20:@46565.4]
  wire  regs_346_reset; // @[RegFile.scala 66:20:@46565.4]
  wire [63:0] regs_346_io_in; // @[RegFile.scala 66:20:@46565.4]
  wire  regs_346_io_reset; // @[RegFile.scala 66:20:@46565.4]
  wire [63:0] regs_346_io_out; // @[RegFile.scala 66:20:@46565.4]
  wire  regs_346_io_enable; // @[RegFile.scala 66:20:@46565.4]
  wire  regs_347_clock; // @[RegFile.scala 66:20:@46579.4]
  wire  regs_347_reset; // @[RegFile.scala 66:20:@46579.4]
  wire [63:0] regs_347_io_in; // @[RegFile.scala 66:20:@46579.4]
  wire  regs_347_io_reset; // @[RegFile.scala 66:20:@46579.4]
  wire [63:0] regs_347_io_out; // @[RegFile.scala 66:20:@46579.4]
  wire  regs_347_io_enable; // @[RegFile.scala 66:20:@46579.4]
  wire  regs_348_clock; // @[RegFile.scala 66:20:@46593.4]
  wire  regs_348_reset; // @[RegFile.scala 66:20:@46593.4]
  wire [63:0] regs_348_io_in; // @[RegFile.scala 66:20:@46593.4]
  wire  regs_348_io_reset; // @[RegFile.scala 66:20:@46593.4]
  wire [63:0] regs_348_io_out; // @[RegFile.scala 66:20:@46593.4]
  wire  regs_348_io_enable; // @[RegFile.scala 66:20:@46593.4]
  wire  regs_349_clock; // @[RegFile.scala 66:20:@46607.4]
  wire  regs_349_reset; // @[RegFile.scala 66:20:@46607.4]
  wire [63:0] regs_349_io_in; // @[RegFile.scala 66:20:@46607.4]
  wire  regs_349_io_reset; // @[RegFile.scala 66:20:@46607.4]
  wire [63:0] regs_349_io_out; // @[RegFile.scala 66:20:@46607.4]
  wire  regs_349_io_enable; // @[RegFile.scala 66:20:@46607.4]
  wire  regs_350_clock; // @[RegFile.scala 66:20:@46621.4]
  wire  regs_350_reset; // @[RegFile.scala 66:20:@46621.4]
  wire [63:0] regs_350_io_in; // @[RegFile.scala 66:20:@46621.4]
  wire  regs_350_io_reset; // @[RegFile.scala 66:20:@46621.4]
  wire [63:0] regs_350_io_out; // @[RegFile.scala 66:20:@46621.4]
  wire  regs_350_io_enable; // @[RegFile.scala 66:20:@46621.4]
  wire  regs_351_clock; // @[RegFile.scala 66:20:@46635.4]
  wire  regs_351_reset; // @[RegFile.scala 66:20:@46635.4]
  wire [63:0] regs_351_io_in; // @[RegFile.scala 66:20:@46635.4]
  wire  regs_351_io_reset; // @[RegFile.scala 66:20:@46635.4]
  wire [63:0] regs_351_io_out; // @[RegFile.scala 66:20:@46635.4]
  wire  regs_351_io_enable; // @[RegFile.scala 66:20:@46635.4]
  wire  regs_352_clock; // @[RegFile.scala 66:20:@46649.4]
  wire  regs_352_reset; // @[RegFile.scala 66:20:@46649.4]
  wire [63:0] regs_352_io_in; // @[RegFile.scala 66:20:@46649.4]
  wire  regs_352_io_reset; // @[RegFile.scala 66:20:@46649.4]
  wire [63:0] regs_352_io_out; // @[RegFile.scala 66:20:@46649.4]
  wire  regs_352_io_enable; // @[RegFile.scala 66:20:@46649.4]
  wire  regs_353_clock; // @[RegFile.scala 66:20:@46663.4]
  wire  regs_353_reset; // @[RegFile.scala 66:20:@46663.4]
  wire [63:0] regs_353_io_in; // @[RegFile.scala 66:20:@46663.4]
  wire  regs_353_io_reset; // @[RegFile.scala 66:20:@46663.4]
  wire [63:0] regs_353_io_out; // @[RegFile.scala 66:20:@46663.4]
  wire  regs_353_io_enable; // @[RegFile.scala 66:20:@46663.4]
  wire  regs_354_clock; // @[RegFile.scala 66:20:@46677.4]
  wire  regs_354_reset; // @[RegFile.scala 66:20:@46677.4]
  wire [63:0] regs_354_io_in; // @[RegFile.scala 66:20:@46677.4]
  wire  regs_354_io_reset; // @[RegFile.scala 66:20:@46677.4]
  wire [63:0] regs_354_io_out; // @[RegFile.scala 66:20:@46677.4]
  wire  regs_354_io_enable; // @[RegFile.scala 66:20:@46677.4]
  wire  regs_355_clock; // @[RegFile.scala 66:20:@46691.4]
  wire  regs_355_reset; // @[RegFile.scala 66:20:@46691.4]
  wire [63:0] regs_355_io_in; // @[RegFile.scala 66:20:@46691.4]
  wire  regs_355_io_reset; // @[RegFile.scala 66:20:@46691.4]
  wire [63:0] regs_355_io_out; // @[RegFile.scala 66:20:@46691.4]
  wire  regs_355_io_enable; // @[RegFile.scala 66:20:@46691.4]
  wire  regs_356_clock; // @[RegFile.scala 66:20:@46705.4]
  wire  regs_356_reset; // @[RegFile.scala 66:20:@46705.4]
  wire [63:0] regs_356_io_in; // @[RegFile.scala 66:20:@46705.4]
  wire  regs_356_io_reset; // @[RegFile.scala 66:20:@46705.4]
  wire [63:0] regs_356_io_out; // @[RegFile.scala 66:20:@46705.4]
  wire  regs_356_io_enable; // @[RegFile.scala 66:20:@46705.4]
  wire  regs_357_clock; // @[RegFile.scala 66:20:@46719.4]
  wire  regs_357_reset; // @[RegFile.scala 66:20:@46719.4]
  wire [63:0] regs_357_io_in; // @[RegFile.scala 66:20:@46719.4]
  wire  regs_357_io_reset; // @[RegFile.scala 66:20:@46719.4]
  wire [63:0] regs_357_io_out; // @[RegFile.scala 66:20:@46719.4]
  wire  regs_357_io_enable; // @[RegFile.scala 66:20:@46719.4]
  wire  regs_358_clock; // @[RegFile.scala 66:20:@46733.4]
  wire  regs_358_reset; // @[RegFile.scala 66:20:@46733.4]
  wire [63:0] regs_358_io_in; // @[RegFile.scala 66:20:@46733.4]
  wire  regs_358_io_reset; // @[RegFile.scala 66:20:@46733.4]
  wire [63:0] regs_358_io_out; // @[RegFile.scala 66:20:@46733.4]
  wire  regs_358_io_enable; // @[RegFile.scala 66:20:@46733.4]
  wire  regs_359_clock; // @[RegFile.scala 66:20:@46747.4]
  wire  regs_359_reset; // @[RegFile.scala 66:20:@46747.4]
  wire [63:0] regs_359_io_in; // @[RegFile.scala 66:20:@46747.4]
  wire  regs_359_io_reset; // @[RegFile.scala 66:20:@46747.4]
  wire [63:0] regs_359_io_out; // @[RegFile.scala 66:20:@46747.4]
  wire  regs_359_io_enable; // @[RegFile.scala 66:20:@46747.4]
  wire  regs_360_clock; // @[RegFile.scala 66:20:@46761.4]
  wire  regs_360_reset; // @[RegFile.scala 66:20:@46761.4]
  wire [63:0] regs_360_io_in; // @[RegFile.scala 66:20:@46761.4]
  wire  regs_360_io_reset; // @[RegFile.scala 66:20:@46761.4]
  wire [63:0] regs_360_io_out; // @[RegFile.scala 66:20:@46761.4]
  wire  regs_360_io_enable; // @[RegFile.scala 66:20:@46761.4]
  wire  regs_361_clock; // @[RegFile.scala 66:20:@46775.4]
  wire  regs_361_reset; // @[RegFile.scala 66:20:@46775.4]
  wire [63:0] regs_361_io_in; // @[RegFile.scala 66:20:@46775.4]
  wire  regs_361_io_reset; // @[RegFile.scala 66:20:@46775.4]
  wire [63:0] regs_361_io_out; // @[RegFile.scala 66:20:@46775.4]
  wire  regs_361_io_enable; // @[RegFile.scala 66:20:@46775.4]
  wire  regs_362_clock; // @[RegFile.scala 66:20:@46789.4]
  wire  regs_362_reset; // @[RegFile.scala 66:20:@46789.4]
  wire [63:0] regs_362_io_in; // @[RegFile.scala 66:20:@46789.4]
  wire  regs_362_io_reset; // @[RegFile.scala 66:20:@46789.4]
  wire [63:0] regs_362_io_out; // @[RegFile.scala 66:20:@46789.4]
  wire  regs_362_io_enable; // @[RegFile.scala 66:20:@46789.4]
  wire  regs_363_clock; // @[RegFile.scala 66:20:@46803.4]
  wire  regs_363_reset; // @[RegFile.scala 66:20:@46803.4]
  wire [63:0] regs_363_io_in; // @[RegFile.scala 66:20:@46803.4]
  wire  regs_363_io_reset; // @[RegFile.scala 66:20:@46803.4]
  wire [63:0] regs_363_io_out; // @[RegFile.scala 66:20:@46803.4]
  wire  regs_363_io_enable; // @[RegFile.scala 66:20:@46803.4]
  wire  regs_364_clock; // @[RegFile.scala 66:20:@46817.4]
  wire  regs_364_reset; // @[RegFile.scala 66:20:@46817.4]
  wire [63:0] regs_364_io_in; // @[RegFile.scala 66:20:@46817.4]
  wire  regs_364_io_reset; // @[RegFile.scala 66:20:@46817.4]
  wire [63:0] regs_364_io_out; // @[RegFile.scala 66:20:@46817.4]
  wire  regs_364_io_enable; // @[RegFile.scala 66:20:@46817.4]
  wire  regs_365_clock; // @[RegFile.scala 66:20:@46831.4]
  wire  regs_365_reset; // @[RegFile.scala 66:20:@46831.4]
  wire [63:0] regs_365_io_in; // @[RegFile.scala 66:20:@46831.4]
  wire  regs_365_io_reset; // @[RegFile.scala 66:20:@46831.4]
  wire [63:0] regs_365_io_out; // @[RegFile.scala 66:20:@46831.4]
  wire  regs_365_io_enable; // @[RegFile.scala 66:20:@46831.4]
  wire  regs_366_clock; // @[RegFile.scala 66:20:@46845.4]
  wire  regs_366_reset; // @[RegFile.scala 66:20:@46845.4]
  wire [63:0] regs_366_io_in; // @[RegFile.scala 66:20:@46845.4]
  wire  regs_366_io_reset; // @[RegFile.scala 66:20:@46845.4]
  wire [63:0] regs_366_io_out; // @[RegFile.scala 66:20:@46845.4]
  wire  regs_366_io_enable; // @[RegFile.scala 66:20:@46845.4]
  wire  regs_367_clock; // @[RegFile.scala 66:20:@46859.4]
  wire  regs_367_reset; // @[RegFile.scala 66:20:@46859.4]
  wire [63:0] regs_367_io_in; // @[RegFile.scala 66:20:@46859.4]
  wire  regs_367_io_reset; // @[RegFile.scala 66:20:@46859.4]
  wire [63:0] regs_367_io_out; // @[RegFile.scala 66:20:@46859.4]
  wire  regs_367_io_enable; // @[RegFile.scala 66:20:@46859.4]
  wire  regs_368_clock; // @[RegFile.scala 66:20:@46873.4]
  wire  regs_368_reset; // @[RegFile.scala 66:20:@46873.4]
  wire [63:0] regs_368_io_in; // @[RegFile.scala 66:20:@46873.4]
  wire  regs_368_io_reset; // @[RegFile.scala 66:20:@46873.4]
  wire [63:0] regs_368_io_out; // @[RegFile.scala 66:20:@46873.4]
  wire  regs_368_io_enable; // @[RegFile.scala 66:20:@46873.4]
  wire  regs_369_clock; // @[RegFile.scala 66:20:@46887.4]
  wire  regs_369_reset; // @[RegFile.scala 66:20:@46887.4]
  wire [63:0] regs_369_io_in; // @[RegFile.scala 66:20:@46887.4]
  wire  regs_369_io_reset; // @[RegFile.scala 66:20:@46887.4]
  wire [63:0] regs_369_io_out; // @[RegFile.scala 66:20:@46887.4]
  wire  regs_369_io_enable; // @[RegFile.scala 66:20:@46887.4]
  wire  regs_370_clock; // @[RegFile.scala 66:20:@46901.4]
  wire  regs_370_reset; // @[RegFile.scala 66:20:@46901.4]
  wire [63:0] regs_370_io_in; // @[RegFile.scala 66:20:@46901.4]
  wire  regs_370_io_reset; // @[RegFile.scala 66:20:@46901.4]
  wire [63:0] regs_370_io_out; // @[RegFile.scala 66:20:@46901.4]
  wire  regs_370_io_enable; // @[RegFile.scala 66:20:@46901.4]
  wire  regs_371_clock; // @[RegFile.scala 66:20:@46915.4]
  wire  regs_371_reset; // @[RegFile.scala 66:20:@46915.4]
  wire [63:0] regs_371_io_in; // @[RegFile.scala 66:20:@46915.4]
  wire  regs_371_io_reset; // @[RegFile.scala 66:20:@46915.4]
  wire [63:0] regs_371_io_out; // @[RegFile.scala 66:20:@46915.4]
  wire  regs_371_io_enable; // @[RegFile.scala 66:20:@46915.4]
  wire  regs_372_clock; // @[RegFile.scala 66:20:@46929.4]
  wire  regs_372_reset; // @[RegFile.scala 66:20:@46929.4]
  wire [63:0] regs_372_io_in; // @[RegFile.scala 66:20:@46929.4]
  wire  regs_372_io_reset; // @[RegFile.scala 66:20:@46929.4]
  wire [63:0] regs_372_io_out; // @[RegFile.scala 66:20:@46929.4]
  wire  regs_372_io_enable; // @[RegFile.scala 66:20:@46929.4]
  wire  regs_373_clock; // @[RegFile.scala 66:20:@46943.4]
  wire  regs_373_reset; // @[RegFile.scala 66:20:@46943.4]
  wire [63:0] regs_373_io_in; // @[RegFile.scala 66:20:@46943.4]
  wire  regs_373_io_reset; // @[RegFile.scala 66:20:@46943.4]
  wire [63:0] regs_373_io_out; // @[RegFile.scala 66:20:@46943.4]
  wire  regs_373_io_enable; // @[RegFile.scala 66:20:@46943.4]
  wire  regs_374_clock; // @[RegFile.scala 66:20:@46957.4]
  wire  regs_374_reset; // @[RegFile.scala 66:20:@46957.4]
  wire [63:0] regs_374_io_in; // @[RegFile.scala 66:20:@46957.4]
  wire  regs_374_io_reset; // @[RegFile.scala 66:20:@46957.4]
  wire [63:0] regs_374_io_out; // @[RegFile.scala 66:20:@46957.4]
  wire  regs_374_io_enable; // @[RegFile.scala 66:20:@46957.4]
  wire  regs_375_clock; // @[RegFile.scala 66:20:@46971.4]
  wire  regs_375_reset; // @[RegFile.scala 66:20:@46971.4]
  wire [63:0] regs_375_io_in; // @[RegFile.scala 66:20:@46971.4]
  wire  regs_375_io_reset; // @[RegFile.scala 66:20:@46971.4]
  wire [63:0] regs_375_io_out; // @[RegFile.scala 66:20:@46971.4]
  wire  regs_375_io_enable; // @[RegFile.scala 66:20:@46971.4]
  wire  regs_376_clock; // @[RegFile.scala 66:20:@46985.4]
  wire  regs_376_reset; // @[RegFile.scala 66:20:@46985.4]
  wire [63:0] regs_376_io_in; // @[RegFile.scala 66:20:@46985.4]
  wire  regs_376_io_reset; // @[RegFile.scala 66:20:@46985.4]
  wire [63:0] regs_376_io_out; // @[RegFile.scala 66:20:@46985.4]
  wire  regs_376_io_enable; // @[RegFile.scala 66:20:@46985.4]
  wire  regs_377_clock; // @[RegFile.scala 66:20:@46999.4]
  wire  regs_377_reset; // @[RegFile.scala 66:20:@46999.4]
  wire [63:0] regs_377_io_in; // @[RegFile.scala 66:20:@46999.4]
  wire  regs_377_io_reset; // @[RegFile.scala 66:20:@46999.4]
  wire [63:0] regs_377_io_out; // @[RegFile.scala 66:20:@46999.4]
  wire  regs_377_io_enable; // @[RegFile.scala 66:20:@46999.4]
  wire  regs_378_clock; // @[RegFile.scala 66:20:@47013.4]
  wire  regs_378_reset; // @[RegFile.scala 66:20:@47013.4]
  wire [63:0] regs_378_io_in; // @[RegFile.scala 66:20:@47013.4]
  wire  regs_378_io_reset; // @[RegFile.scala 66:20:@47013.4]
  wire [63:0] regs_378_io_out; // @[RegFile.scala 66:20:@47013.4]
  wire  regs_378_io_enable; // @[RegFile.scala 66:20:@47013.4]
  wire  regs_379_clock; // @[RegFile.scala 66:20:@47027.4]
  wire  regs_379_reset; // @[RegFile.scala 66:20:@47027.4]
  wire [63:0] regs_379_io_in; // @[RegFile.scala 66:20:@47027.4]
  wire  regs_379_io_reset; // @[RegFile.scala 66:20:@47027.4]
  wire [63:0] regs_379_io_out; // @[RegFile.scala 66:20:@47027.4]
  wire  regs_379_io_enable; // @[RegFile.scala 66:20:@47027.4]
  wire  regs_380_clock; // @[RegFile.scala 66:20:@47041.4]
  wire  regs_380_reset; // @[RegFile.scala 66:20:@47041.4]
  wire [63:0] regs_380_io_in; // @[RegFile.scala 66:20:@47041.4]
  wire  regs_380_io_reset; // @[RegFile.scala 66:20:@47041.4]
  wire [63:0] regs_380_io_out; // @[RegFile.scala 66:20:@47041.4]
  wire  regs_380_io_enable; // @[RegFile.scala 66:20:@47041.4]
  wire  regs_381_clock; // @[RegFile.scala 66:20:@47055.4]
  wire  regs_381_reset; // @[RegFile.scala 66:20:@47055.4]
  wire [63:0] regs_381_io_in; // @[RegFile.scala 66:20:@47055.4]
  wire  regs_381_io_reset; // @[RegFile.scala 66:20:@47055.4]
  wire [63:0] regs_381_io_out; // @[RegFile.scala 66:20:@47055.4]
  wire  regs_381_io_enable; // @[RegFile.scala 66:20:@47055.4]
  wire  regs_382_clock; // @[RegFile.scala 66:20:@47069.4]
  wire  regs_382_reset; // @[RegFile.scala 66:20:@47069.4]
  wire [63:0] regs_382_io_in; // @[RegFile.scala 66:20:@47069.4]
  wire  regs_382_io_reset; // @[RegFile.scala 66:20:@47069.4]
  wire [63:0] regs_382_io_out; // @[RegFile.scala 66:20:@47069.4]
  wire  regs_382_io_enable; // @[RegFile.scala 66:20:@47069.4]
  wire  regs_383_clock; // @[RegFile.scala 66:20:@47083.4]
  wire  regs_383_reset; // @[RegFile.scala 66:20:@47083.4]
  wire [63:0] regs_383_io_in; // @[RegFile.scala 66:20:@47083.4]
  wire  regs_383_io_reset; // @[RegFile.scala 66:20:@47083.4]
  wire [63:0] regs_383_io_out; // @[RegFile.scala 66:20:@47083.4]
  wire  regs_383_io_enable; // @[RegFile.scala 66:20:@47083.4]
  wire  regs_384_clock; // @[RegFile.scala 66:20:@47097.4]
  wire  regs_384_reset; // @[RegFile.scala 66:20:@47097.4]
  wire [63:0] regs_384_io_in; // @[RegFile.scala 66:20:@47097.4]
  wire  regs_384_io_reset; // @[RegFile.scala 66:20:@47097.4]
  wire [63:0] regs_384_io_out; // @[RegFile.scala 66:20:@47097.4]
  wire  regs_384_io_enable; // @[RegFile.scala 66:20:@47097.4]
  wire  regs_385_clock; // @[RegFile.scala 66:20:@47111.4]
  wire  regs_385_reset; // @[RegFile.scala 66:20:@47111.4]
  wire [63:0] regs_385_io_in; // @[RegFile.scala 66:20:@47111.4]
  wire  regs_385_io_reset; // @[RegFile.scala 66:20:@47111.4]
  wire [63:0] regs_385_io_out; // @[RegFile.scala 66:20:@47111.4]
  wire  regs_385_io_enable; // @[RegFile.scala 66:20:@47111.4]
  wire  regs_386_clock; // @[RegFile.scala 66:20:@47125.4]
  wire  regs_386_reset; // @[RegFile.scala 66:20:@47125.4]
  wire [63:0] regs_386_io_in; // @[RegFile.scala 66:20:@47125.4]
  wire  regs_386_io_reset; // @[RegFile.scala 66:20:@47125.4]
  wire [63:0] regs_386_io_out; // @[RegFile.scala 66:20:@47125.4]
  wire  regs_386_io_enable; // @[RegFile.scala 66:20:@47125.4]
  wire  regs_387_clock; // @[RegFile.scala 66:20:@47139.4]
  wire  regs_387_reset; // @[RegFile.scala 66:20:@47139.4]
  wire [63:0] regs_387_io_in; // @[RegFile.scala 66:20:@47139.4]
  wire  regs_387_io_reset; // @[RegFile.scala 66:20:@47139.4]
  wire [63:0] regs_387_io_out; // @[RegFile.scala 66:20:@47139.4]
  wire  regs_387_io_enable; // @[RegFile.scala 66:20:@47139.4]
  wire  regs_388_clock; // @[RegFile.scala 66:20:@47153.4]
  wire  regs_388_reset; // @[RegFile.scala 66:20:@47153.4]
  wire [63:0] regs_388_io_in; // @[RegFile.scala 66:20:@47153.4]
  wire  regs_388_io_reset; // @[RegFile.scala 66:20:@47153.4]
  wire [63:0] regs_388_io_out; // @[RegFile.scala 66:20:@47153.4]
  wire  regs_388_io_enable; // @[RegFile.scala 66:20:@47153.4]
  wire  regs_389_clock; // @[RegFile.scala 66:20:@47167.4]
  wire  regs_389_reset; // @[RegFile.scala 66:20:@47167.4]
  wire [63:0] regs_389_io_in; // @[RegFile.scala 66:20:@47167.4]
  wire  regs_389_io_reset; // @[RegFile.scala 66:20:@47167.4]
  wire [63:0] regs_389_io_out; // @[RegFile.scala 66:20:@47167.4]
  wire  regs_389_io_enable; // @[RegFile.scala 66:20:@47167.4]
  wire  regs_390_clock; // @[RegFile.scala 66:20:@47181.4]
  wire  regs_390_reset; // @[RegFile.scala 66:20:@47181.4]
  wire [63:0] regs_390_io_in; // @[RegFile.scala 66:20:@47181.4]
  wire  regs_390_io_reset; // @[RegFile.scala 66:20:@47181.4]
  wire [63:0] regs_390_io_out; // @[RegFile.scala 66:20:@47181.4]
  wire  regs_390_io_enable; // @[RegFile.scala 66:20:@47181.4]
  wire  regs_391_clock; // @[RegFile.scala 66:20:@47195.4]
  wire  regs_391_reset; // @[RegFile.scala 66:20:@47195.4]
  wire [63:0] regs_391_io_in; // @[RegFile.scala 66:20:@47195.4]
  wire  regs_391_io_reset; // @[RegFile.scala 66:20:@47195.4]
  wire [63:0] regs_391_io_out; // @[RegFile.scala 66:20:@47195.4]
  wire  regs_391_io_enable; // @[RegFile.scala 66:20:@47195.4]
  wire  regs_392_clock; // @[RegFile.scala 66:20:@47209.4]
  wire  regs_392_reset; // @[RegFile.scala 66:20:@47209.4]
  wire [63:0] regs_392_io_in; // @[RegFile.scala 66:20:@47209.4]
  wire  regs_392_io_reset; // @[RegFile.scala 66:20:@47209.4]
  wire [63:0] regs_392_io_out; // @[RegFile.scala 66:20:@47209.4]
  wire  regs_392_io_enable; // @[RegFile.scala 66:20:@47209.4]
  wire  regs_393_clock; // @[RegFile.scala 66:20:@47223.4]
  wire  regs_393_reset; // @[RegFile.scala 66:20:@47223.4]
  wire [63:0] regs_393_io_in; // @[RegFile.scala 66:20:@47223.4]
  wire  regs_393_io_reset; // @[RegFile.scala 66:20:@47223.4]
  wire [63:0] regs_393_io_out; // @[RegFile.scala 66:20:@47223.4]
  wire  regs_393_io_enable; // @[RegFile.scala 66:20:@47223.4]
  wire  regs_394_clock; // @[RegFile.scala 66:20:@47237.4]
  wire  regs_394_reset; // @[RegFile.scala 66:20:@47237.4]
  wire [63:0] regs_394_io_in; // @[RegFile.scala 66:20:@47237.4]
  wire  regs_394_io_reset; // @[RegFile.scala 66:20:@47237.4]
  wire [63:0] regs_394_io_out; // @[RegFile.scala 66:20:@47237.4]
  wire  regs_394_io_enable; // @[RegFile.scala 66:20:@47237.4]
  wire  regs_395_clock; // @[RegFile.scala 66:20:@47251.4]
  wire  regs_395_reset; // @[RegFile.scala 66:20:@47251.4]
  wire [63:0] regs_395_io_in; // @[RegFile.scala 66:20:@47251.4]
  wire  regs_395_io_reset; // @[RegFile.scala 66:20:@47251.4]
  wire [63:0] regs_395_io_out; // @[RegFile.scala 66:20:@47251.4]
  wire  regs_395_io_enable; // @[RegFile.scala 66:20:@47251.4]
  wire  regs_396_clock; // @[RegFile.scala 66:20:@47265.4]
  wire  regs_396_reset; // @[RegFile.scala 66:20:@47265.4]
  wire [63:0] regs_396_io_in; // @[RegFile.scala 66:20:@47265.4]
  wire  regs_396_io_reset; // @[RegFile.scala 66:20:@47265.4]
  wire [63:0] regs_396_io_out; // @[RegFile.scala 66:20:@47265.4]
  wire  regs_396_io_enable; // @[RegFile.scala 66:20:@47265.4]
  wire  regs_397_clock; // @[RegFile.scala 66:20:@47279.4]
  wire  regs_397_reset; // @[RegFile.scala 66:20:@47279.4]
  wire [63:0] regs_397_io_in; // @[RegFile.scala 66:20:@47279.4]
  wire  regs_397_io_reset; // @[RegFile.scala 66:20:@47279.4]
  wire [63:0] regs_397_io_out; // @[RegFile.scala 66:20:@47279.4]
  wire  regs_397_io_enable; // @[RegFile.scala 66:20:@47279.4]
  wire  regs_398_clock; // @[RegFile.scala 66:20:@47293.4]
  wire  regs_398_reset; // @[RegFile.scala 66:20:@47293.4]
  wire [63:0] regs_398_io_in; // @[RegFile.scala 66:20:@47293.4]
  wire  regs_398_io_reset; // @[RegFile.scala 66:20:@47293.4]
  wire [63:0] regs_398_io_out; // @[RegFile.scala 66:20:@47293.4]
  wire  regs_398_io_enable; // @[RegFile.scala 66:20:@47293.4]
  wire  regs_399_clock; // @[RegFile.scala 66:20:@47307.4]
  wire  regs_399_reset; // @[RegFile.scala 66:20:@47307.4]
  wire [63:0] regs_399_io_in; // @[RegFile.scala 66:20:@47307.4]
  wire  regs_399_io_reset; // @[RegFile.scala 66:20:@47307.4]
  wire [63:0] regs_399_io_out; // @[RegFile.scala 66:20:@47307.4]
  wire  regs_399_io_enable; // @[RegFile.scala 66:20:@47307.4]
  wire  regs_400_clock; // @[RegFile.scala 66:20:@47321.4]
  wire  regs_400_reset; // @[RegFile.scala 66:20:@47321.4]
  wire [63:0] regs_400_io_in; // @[RegFile.scala 66:20:@47321.4]
  wire  regs_400_io_reset; // @[RegFile.scala 66:20:@47321.4]
  wire [63:0] regs_400_io_out; // @[RegFile.scala 66:20:@47321.4]
  wire  regs_400_io_enable; // @[RegFile.scala 66:20:@47321.4]
  wire  regs_401_clock; // @[RegFile.scala 66:20:@47335.4]
  wire  regs_401_reset; // @[RegFile.scala 66:20:@47335.4]
  wire [63:0] regs_401_io_in; // @[RegFile.scala 66:20:@47335.4]
  wire  regs_401_io_reset; // @[RegFile.scala 66:20:@47335.4]
  wire [63:0] regs_401_io_out; // @[RegFile.scala 66:20:@47335.4]
  wire  regs_401_io_enable; // @[RegFile.scala 66:20:@47335.4]
  wire  regs_402_clock; // @[RegFile.scala 66:20:@47349.4]
  wire  regs_402_reset; // @[RegFile.scala 66:20:@47349.4]
  wire [63:0] regs_402_io_in; // @[RegFile.scala 66:20:@47349.4]
  wire  regs_402_io_reset; // @[RegFile.scala 66:20:@47349.4]
  wire [63:0] regs_402_io_out; // @[RegFile.scala 66:20:@47349.4]
  wire  regs_402_io_enable; // @[RegFile.scala 66:20:@47349.4]
  wire  regs_403_clock; // @[RegFile.scala 66:20:@47363.4]
  wire  regs_403_reset; // @[RegFile.scala 66:20:@47363.4]
  wire [63:0] regs_403_io_in; // @[RegFile.scala 66:20:@47363.4]
  wire  regs_403_io_reset; // @[RegFile.scala 66:20:@47363.4]
  wire [63:0] regs_403_io_out; // @[RegFile.scala 66:20:@47363.4]
  wire  regs_403_io_enable; // @[RegFile.scala 66:20:@47363.4]
  wire  regs_404_clock; // @[RegFile.scala 66:20:@47377.4]
  wire  regs_404_reset; // @[RegFile.scala 66:20:@47377.4]
  wire [63:0] regs_404_io_in; // @[RegFile.scala 66:20:@47377.4]
  wire  regs_404_io_reset; // @[RegFile.scala 66:20:@47377.4]
  wire [63:0] regs_404_io_out; // @[RegFile.scala 66:20:@47377.4]
  wire  regs_404_io_enable; // @[RegFile.scala 66:20:@47377.4]
  wire  regs_405_clock; // @[RegFile.scala 66:20:@47391.4]
  wire  regs_405_reset; // @[RegFile.scala 66:20:@47391.4]
  wire [63:0] regs_405_io_in; // @[RegFile.scala 66:20:@47391.4]
  wire  regs_405_io_reset; // @[RegFile.scala 66:20:@47391.4]
  wire [63:0] regs_405_io_out; // @[RegFile.scala 66:20:@47391.4]
  wire  regs_405_io_enable; // @[RegFile.scala 66:20:@47391.4]
  wire  regs_406_clock; // @[RegFile.scala 66:20:@47405.4]
  wire  regs_406_reset; // @[RegFile.scala 66:20:@47405.4]
  wire [63:0] regs_406_io_in; // @[RegFile.scala 66:20:@47405.4]
  wire  regs_406_io_reset; // @[RegFile.scala 66:20:@47405.4]
  wire [63:0] regs_406_io_out; // @[RegFile.scala 66:20:@47405.4]
  wire  regs_406_io_enable; // @[RegFile.scala 66:20:@47405.4]
  wire  regs_407_clock; // @[RegFile.scala 66:20:@47419.4]
  wire  regs_407_reset; // @[RegFile.scala 66:20:@47419.4]
  wire [63:0] regs_407_io_in; // @[RegFile.scala 66:20:@47419.4]
  wire  regs_407_io_reset; // @[RegFile.scala 66:20:@47419.4]
  wire [63:0] regs_407_io_out; // @[RegFile.scala 66:20:@47419.4]
  wire  regs_407_io_enable; // @[RegFile.scala 66:20:@47419.4]
  wire  regs_408_clock; // @[RegFile.scala 66:20:@47433.4]
  wire  regs_408_reset; // @[RegFile.scala 66:20:@47433.4]
  wire [63:0] regs_408_io_in; // @[RegFile.scala 66:20:@47433.4]
  wire  regs_408_io_reset; // @[RegFile.scala 66:20:@47433.4]
  wire [63:0] regs_408_io_out; // @[RegFile.scala 66:20:@47433.4]
  wire  regs_408_io_enable; // @[RegFile.scala 66:20:@47433.4]
  wire  regs_409_clock; // @[RegFile.scala 66:20:@47447.4]
  wire  regs_409_reset; // @[RegFile.scala 66:20:@47447.4]
  wire [63:0] regs_409_io_in; // @[RegFile.scala 66:20:@47447.4]
  wire  regs_409_io_reset; // @[RegFile.scala 66:20:@47447.4]
  wire [63:0] regs_409_io_out; // @[RegFile.scala 66:20:@47447.4]
  wire  regs_409_io_enable; // @[RegFile.scala 66:20:@47447.4]
  wire  regs_410_clock; // @[RegFile.scala 66:20:@47461.4]
  wire  regs_410_reset; // @[RegFile.scala 66:20:@47461.4]
  wire [63:0] regs_410_io_in; // @[RegFile.scala 66:20:@47461.4]
  wire  regs_410_io_reset; // @[RegFile.scala 66:20:@47461.4]
  wire [63:0] regs_410_io_out; // @[RegFile.scala 66:20:@47461.4]
  wire  regs_410_io_enable; // @[RegFile.scala 66:20:@47461.4]
  wire  regs_411_clock; // @[RegFile.scala 66:20:@47475.4]
  wire  regs_411_reset; // @[RegFile.scala 66:20:@47475.4]
  wire [63:0] regs_411_io_in; // @[RegFile.scala 66:20:@47475.4]
  wire  regs_411_io_reset; // @[RegFile.scala 66:20:@47475.4]
  wire [63:0] regs_411_io_out; // @[RegFile.scala 66:20:@47475.4]
  wire  regs_411_io_enable; // @[RegFile.scala 66:20:@47475.4]
  wire  regs_412_clock; // @[RegFile.scala 66:20:@47489.4]
  wire  regs_412_reset; // @[RegFile.scala 66:20:@47489.4]
  wire [63:0] regs_412_io_in; // @[RegFile.scala 66:20:@47489.4]
  wire  regs_412_io_reset; // @[RegFile.scala 66:20:@47489.4]
  wire [63:0] regs_412_io_out; // @[RegFile.scala 66:20:@47489.4]
  wire  regs_412_io_enable; // @[RegFile.scala 66:20:@47489.4]
  wire  regs_413_clock; // @[RegFile.scala 66:20:@47503.4]
  wire  regs_413_reset; // @[RegFile.scala 66:20:@47503.4]
  wire [63:0] regs_413_io_in; // @[RegFile.scala 66:20:@47503.4]
  wire  regs_413_io_reset; // @[RegFile.scala 66:20:@47503.4]
  wire [63:0] regs_413_io_out; // @[RegFile.scala 66:20:@47503.4]
  wire  regs_413_io_enable; // @[RegFile.scala 66:20:@47503.4]
  wire  regs_414_clock; // @[RegFile.scala 66:20:@47517.4]
  wire  regs_414_reset; // @[RegFile.scala 66:20:@47517.4]
  wire [63:0] regs_414_io_in; // @[RegFile.scala 66:20:@47517.4]
  wire  regs_414_io_reset; // @[RegFile.scala 66:20:@47517.4]
  wire [63:0] regs_414_io_out; // @[RegFile.scala 66:20:@47517.4]
  wire  regs_414_io_enable; // @[RegFile.scala 66:20:@47517.4]
  wire  regs_415_clock; // @[RegFile.scala 66:20:@47531.4]
  wire  regs_415_reset; // @[RegFile.scala 66:20:@47531.4]
  wire [63:0] regs_415_io_in; // @[RegFile.scala 66:20:@47531.4]
  wire  regs_415_io_reset; // @[RegFile.scala 66:20:@47531.4]
  wire [63:0] regs_415_io_out; // @[RegFile.scala 66:20:@47531.4]
  wire  regs_415_io_enable; // @[RegFile.scala 66:20:@47531.4]
  wire  regs_416_clock; // @[RegFile.scala 66:20:@47545.4]
  wire  regs_416_reset; // @[RegFile.scala 66:20:@47545.4]
  wire [63:0] regs_416_io_in; // @[RegFile.scala 66:20:@47545.4]
  wire  regs_416_io_reset; // @[RegFile.scala 66:20:@47545.4]
  wire [63:0] regs_416_io_out; // @[RegFile.scala 66:20:@47545.4]
  wire  regs_416_io_enable; // @[RegFile.scala 66:20:@47545.4]
  wire  regs_417_clock; // @[RegFile.scala 66:20:@47559.4]
  wire  regs_417_reset; // @[RegFile.scala 66:20:@47559.4]
  wire [63:0] regs_417_io_in; // @[RegFile.scala 66:20:@47559.4]
  wire  regs_417_io_reset; // @[RegFile.scala 66:20:@47559.4]
  wire [63:0] regs_417_io_out; // @[RegFile.scala 66:20:@47559.4]
  wire  regs_417_io_enable; // @[RegFile.scala 66:20:@47559.4]
  wire  regs_418_clock; // @[RegFile.scala 66:20:@47573.4]
  wire  regs_418_reset; // @[RegFile.scala 66:20:@47573.4]
  wire [63:0] regs_418_io_in; // @[RegFile.scala 66:20:@47573.4]
  wire  regs_418_io_reset; // @[RegFile.scala 66:20:@47573.4]
  wire [63:0] regs_418_io_out; // @[RegFile.scala 66:20:@47573.4]
  wire  regs_418_io_enable; // @[RegFile.scala 66:20:@47573.4]
  wire  regs_419_clock; // @[RegFile.scala 66:20:@47587.4]
  wire  regs_419_reset; // @[RegFile.scala 66:20:@47587.4]
  wire [63:0] regs_419_io_in; // @[RegFile.scala 66:20:@47587.4]
  wire  regs_419_io_reset; // @[RegFile.scala 66:20:@47587.4]
  wire [63:0] regs_419_io_out; // @[RegFile.scala 66:20:@47587.4]
  wire  regs_419_io_enable; // @[RegFile.scala 66:20:@47587.4]
  wire  regs_420_clock; // @[RegFile.scala 66:20:@47601.4]
  wire  regs_420_reset; // @[RegFile.scala 66:20:@47601.4]
  wire [63:0] regs_420_io_in; // @[RegFile.scala 66:20:@47601.4]
  wire  regs_420_io_reset; // @[RegFile.scala 66:20:@47601.4]
  wire [63:0] regs_420_io_out; // @[RegFile.scala 66:20:@47601.4]
  wire  regs_420_io_enable; // @[RegFile.scala 66:20:@47601.4]
  wire  regs_421_clock; // @[RegFile.scala 66:20:@47615.4]
  wire  regs_421_reset; // @[RegFile.scala 66:20:@47615.4]
  wire [63:0] regs_421_io_in; // @[RegFile.scala 66:20:@47615.4]
  wire  regs_421_io_reset; // @[RegFile.scala 66:20:@47615.4]
  wire [63:0] regs_421_io_out; // @[RegFile.scala 66:20:@47615.4]
  wire  regs_421_io_enable; // @[RegFile.scala 66:20:@47615.4]
  wire  regs_422_clock; // @[RegFile.scala 66:20:@47629.4]
  wire  regs_422_reset; // @[RegFile.scala 66:20:@47629.4]
  wire [63:0] regs_422_io_in; // @[RegFile.scala 66:20:@47629.4]
  wire  regs_422_io_reset; // @[RegFile.scala 66:20:@47629.4]
  wire [63:0] regs_422_io_out; // @[RegFile.scala 66:20:@47629.4]
  wire  regs_422_io_enable; // @[RegFile.scala 66:20:@47629.4]
  wire  regs_423_clock; // @[RegFile.scala 66:20:@47643.4]
  wire  regs_423_reset; // @[RegFile.scala 66:20:@47643.4]
  wire [63:0] regs_423_io_in; // @[RegFile.scala 66:20:@47643.4]
  wire  regs_423_io_reset; // @[RegFile.scala 66:20:@47643.4]
  wire [63:0] regs_423_io_out; // @[RegFile.scala 66:20:@47643.4]
  wire  regs_423_io_enable; // @[RegFile.scala 66:20:@47643.4]
  wire  regs_424_clock; // @[RegFile.scala 66:20:@47657.4]
  wire  regs_424_reset; // @[RegFile.scala 66:20:@47657.4]
  wire [63:0] regs_424_io_in; // @[RegFile.scala 66:20:@47657.4]
  wire  regs_424_io_reset; // @[RegFile.scala 66:20:@47657.4]
  wire [63:0] regs_424_io_out; // @[RegFile.scala 66:20:@47657.4]
  wire  regs_424_io_enable; // @[RegFile.scala 66:20:@47657.4]
  wire  regs_425_clock; // @[RegFile.scala 66:20:@47671.4]
  wire  regs_425_reset; // @[RegFile.scala 66:20:@47671.4]
  wire [63:0] regs_425_io_in; // @[RegFile.scala 66:20:@47671.4]
  wire  regs_425_io_reset; // @[RegFile.scala 66:20:@47671.4]
  wire [63:0] regs_425_io_out; // @[RegFile.scala 66:20:@47671.4]
  wire  regs_425_io_enable; // @[RegFile.scala 66:20:@47671.4]
  wire  regs_426_clock; // @[RegFile.scala 66:20:@47685.4]
  wire  regs_426_reset; // @[RegFile.scala 66:20:@47685.4]
  wire [63:0] regs_426_io_in; // @[RegFile.scala 66:20:@47685.4]
  wire  regs_426_io_reset; // @[RegFile.scala 66:20:@47685.4]
  wire [63:0] regs_426_io_out; // @[RegFile.scala 66:20:@47685.4]
  wire  regs_426_io_enable; // @[RegFile.scala 66:20:@47685.4]
  wire  regs_427_clock; // @[RegFile.scala 66:20:@47699.4]
  wire  regs_427_reset; // @[RegFile.scala 66:20:@47699.4]
  wire [63:0] regs_427_io_in; // @[RegFile.scala 66:20:@47699.4]
  wire  regs_427_io_reset; // @[RegFile.scala 66:20:@47699.4]
  wire [63:0] regs_427_io_out; // @[RegFile.scala 66:20:@47699.4]
  wire  regs_427_io_enable; // @[RegFile.scala 66:20:@47699.4]
  wire  regs_428_clock; // @[RegFile.scala 66:20:@47713.4]
  wire  regs_428_reset; // @[RegFile.scala 66:20:@47713.4]
  wire [63:0] regs_428_io_in; // @[RegFile.scala 66:20:@47713.4]
  wire  regs_428_io_reset; // @[RegFile.scala 66:20:@47713.4]
  wire [63:0] regs_428_io_out; // @[RegFile.scala 66:20:@47713.4]
  wire  regs_428_io_enable; // @[RegFile.scala 66:20:@47713.4]
  wire  regs_429_clock; // @[RegFile.scala 66:20:@47727.4]
  wire  regs_429_reset; // @[RegFile.scala 66:20:@47727.4]
  wire [63:0] regs_429_io_in; // @[RegFile.scala 66:20:@47727.4]
  wire  regs_429_io_reset; // @[RegFile.scala 66:20:@47727.4]
  wire [63:0] regs_429_io_out; // @[RegFile.scala 66:20:@47727.4]
  wire  regs_429_io_enable; // @[RegFile.scala 66:20:@47727.4]
  wire  regs_430_clock; // @[RegFile.scala 66:20:@47741.4]
  wire  regs_430_reset; // @[RegFile.scala 66:20:@47741.4]
  wire [63:0] regs_430_io_in; // @[RegFile.scala 66:20:@47741.4]
  wire  regs_430_io_reset; // @[RegFile.scala 66:20:@47741.4]
  wire [63:0] regs_430_io_out; // @[RegFile.scala 66:20:@47741.4]
  wire  regs_430_io_enable; // @[RegFile.scala 66:20:@47741.4]
  wire  regs_431_clock; // @[RegFile.scala 66:20:@47755.4]
  wire  regs_431_reset; // @[RegFile.scala 66:20:@47755.4]
  wire [63:0] regs_431_io_in; // @[RegFile.scala 66:20:@47755.4]
  wire  regs_431_io_reset; // @[RegFile.scala 66:20:@47755.4]
  wire [63:0] regs_431_io_out; // @[RegFile.scala 66:20:@47755.4]
  wire  regs_431_io_enable; // @[RegFile.scala 66:20:@47755.4]
  wire  regs_432_clock; // @[RegFile.scala 66:20:@47769.4]
  wire  regs_432_reset; // @[RegFile.scala 66:20:@47769.4]
  wire [63:0] regs_432_io_in; // @[RegFile.scala 66:20:@47769.4]
  wire  regs_432_io_reset; // @[RegFile.scala 66:20:@47769.4]
  wire [63:0] regs_432_io_out; // @[RegFile.scala 66:20:@47769.4]
  wire  regs_432_io_enable; // @[RegFile.scala 66:20:@47769.4]
  wire  regs_433_clock; // @[RegFile.scala 66:20:@47783.4]
  wire  regs_433_reset; // @[RegFile.scala 66:20:@47783.4]
  wire [63:0] regs_433_io_in; // @[RegFile.scala 66:20:@47783.4]
  wire  regs_433_io_reset; // @[RegFile.scala 66:20:@47783.4]
  wire [63:0] regs_433_io_out; // @[RegFile.scala 66:20:@47783.4]
  wire  regs_433_io_enable; // @[RegFile.scala 66:20:@47783.4]
  wire  regs_434_clock; // @[RegFile.scala 66:20:@47797.4]
  wire  regs_434_reset; // @[RegFile.scala 66:20:@47797.4]
  wire [63:0] regs_434_io_in; // @[RegFile.scala 66:20:@47797.4]
  wire  regs_434_io_reset; // @[RegFile.scala 66:20:@47797.4]
  wire [63:0] regs_434_io_out; // @[RegFile.scala 66:20:@47797.4]
  wire  regs_434_io_enable; // @[RegFile.scala 66:20:@47797.4]
  wire  regs_435_clock; // @[RegFile.scala 66:20:@47811.4]
  wire  regs_435_reset; // @[RegFile.scala 66:20:@47811.4]
  wire [63:0] regs_435_io_in; // @[RegFile.scala 66:20:@47811.4]
  wire  regs_435_io_reset; // @[RegFile.scala 66:20:@47811.4]
  wire [63:0] regs_435_io_out; // @[RegFile.scala 66:20:@47811.4]
  wire  regs_435_io_enable; // @[RegFile.scala 66:20:@47811.4]
  wire  regs_436_clock; // @[RegFile.scala 66:20:@47825.4]
  wire  regs_436_reset; // @[RegFile.scala 66:20:@47825.4]
  wire [63:0] regs_436_io_in; // @[RegFile.scala 66:20:@47825.4]
  wire  regs_436_io_reset; // @[RegFile.scala 66:20:@47825.4]
  wire [63:0] regs_436_io_out; // @[RegFile.scala 66:20:@47825.4]
  wire  regs_436_io_enable; // @[RegFile.scala 66:20:@47825.4]
  wire  regs_437_clock; // @[RegFile.scala 66:20:@47839.4]
  wire  regs_437_reset; // @[RegFile.scala 66:20:@47839.4]
  wire [63:0] regs_437_io_in; // @[RegFile.scala 66:20:@47839.4]
  wire  regs_437_io_reset; // @[RegFile.scala 66:20:@47839.4]
  wire [63:0] regs_437_io_out; // @[RegFile.scala 66:20:@47839.4]
  wire  regs_437_io_enable; // @[RegFile.scala 66:20:@47839.4]
  wire  regs_438_clock; // @[RegFile.scala 66:20:@47853.4]
  wire  regs_438_reset; // @[RegFile.scala 66:20:@47853.4]
  wire [63:0] regs_438_io_in; // @[RegFile.scala 66:20:@47853.4]
  wire  regs_438_io_reset; // @[RegFile.scala 66:20:@47853.4]
  wire [63:0] regs_438_io_out; // @[RegFile.scala 66:20:@47853.4]
  wire  regs_438_io_enable; // @[RegFile.scala 66:20:@47853.4]
  wire  regs_439_clock; // @[RegFile.scala 66:20:@47867.4]
  wire  regs_439_reset; // @[RegFile.scala 66:20:@47867.4]
  wire [63:0] regs_439_io_in; // @[RegFile.scala 66:20:@47867.4]
  wire  regs_439_io_reset; // @[RegFile.scala 66:20:@47867.4]
  wire [63:0] regs_439_io_out; // @[RegFile.scala 66:20:@47867.4]
  wire  regs_439_io_enable; // @[RegFile.scala 66:20:@47867.4]
  wire  regs_440_clock; // @[RegFile.scala 66:20:@47881.4]
  wire  regs_440_reset; // @[RegFile.scala 66:20:@47881.4]
  wire [63:0] regs_440_io_in; // @[RegFile.scala 66:20:@47881.4]
  wire  regs_440_io_reset; // @[RegFile.scala 66:20:@47881.4]
  wire [63:0] regs_440_io_out; // @[RegFile.scala 66:20:@47881.4]
  wire  regs_440_io_enable; // @[RegFile.scala 66:20:@47881.4]
  wire  regs_441_clock; // @[RegFile.scala 66:20:@47895.4]
  wire  regs_441_reset; // @[RegFile.scala 66:20:@47895.4]
  wire [63:0] regs_441_io_in; // @[RegFile.scala 66:20:@47895.4]
  wire  regs_441_io_reset; // @[RegFile.scala 66:20:@47895.4]
  wire [63:0] regs_441_io_out; // @[RegFile.scala 66:20:@47895.4]
  wire  regs_441_io_enable; // @[RegFile.scala 66:20:@47895.4]
  wire  regs_442_clock; // @[RegFile.scala 66:20:@47909.4]
  wire  regs_442_reset; // @[RegFile.scala 66:20:@47909.4]
  wire [63:0] regs_442_io_in; // @[RegFile.scala 66:20:@47909.4]
  wire  regs_442_io_reset; // @[RegFile.scala 66:20:@47909.4]
  wire [63:0] regs_442_io_out; // @[RegFile.scala 66:20:@47909.4]
  wire  regs_442_io_enable; // @[RegFile.scala 66:20:@47909.4]
  wire  regs_443_clock; // @[RegFile.scala 66:20:@47923.4]
  wire  regs_443_reset; // @[RegFile.scala 66:20:@47923.4]
  wire [63:0] regs_443_io_in; // @[RegFile.scala 66:20:@47923.4]
  wire  regs_443_io_reset; // @[RegFile.scala 66:20:@47923.4]
  wire [63:0] regs_443_io_out; // @[RegFile.scala 66:20:@47923.4]
  wire  regs_443_io_enable; // @[RegFile.scala 66:20:@47923.4]
  wire  regs_444_clock; // @[RegFile.scala 66:20:@47937.4]
  wire  regs_444_reset; // @[RegFile.scala 66:20:@47937.4]
  wire [63:0] regs_444_io_in; // @[RegFile.scala 66:20:@47937.4]
  wire  regs_444_io_reset; // @[RegFile.scala 66:20:@47937.4]
  wire [63:0] regs_444_io_out; // @[RegFile.scala 66:20:@47937.4]
  wire  regs_444_io_enable; // @[RegFile.scala 66:20:@47937.4]
  wire  regs_445_clock; // @[RegFile.scala 66:20:@47951.4]
  wire  regs_445_reset; // @[RegFile.scala 66:20:@47951.4]
  wire [63:0] regs_445_io_in; // @[RegFile.scala 66:20:@47951.4]
  wire  regs_445_io_reset; // @[RegFile.scala 66:20:@47951.4]
  wire [63:0] regs_445_io_out; // @[RegFile.scala 66:20:@47951.4]
  wire  regs_445_io_enable; // @[RegFile.scala 66:20:@47951.4]
  wire  regs_446_clock; // @[RegFile.scala 66:20:@47965.4]
  wire  regs_446_reset; // @[RegFile.scala 66:20:@47965.4]
  wire [63:0] regs_446_io_in; // @[RegFile.scala 66:20:@47965.4]
  wire  regs_446_io_reset; // @[RegFile.scala 66:20:@47965.4]
  wire [63:0] regs_446_io_out; // @[RegFile.scala 66:20:@47965.4]
  wire  regs_446_io_enable; // @[RegFile.scala 66:20:@47965.4]
  wire  regs_447_clock; // @[RegFile.scala 66:20:@47979.4]
  wire  regs_447_reset; // @[RegFile.scala 66:20:@47979.4]
  wire [63:0] regs_447_io_in; // @[RegFile.scala 66:20:@47979.4]
  wire  regs_447_io_reset; // @[RegFile.scala 66:20:@47979.4]
  wire [63:0] regs_447_io_out; // @[RegFile.scala 66:20:@47979.4]
  wire  regs_447_io_enable; // @[RegFile.scala 66:20:@47979.4]
  wire  regs_448_clock; // @[RegFile.scala 66:20:@47993.4]
  wire  regs_448_reset; // @[RegFile.scala 66:20:@47993.4]
  wire [63:0] regs_448_io_in; // @[RegFile.scala 66:20:@47993.4]
  wire  regs_448_io_reset; // @[RegFile.scala 66:20:@47993.4]
  wire [63:0] regs_448_io_out; // @[RegFile.scala 66:20:@47993.4]
  wire  regs_448_io_enable; // @[RegFile.scala 66:20:@47993.4]
  wire  regs_449_clock; // @[RegFile.scala 66:20:@48007.4]
  wire  regs_449_reset; // @[RegFile.scala 66:20:@48007.4]
  wire [63:0] regs_449_io_in; // @[RegFile.scala 66:20:@48007.4]
  wire  regs_449_io_reset; // @[RegFile.scala 66:20:@48007.4]
  wire [63:0] regs_449_io_out; // @[RegFile.scala 66:20:@48007.4]
  wire  regs_449_io_enable; // @[RegFile.scala 66:20:@48007.4]
  wire  regs_450_clock; // @[RegFile.scala 66:20:@48021.4]
  wire  regs_450_reset; // @[RegFile.scala 66:20:@48021.4]
  wire [63:0] regs_450_io_in; // @[RegFile.scala 66:20:@48021.4]
  wire  regs_450_io_reset; // @[RegFile.scala 66:20:@48021.4]
  wire [63:0] regs_450_io_out; // @[RegFile.scala 66:20:@48021.4]
  wire  regs_450_io_enable; // @[RegFile.scala 66:20:@48021.4]
  wire  regs_451_clock; // @[RegFile.scala 66:20:@48035.4]
  wire  regs_451_reset; // @[RegFile.scala 66:20:@48035.4]
  wire [63:0] regs_451_io_in; // @[RegFile.scala 66:20:@48035.4]
  wire  regs_451_io_reset; // @[RegFile.scala 66:20:@48035.4]
  wire [63:0] regs_451_io_out; // @[RegFile.scala 66:20:@48035.4]
  wire  regs_451_io_enable; // @[RegFile.scala 66:20:@48035.4]
  wire  regs_452_clock; // @[RegFile.scala 66:20:@48049.4]
  wire  regs_452_reset; // @[RegFile.scala 66:20:@48049.4]
  wire [63:0] regs_452_io_in; // @[RegFile.scala 66:20:@48049.4]
  wire  regs_452_io_reset; // @[RegFile.scala 66:20:@48049.4]
  wire [63:0] regs_452_io_out; // @[RegFile.scala 66:20:@48049.4]
  wire  regs_452_io_enable; // @[RegFile.scala 66:20:@48049.4]
  wire  regs_453_clock; // @[RegFile.scala 66:20:@48063.4]
  wire  regs_453_reset; // @[RegFile.scala 66:20:@48063.4]
  wire [63:0] regs_453_io_in; // @[RegFile.scala 66:20:@48063.4]
  wire  regs_453_io_reset; // @[RegFile.scala 66:20:@48063.4]
  wire [63:0] regs_453_io_out; // @[RegFile.scala 66:20:@48063.4]
  wire  regs_453_io_enable; // @[RegFile.scala 66:20:@48063.4]
  wire  regs_454_clock; // @[RegFile.scala 66:20:@48077.4]
  wire  regs_454_reset; // @[RegFile.scala 66:20:@48077.4]
  wire [63:0] regs_454_io_in; // @[RegFile.scala 66:20:@48077.4]
  wire  regs_454_io_reset; // @[RegFile.scala 66:20:@48077.4]
  wire [63:0] regs_454_io_out; // @[RegFile.scala 66:20:@48077.4]
  wire  regs_454_io_enable; // @[RegFile.scala 66:20:@48077.4]
  wire  regs_455_clock; // @[RegFile.scala 66:20:@48091.4]
  wire  regs_455_reset; // @[RegFile.scala 66:20:@48091.4]
  wire [63:0] regs_455_io_in; // @[RegFile.scala 66:20:@48091.4]
  wire  regs_455_io_reset; // @[RegFile.scala 66:20:@48091.4]
  wire [63:0] regs_455_io_out; // @[RegFile.scala 66:20:@48091.4]
  wire  regs_455_io_enable; // @[RegFile.scala 66:20:@48091.4]
  wire  regs_456_clock; // @[RegFile.scala 66:20:@48105.4]
  wire  regs_456_reset; // @[RegFile.scala 66:20:@48105.4]
  wire [63:0] regs_456_io_in; // @[RegFile.scala 66:20:@48105.4]
  wire  regs_456_io_reset; // @[RegFile.scala 66:20:@48105.4]
  wire [63:0] regs_456_io_out; // @[RegFile.scala 66:20:@48105.4]
  wire  regs_456_io_enable; // @[RegFile.scala 66:20:@48105.4]
  wire  regs_457_clock; // @[RegFile.scala 66:20:@48119.4]
  wire  regs_457_reset; // @[RegFile.scala 66:20:@48119.4]
  wire [63:0] regs_457_io_in; // @[RegFile.scala 66:20:@48119.4]
  wire  regs_457_io_reset; // @[RegFile.scala 66:20:@48119.4]
  wire [63:0] regs_457_io_out; // @[RegFile.scala 66:20:@48119.4]
  wire  regs_457_io_enable; // @[RegFile.scala 66:20:@48119.4]
  wire  regs_458_clock; // @[RegFile.scala 66:20:@48133.4]
  wire  regs_458_reset; // @[RegFile.scala 66:20:@48133.4]
  wire [63:0] regs_458_io_in; // @[RegFile.scala 66:20:@48133.4]
  wire  regs_458_io_reset; // @[RegFile.scala 66:20:@48133.4]
  wire [63:0] regs_458_io_out; // @[RegFile.scala 66:20:@48133.4]
  wire  regs_458_io_enable; // @[RegFile.scala 66:20:@48133.4]
  wire  regs_459_clock; // @[RegFile.scala 66:20:@48147.4]
  wire  regs_459_reset; // @[RegFile.scala 66:20:@48147.4]
  wire [63:0] regs_459_io_in; // @[RegFile.scala 66:20:@48147.4]
  wire  regs_459_io_reset; // @[RegFile.scala 66:20:@48147.4]
  wire [63:0] regs_459_io_out; // @[RegFile.scala 66:20:@48147.4]
  wire  regs_459_io_enable; // @[RegFile.scala 66:20:@48147.4]
  wire  regs_460_clock; // @[RegFile.scala 66:20:@48161.4]
  wire  regs_460_reset; // @[RegFile.scala 66:20:@48161.4]
  wire [63:0] regs_460_io_in; // @[RegFile.scala 66:20:@48161.4]
  wire  regs_460_io_reset; // @[RegFile.scala 66:20:@48161.4]
  wire [63:0] regs_460_io_out; // @[RegFile.scala 66:20:@48161.4]
  wire  regs_460_io_enable; // @[RegFile.scala 66:20:@48161.4]
  wire  regs_461_clock; // @[RegFile.scala 66:20:@48175.4]
  wire  regs_461_reset; // @[RegFile.scala 66:20:@48175.4]
  wire [63:0] regs_461_io_in; // @[RegFile.scala 66:20:@48175.4]
  wire  regs_461_io_reset; // @[RegFile.scala 66:20:@48175.4]
  wire [63:0] regs_461_io_out; // @[RegFile.scala 66:20:@48175.4]
  wire  regs_461_io_enable; // @[RegFile.scala 66:20:@48175.4]
  wire  regs_462_clock; // @[RegFile.scala 66:20:@48189.4]
  wire  regs_462_reset; // @[RegFile.scala 66:20:@48189.4]
  wire [63:0] regs_462_io_in; // @[RegFile.scala 66:20:@48189.4]
  wire  regs_462_io_reset; // @[RegFile.scala 66:20:@48189.4]
  wire [63:0] regs_462_io_out; // @[RegFile.scala 66:20:@48189.4]
  wire  regs_462_io_enable; // @[RegFile.scala 66:20:@48189.4]
  wire  regs_463_clock; // @[RegFile.scala 66:20:@48203.4]
  wire  regs_463_reset; // @[RegFile.scala 66:20:@48203.4]
  wire [63:0] regs_463_io_in; // @[RegFile.scala 66:20:@48203.4]
  wire  regs_463_io_reset; // @[RegFile.scala 66:20:@48203.4]
  wire [63:0] regs_463_io_out; // @[RegFile.scala 66:20:@48203.4]
  wire  regs_463_io_enable; // @[RegFile.scala 66:20:@48203.4]
  wire  regs_464_clock; // @[RegFile.scala 66:20:@48217.4]
  wire  regs_464_reset; // @[RegFile.scala 66:20:@48217.4]
  wire [63:0] regs_464_io_in; // @[RegFile.scala 66:20:@48217.4]
  wire  regs_464_io_reset; // @[RegFile.scala 66:20:@48217.4]
  wire [63:0] regs_464_io_out; // @[RegFile.scala 66:20:@48217.4]
  wire  regs_464_io_enable; // @[RegFile.scala 66:20:@48217.4]
  wire  regs_465_clock; // @[RegFile.scala 66:20:@48231.4]
  wire  regs_465_reset; // @[RegFile.scala 66:20:@48231.4]
  wire [63:0] regs_465_io_in; // @[RegFile.scala 66:20:@48231.4]
  wire  regs_465_io_reset; // @[RegFile.scala 66:20:@48231.4]
  wire [63:0] regs_465_io_out; // @[RegFile.scala 66:20:@48231.4]
  wire  regs_465_io_enable; // @[RegFile.scala 66:20:@48231.4]
  wire  regs_466_clock; // @[RegFile.scala 66:20:@48245.4]
  wire  regs_466_reset; // @[RegFile.scala 66:20:@48245.4]
  wire [63:0] regs_466_io_in; // @[RegFile.scala 66:20:@48245.4]
  wire  regs_466_io_reset; // @[RegFile.scala 66:20:@48245.4]
  wire [63:0] regs_466_io_out; // @[RegFile.scala 66:20:@48245.4]
  wire  regs_466_io_enable; // @[RegFile.scala 66:20:@48245.4]
  wire  regs_467_clock; // @[RegFile.scala 66:20:@48259.4]
  wire  regs_467_reset; // @[RegFile.scala 66:20:@48259.4]
  wire [63:0] regs_467_io_in; // @[RegFile.scala 66:20:@48259.4]
  wire  regs_467_io_reset; // @[RegFile.scala 66:20:@48259.4]
  wire [63:0] regs_467_io_out; // @[RegFile.scala 66:20:@48259.4]
  wire  regs_467_io_enable; // @[RegFile.scala 66:20:@48259.4]
  wire  regs_468_clock; // @[RegFile.scala 66:20:@48273.4]
  wire  regs_468_reset; // @[RegFile.scala 66:20:@48273.4]
  wire [63:0] regs_468_io_in; // @[RegFile.scala 66:20:@48273.4]
  wire  regs_468_io_reset; // @[RegFile.scala 66:20:@48273.4]
  wire [63:0] regs_468_io_out; // @[RegFile.scala 66:20:@48273.4]
  wire  regs_468_io_enable; // @[RegFile.scala 66:20:@48273.4]
  wire  regs_469_clock; // @[RegFile.scala 66:20:@48287.4]
  wire  regs_469_reset; // @[RegFile.scala 66:20:@48287.4]
  wire [63:0] regs_469_io_in; // @[RegFile.scala 66:20:@48287.4]
  wire  regs_469_io_reset; // @[RegFile.scala 66:20:@48287.4]
  wire [63:0] regs_469_io_out; // @[RegFile.scala 66:20:@48287.4]
  wire  regs_469_io_enable; // @[RegFile.scala 66:20:@48287.4]
  wire  regs_470_clock; // @[RegFile.scala 66:20:@48301.4]
  wire  regs_470_reset; // @[RegFile.scala 66:20:@48301.4]
  wire [63:0] regs_470_io_in; // @[RegFile.scala 66:20:@48301.4]
  wire  regs_470_io_reset; // @[RegFile.scala 66:20:@48301.4]
  wire [63:0] regs_470_io_out; // @[RegFile.scala 66:20:@48301.4]
  wire  regs_470_io_enable; // @[RegFile.scala 66:20:@48301.4]
  wire  regs_471_clock; // @[RegFile.scala 66:20:@48315.4]
  wire  regs_471_reset; // @[RegFile.scala 66:20:@48315.4]
  wire [63:0] regs_471_io_in; // @[RegFile.scala 66:20:@48315.4]
  wire  regs_471_io_reset; // @[RegFile.scala 66:20:@48315.4]
  wire [63:0] regs_471_io_out; // @[RegFile.scala 66:20:@48315.4]
  wire  regs_471_io_enable; // @[RegFile.scala 66:20:@48315.4]
  wire  regs_472_clock; // @[RegFile.scala 66:20:@48329.4]
  wire  regs_472_reset; // @[RegFile.scala 66:20:@48329.4]
  wire [63:0] regs_472_io_in; // @[RegFile.scala 66:20:@48329.4]
  wire  regs_472_io_reset; // @[RegFile.scala 66:20:@48329.4]
  wire [63:0] regs_472_io_out; // @[RegFile.scala 66:20:@48329.4]
  wire  regs_472_io_enable; // @[RegFile.scala 66:20:@48329.4]
  wire  regs_473_clock; // @[RegFile.scala 66:20:@48343.4]
  wire  regs_473_reset; // @[RegFile.scala 66:20:@48343.4]
  wire [63:0] regs_473_io_in; // @[RegFile.scala 66:20:@48343.4]
  wire  regs_473_io_reset; // @[RegFile.scala 66:20:@48343.4]
  wire [63:0] regs_473_io_out; // @[RegFile.scala 66:20:@48343.4]
  wire  regs_473_io_enable; // @[RegFile.scala 66:20:@48343.4]
  wire  regs_474_clock; // @[RegFile.scala 66:20:@48357.4]
  wire  regs_474_reset; // @[RegFile.scala 66:20:@48357.4]
  wire [63:0] regs_474_io_in; // @[RegFile.scala 66:20:@48357.4]
  wire  regs_474_io_reset; // @[RegFile.scala 66:20:@48357.4]
  wire [63:0] regs_474_io_out; // @[RegFile.scala 66:20:@48357.4]
  wire  regs_474_io_enable; // @[RegFile.scala 66:20:@48357.4]
  wire  regs_475_clock; // @[RegFile.scala 66:20:@48371.4]
  wire  regs_475_reset; // @[RegFile.scala 66:20:@48371.4]
  wire [63:0] regs_475_io_in; // @[RegFile.scala 66:20:@48371.4]
  wire  regs_475_io_reset; // @[RegFile.scala 66:20:@48371.4]
  wire [63:0] regs_475_io_out; // @[RegFile.scala 66:20:@48371.4]
  wire  regs_475_io_enable; // @[RegFile.scala 66:20:@48371.4]
  wire  regs_476_clock; // @[RegFile.scala 66:20:@48385.4]
  wire  regs_476_reset; // @[RegFile.scala 66:20:@48385.4]
  wire [63:0] regs_476_io_in; // @[RegFile.scala 66:20:@48385.4]
  wire  regs_476_io_reset; // @[RegFile.scala 66:20:@48385.4]
  wire [63:0] regs_476_io_out; // @[RegFile.scala 66:20:@48385.4]
  wire  regs_476_io_enable; // @[RegFile.scala 66:20:@48385.4]
  wire  regs_477_clock; // @[RegFile.scala 66:20:@48399.4]
  wire  regs_477_reset; // @[RegFile.scala 66:20:@48399.4]
  wire [63:0] regs_477_io_in; // @[RegFile.scala 66:20:@48399.4]
  wire  regs_477_io_reset; // @[RegFile.scala 66:20:@48399.4]
  wire [63:0] regs_477_io_out; // @[RegFile.scala 66:20:@48399.4]
  wire  regs_477_io_enable; // @[RegFile.scala 66:20:@48399.4]
  wire  regs_478_clock; // @[RegFile.scala 66:20:@48413.4]
  wire  regs_478_reset; // @[RegFile.scala 66:20:@48413.4]
  wire [63:0] regs_478_io_in; // @[RegFile.scala 66:20:@48413.4]
  wire  regs_478_io_reset; // @[RegFile.scala 66:20:@48413.4]
  wire [63:0] regs_478_io_out; // @[RegFile.scala 66:20:@48413.4]
  wire  regs_478_io_enable; // @[RegFile.scala 66:20:@48413.4]
  wire  regs_479_clock; // @[RegFile.scala 66:20:@48427.4]
  wire  regs_479_reset; // @[RegFile.scala 66:20:@48427.4]
  wire [63:0] regs_479_io_in; // @[RegFile.scala 66:20:@48427.4]
  wire  regs_479_io_reset; // @[RegFile.scala 66:20:@48427.4]
  wire [63:0] regs_479_io_out; // @[RegFile.scala 66:20:@48427.4]
  wire  regs_479_io_enable; // @[RegFile.scala 66:20:@48427.4]
  wire  regs_480_clock; // @[RegFile.scala 66:20:@48441.4]
  wire  regs_480_reset; // @[RegFile.scala 66:20:@48441.4]
  wire [63:0] regs_480_io_in; // @[RegFile.scala 66:20:@48441.4]
  wire  regs_480_io_reset; // @[RegFile.scala 66:20:@48441.4]
  wire [63:0] regs_480_io_out; // @[RegFile.scala 66:20:@48441.4]
  wire  regs_480_io_enable; // @[RegFile.scala 66:20:@48441.4]
  wire  regs_481_clock; // @[RegFile.scala 66:20:@48455.4]
  wire  regs_481_reset; // @[RegFile.scala 66:20:@48455.4]
  wire [63:0] regs_481_io_in; // @[RegFile.scala 66:20:@48455.4]
  wire  regs_481_io_reset; // @[RegFile.scala 66:20:@48455.4]
  wire [63:0] regs_481_io_out; // @[RegFile.scala 66:20:@48455.4]
  wire  regs_481_io_enable; // @[RegFile.scala 66:20:@48455.4]
  wire  regs_482_clock; // @[RegFile.scala 66:20:@48469.4]
  wire  regs_482_reset; // @[RegFile.scala 66:20:@48469.4]
  wire [63:0] regs_482_io_in; // @[RegFile.scala 66:20:@48469.4]
  wire  regs_482_io_reset; // @[RegFile.scala 66:20:@48469.4]
  wire [63:0] regs_482_io_out; // @[RegFile.scala 66:20:@48469.4]
  wire  regs_482_io_enable; // @[RegFile.scala 66:20:@48469.4]
  wire  regs_483_clock; // @[RegFile.scala 66:20:@48483.4]
  wire  regs_483_reset; // @[RegFile.scala 66:20:@48483.4]
  wire [63:0] regs_483_io_in; // @[RegFile.scala 66:20:@48483.4]
  wire  regs_483_io_reset; // @[RegFile.scala 66:20:@48483.4]
  wire [63:0] regs_483_io_out; // @[RegFile.scala 66:20:@48483.4]
  wire  regs_483_io_enable; // @[RegFile.scala 66:20:@48483.4]
  wire  regs_484_clock; // @[RegFile.scala 66:20:@48497.4]
  wire  regs_484_reset; // @[RegFile.scala 66:20:@48497.4]
  wire [63:0] regs_484_io_in; // @[RegFile.scala 66:20:@48497.4]
  wire  regs_484_io_reset; // @[RegFile.scala 66:20:@48497.4]
  wire [63:0] regs_484_io_out; // @[RegFile.scala 66:20:@48497.4]
  wire  regs_484_io_enable; // @[RegFile.scala 66:20:@48497.4]
  wire  regs_485_clock; // @[RegFile.scala 66:20:@48511.4]
  wire  regs_485_reset; // @[RegFile.scala 66:20:@48511.4]
  wire [63:0] regs_485_io_in; // @[RegFile.scala 66:20:@48511.4]
  wire  regs_485_io_reset; // @[RegFile.scala 66:20:@48511.4]
  wire [63:0] regs_485_io_out; // @[RegFile.scala 66:20:@48511.4]
  wire  regs_485_io_enable; // @[RegFile.scala 66:20:@48511.4]
  wire  regs_486_clock; // @[RegFile.scala 66:20:@48525.4]
  wire  regs_486_reset; // @[RegFile.scala 66:20:@48525.4]
  wire [63:0] regs_486_io_in; // @[RegFile.scala 66:20:@48525.4]
  wire  regs_486_io_reset; // @[RegFile.scala 66:20:@48525.4]
  wire [63:0] regs_486_io_out; // @[RegFile.scala 66:20:@48525.4]
  wire  regs_486_io_enable; // @[RegFile.scala 66:20:@48525.4]
  wire  regs_487_clock; // @[RegFile.scala 66:20:@48539.4]
  wire  regs_487_reset; // @[RegFile.scala 66:20:@48539.4]
  wire [63:0] regs_487_io_in; // @[RegFile.scala 66:20:@48539.4]
  wire  regs_487_io_reset; // @[RegFile.scala 66:20:@48539.4]
  wire [63:0] regs_487_io_out; // @[RegFile.scala 66:20:@48539.4]
  wire  regs_487_io_enable; // @[RegFile.scala 66:20:@48539.4]
  wire  regs_488_clock; // @[RegFile.scala 66:20:@48553.4]
  wire  regs_488_reset; // @[RegFile.scala 66:20:@48553.4]
  wire [63:0] regs_488_io_in; // @[RegFile.scala 66:20:@48553.4]
  wire  regs_488_io_reset; // @[RegFile.scala 66:20:@48553.4]
  wire [63:0] regs_488_io_out; // @[RegFile.scala 66:20:@48553.4]
  wire  regs_488_io_enable; // @[RegFile.scala 66:20:@48553.4]
  wire  regs_489_clock; // @[RegFile.scala 66:20:@48567.4]
  wire  regs_489_reset; // @[RegFile.scala 66:20:@48567.4]
  wire [63:0] regs_489_io_in; // @[RegFile.scala 66:20:@48567.4]
  wire  regs_489_io_reset; // @[RegFile.scala 66:20:@48567.4]
  wire [63:0] regs_489_io_out; // @[RegFile.scala 66:20:@48567.4]
  wire  regs_489_io_enable; // @[RegFile.scala 66:20:@48567.4]
  wire  regs_490_clock; // @[RegFile.scala 66:20:@48581.4]
  wire  regs_490_reset; // @[RegFile.scala 66:20:@48581.4]
  wire [63:0] regs_490_io_in; // @[RegFile.scala 66:20:@48581.4]
  wire  regs_490_io_reset; // @[RegFile.scala 66:20:@48581.4]
  wire [63:0] regs_490_io_out; // @[RegFile.scala 66:20:@48581.4]
  wire  regs_490_io_enable; // @[RegFile.scala 66:20:@48581.4]
  wire  regs_491_clock; // @[RegFile.scala 66:20:@48595.4]
  wire  regs_491_reset; // @[RegFile.scala 66:20:@48595.4]
  wire [63:0] regs_491_io_in; // @[RegFile.scala 66:20:@48595.4]
  wire  regs_491_io_reset; // @[RegFile.scala 66:20:@48595.4]
  wire [63:0] regs_491_io_out; // @[RegFile.scala 66:20:@48595.4]
  wire  regs_491_io_enable; // @[RegFile.scala 66:20:@48595.4]
  wire  regs_492_clock; // @[RegFile.scala 66:20:@48609.4]
  wire  regs_492_reset; // @[RegFile.scala 66:20:@48609.4]
  wire [63:0] regs_492_io_in; // @[RegFile.scala 66:20:@48609.4]
  wire  regs_492_io_reset; // @[RegFile.scala 66:20:@48609.4]
  wire [63:0] regs_492_io_out; // @[RegFile.scala 66:20:@48609.4]
  wire  regs_492_io_enable; // @[RegFile.scala 66:20:@48609.4]
  wire  regs_493_clock; // @[RegFile.scala 66:20:@48623.4]
  wire  regs_493_reset; // @[RegFile.scala 66:20:@48623.4]
  wire [63:0] regs_493_io_in; // @[RegFile.scala 66:20:@48623.4]
  wire  regs_493_io_reset; // @[RegFile.scala 66:20:@48623.4]
  wire [63:0] regs_493_io_out; // @[RegFile.scala 66:20:@48623.4]
  wire  regs_493_io_enable; // @[RegFile.scala 66:20:@48623.4]
  wire  regs_494_clock; // @[RegFile.scala 66:20:@48637.4]
  wire  regs_494_reset; // @[RegFile.scala 66:20:@48637.4]
  wire [63:0] regs_494_io_in; // @[RegFile.scala 66:20:@48637.4]
  wire  regs_494_io_reset; // @[RegFile.scala 66:20:@48637.4]
  wire [63:0] regs_494_io_out; // @[RegFile.scala 66:20:@48637.4]
  wire  regs_494_io_enable; // @[RegFile.scala 66:20:@48637.4]
  wire  regs_495_clock; // @[RegFile.scala 66:20:@48651.4]
  wire  regs_495_reset; // @[RegFile.scala 66:20:@48651.4]
  wire [63:0] regs_495_io_in; // @[RegFile.scala 66:20:@48651.4]
  wire  regs_495_io_reset; // @[RegFile.scala 66:20:@48651.4]
  wire [63:0] regs_495_io_out; // @[RegFile.scala 66:20:@48651.4]
  wire  regs_495_io_enable; // @[RegFile.scala 66:20:@48651.4]
  wire  regs_496_clock; // @[RegFile.scala 66:20:@48665.4]
  wire  regs_496_reset; // @[RegFile.scala 66:20:@48665.4]
  wire [63:0] regs_496_io_in; // @[RegFile.scala 66:20:@48665.4]
  wire  regs_496_io_reset; // @[RegFile.scala 66:20:@48665.4]
  wire [63:0] regs_496_io_out; // @[RegFile.scala 66:20:@48665.4]
  wire  regs_496_io_enable; // @[RegFile.scala 66:20:@48665.4]
  wire  regs_497_clock; // @[RegFile.scala 66:20:@48679.4]
  wire  regs_497_reset; // @[RegFile.scala 66:20:@48679.4]
  wire [63:0] regs_497_io_in; // @[RegFile.scala 66:20:@48679.4]
  wire  regs_497_io_reset; // @[RegFile.scala 66:20:@48679.4]
  wire [63:0] regs_497_io_out; // @[RegFile.scala 66:20:@48679.4]
  wire  regs_497_io_enable; // @[RegFile.scala 66:20:@48679.4]
  wire  regs_498_clock; // @[RegFile.scala 66:20:@48693.4]
  wire  regs_498_reset; // @[RegFile.scala 66:20:@48693.4]
  wire [63:0] regs_498_io_in; // @[RegFile.scala 66:20:@48693.4]
  wire  regs_498_io_reset; // @[RegFile.scala 66:20:@48693.4]
  wire [63:0] regs_498_io_out; // @[RegFile.scala 66:20:@48693.4]
  wire  regs_498_io_enable; // @[RegFile.scala 66:20:@48693.4]
  wire  regs_499_clock; // @[RegFile.scala 66:20:@48707.4]
  wire  regs_499_reset; // @[RegFile.scala 66:20:@48707.4]
  wire [63:0] regs_499_io_in; // @[RegFile.scala 66:20:@48707.4]
  wire  regs_499_io_reset; // @[RegFile.scala 66:20:@48707.4]
  wire [63:0] regs_499_io_out; // @[RegFile.scala 66:20:@48707.4]
  wire  regs_499_io_enable; // @[RegFile.scala 66:20:@48707.4]
  wire  regs_500_clock; // @[RegFile.scala 66:20:@48721.4]
  wire  regs_500_reset; // @[RegFile.scala 66:20:@48721.4]
  wire [63:0] regs_500_io_in; // @[RegFile.scala 66:20:@48721.4]
  wire  regs_500_io_reset; // @[RegFile.scala 66:20:@48721.4]
  wire [63:0] regs_500_io_out; // @[RegFile.scala 66:20:@48721.4]
  wire  regs_500_io_enable; // @[RegFile.scala 66:20:@48721.4]
  wire  regs_501_clock; // @[RegFile.scala 66:20:@48735.4]
  wire  regs_501_reset; // @[RegFile.scala 66:20:@48735.4]
  wire [63:0] regs_501_io_in; // @[RegFile.scala 66:20:@48735.4]
  wire  regs_501_io_reset; // @[RegFile.scala 66:20:@48735.4]
  wire [63:0] regs_501_io_out; // @[RegFile.scala 66:20:@48735.4]
  wire  regs_501_io_enable; // @[RegFile.scala 66:20:@48735.4]
  wire  regs_502_clock; // @[RegFile.scala 66:20:@48749.4]
  wire  regs_502_reset; // @[RegFile.scala 66:20:@48749.4]
  wire [63:0] regs_502_io_in; // @[RegFile.scala 66:20:@48749.4]
  wire  regs_502_io_reset; // @[RegFile.scala 66:20:@48749.4]
  wire [63:0] regs_502_io_out; // @[RegFile.scala 66:20:@48749.4]
  wire  regs_502_io_enable; // @[RegFile.scala 66:20:@48749.4]
  wire  regs_503_clock; // @[RegFile.scala 66:20:@48763.4]
  wire  regs_503_reset; // @[RegFile.scala 66:20:@48763.4]
  wire [63:0] regs_503_io_in; // @[RegFile.scala 66:20:@48763.4]
  wire  regs_503_io_reset; // @[RegFile.scala 66:20:@48763.4]
  wire [63:0] regs_503_io_out; // @[RegFile.scala 66:20:@48763.4]
  wire  regs_503_io_enable; // @[RegFile.scala 66:20:@48763.4]
  wire  regs_504_clock; // @[RegFile.scala 66:20:@48777.4]
  wire  regs_504_reset; // @[RegFile.scala 66:20:@48777.4]
  wire [63:0] regs_504_io_in; // @[RegFile.scala 66:20:@48777.4]
  wire  regs_504_io_reset; // @[RegFile.scala 66:20:@48777.4]
  wire [63:0] regs_504_io_out; // @[RegFile.scala 66:20:@48777.4]
  wire  regs_504_io_enable; // @[RegFile.scala 66:20:@48777.4]
  wire  regs_505_clock; // @[RegFile.scala 66:20:@48791.4]
  wire  regs_505_reset; // @[RegFile.scala 66:20:@48791.4]
  wire [63:0] regs_505_io_in; // @[RegFile.scala 66:20:@48791.4]
  wire  regs_505_io_reset; // @[RegFile.scala 66:20:@48791.4]
  wire [63:0] regs_505_io_out; // @[RegFile.scala 66:20:@48791.4]
  wire  regs_505_io_enable; // @[RegFile.scala 66:20:@48791.4]
  wire  regs_506_clock; // @[RegFile.scala 66:20:@48805.4]
  wire  regs_506_reset; // @[RegFile.scala 66:20:@48805.4]
  wire [63:0] regs_506_io_in; // @[RegFile.scala 66:20:@48805.4]
  wire  regs_506_io_reset; // @[RegFile.scala 66:20:@48805.4]
  wire [63:0] regs_506_io_out; // @[RegFile.scala 66:20:@48805.4]
  wire  regs_506_io_enable; // @[RegFile.scala 66:20:@48805.4]
  wire  regs_507_clock; // @[RegFile.scala 66:20:@48819.4]
  wire  regs_507_reset; // @[RegFile.scala 66:20:@48819.4]
  wire [63:0] regs_507_io_in; // @[RegFile.scala 66:20:@48819.4]
  wire  regs_507_io_reset; // @[RegFile.scala 66:20:@48819.4]
  wire [63:0] regs_507_io_out; // @[RegFile.scala 66:20:@48819.4]
  wire  regs_507_io_enable; // @[RegFile.scala 66:20:@48819.4]
  wire  regs_508_clock; // @[RegFile.scala 66:20:@48833.4]
  wire  regs_508_reset; // @[RegFile.scala 66:20:@48833.4]
  wire [63:0] regs_508_io_in; // @[RegFile.scala 66:20:@48833.4]
  wire  regs_508_io_reset; // @[RegFile.scala 66:20:@48833.4]
  wire [63:0] regs_508_io_out; // @[RegFile.scala 66:20:@48833.4]
  wire  regs_508_io_enable; // @[RegFile.scala 66:20:@48833.4]
  wire  regs_509_clock; // @[RegFile.scala 66:20:@48847.4]
  wire  regs_509_reset; // @[RegFile.scala 66:20:@48847.4]
  wire [63:0] regs_509_io_in; // @[RegFile.scala 66:20:@48847.4]
  wire  regs_509_io_reset; // @[RegFile.scala 66:20:@48847.4]
  wire [63:0] regs_509_io_out; // @[RegFile.scala 66:20:@48847.4]
  wire  regs_509_io_enable; // @[RegFile.scala 66:20:@48847.4]
  wire  regs_510_clock; // @[RegFile.scala 66:20:@48861.4]
  wire  regs_510_reset; // @[RegFile.scala 66:20:@48861.4]
  wire [63:0] regs_510_io_in; // @[RegFile.scala 66:20:@48861.4]
  wire  regs_510_io_reset; // @[RegFile.scala 66:20:@48861.4]
  wire [63:0] regs_510_io_out; // @[RegFile.scala 66:20:@48861.4]
  wire  regs_510_io_enable; // @[RegFile.scala 66:20:@48861.4]
  wire  regs_511_clock; // @[RegFile.scala 66:20:@48875.4]
  wire  regs_511_reset; // @[RegFile.scala 66:20:@48875.4]
  wire [63:0] regs_511_io_in; // @[RegFile.scala 66:20:@48875.4]
  wire  regs_511_io_reset; // @[RegFile.scala 66:20:@48875.4]
  wire [63:0] regs_511_io_out; // @[RegFile.scala 66:20:@48875.4]
  wire  regs_511_io_enable; // @[RegFile.scala 66:20:@48875.4]
  wire  regs_512_clock; // @[RegFile.scala 66:20:@48889.4]
  wire  regs_512_reset; // @[RegFile.scala 66:20:@48889.4]
  wire [63:0] regs_512_io_in; // @[RegFile.scala 66:20:@48889.4]
  wire  regs_512_io_reset; // @[RegFile.scala 66:20:@48889.4]
  wire [63:0] regs_512_io_out; // @[RegFile.scala 66:20:@48889.4]
  wire  regs_512_io_enable; // @[RegFile.scala 66:20:@48889.4]
  wire  regs_513_clock; // @[RegFile.scala 66:20:@48903.4]
  wire  regs_513_reset; // @[RegFile.scala 66:20:@48903.4]
  wire [63:0] regs_513_io_in; // @[RegFile.scala 66:20:@48903.4]
  wire  regs_513_io_reset; // @[RegFile.scala 66:20:@48903.4]
  wire [63:0] regs_513_io_out; // @[RegFile.scala 66:20:@48903.4]
  wire  regs_513_io_enable; // @[RegFile.scala 66:20:@48903.4]
  wire  regs_514_clock; // @[RegFile.scala 66:20:@48917.4]
  wire  regs_514_reset; // @[RegFile.scala 66:20:@48917.4]
  wire [63:0] regs_514_io_in; // @[RegFile.scala 66:20:@48917.4]
  wire  regs_514_io_reset; // @[RegFile.scala 66:20:@48917.4]
  wire [63:0] regs_514_io_out; // @[RegFile.scala 66:20:@48917.4]
  wire  regs_514_io_enable; // @[RegFile.scala 66:20:@48917.4]
  wire  regs_515_clock; // @[RegFile.scala 66:20:@48931.4]
  wire  regs_515_reset; // @[RegFile.scala 66:20:@48931.4]
  wire [63:0] regs_515_io_in; // @[RegFile.scala 66:20:@48931.4]
  wire  regs_515_io_reset; // @[RegFile.scala 66:20:@48931.4]
  wire [63:0] regs_515_io_out; // @[RegFile.scala 66:20:@48931.4]
  wire  regs_515_io_enable; // @[RegFile.scala 66:20:@48931.4]
  wire  regs_516_clock; // @[RegFile.scala 66:20:@48945.4]
  wire  regs_516_reset; // @[RegFile.scala 66:20:@48945.4]
  wire [63:0] regs_516_io_in; // @[RegFile.scala 66:20:@48945.4]
  wire  regs_516_io_reset; // @[RegFile.scala 66:20:@48945.4]
  wire [63:0] regs_516_io_out; // @[RegFile.scala 66:20:@48945.4]
  wire  regs_516_io_enable; // @[RegFile.scala 66:20:@48945.4]
  wire  regs_517_clock; // @[RegFile.scala 66:20:@48959.4]
  wire  regs_517_reset; // @[RegFile.scala 66:20:@48959.4]
  wire [63:0] regs_517_io_in; // @[RegFile.scala 66:20:@48959.4]
  wire  regs_517_io_reset; // @[RegFile.scala 66:20:@48959.4]
  wire [63:0] regs_517_io_out; // @[RegFile.scala 66:20:@48959.4]
  wire  regs_517_io_enable; // @[RegFile.scala 66:20:@48959.4]
  wire  regs_518_clock; // @[RegFile.scala 66:20:@48973.4]
  wire  regs_518_reset; // @[RegFile.scala 66:20:@48973.4]
  wire [63:0] regs_518_io_in; // @[RegFile.scala 66:20:@48973.4]
  wire  regs_518_io_reset; // @[RegFile.scala 66:20:@48973.4]
  wire [63:0] regs_518_io_out; // @[RegFile.scala 66:20:@48973.4]
  wire  regs_518_io_enable; // @[RegFile.scala 66:20:@48973.4]
  wire  regs_519_clock; // @[RegFile.scala 66:20:@48987.4]
  wire  regs_519_reset; // @[RegFile.scala 66:20:@48987.4]
  wire [63:0] regs_519_io_in; // @[RegFile.scala 66:20:@48987.4]
  wire  regs_519_io_reset; // @[RegFile.scala 66:20:@48987.4]
  wire [63:0] regs_519_io_out; // @[RegFile.scala 66:20:@48987.4]
  wire  regs_519_io_enable; // @[RegFile.scala 66:20:@48987.4]
  wire  regs_520_clock; // @[RegFile.scala 66:20:@49001.4]
  wire  regs_520_reset; // @[RegFile.scala 66:20:@49001.4]
  wire [63:0] regs_520_io_in; // @[RegFile.scala 66:20:@49001.4]
  wire  regs_520_io_reset; // @[RegFile.scala 66:20:@49001.4]
  wire [63:0] regs_520_io_out; // @[RegFile.scala 66:20:@49001.4]
  wire  regs_520_io_enable; // @[RegFile.scala 66:20:@49001.4]
  wire  regs_521_clock; // @[RegFile.scala 66:20:@49015.4]
  wire  regs_521_reset; // @[RegFile.scala 66:20:@49015.4]
  wire [63:0] regs_521_io_in; // @[RegFile.scala 66:20:@49015.4]
  wire  regs_521_io_reset; // @[RegFile.scala 66:20:@49015.4]
  wire [63:0] regs_521_io_out; // @[RegFile.scala 66:20:@49015.4]
  wire  regs_521_io_enable; // @[RegFile.scala 66:20:@49015.4]
  wire  regs_522_clock; // @[RegFile.scala 66:20:@49029.4]
  wire  regs_522_reset; // @[RegFile.scala 66:20:@49029.4]
  wire [63:0] regs_522_io_in; // @[RegFile.scala 66:20:@49029.4]
  wire  regs_522_io_reset; // @[RegFile.scala 66:20:@49029.4]
  wire [63:0] regs_522_io_out; // @[RegFile.scala 66:20:@49029.4]
  wire  regs_522_io_enable; // @[RegFile.scala 66:20:@49029.4]
  wire  regs_523_clock; // @[RegFile.scala 66:20:@49043.4]
  wire  regs_523_reset; // @[RegFile.scala 66:20:@49043.4]
  wire [63:0] regs_523_io_in; // @[RegFile.scala 66:20:@49043.4]
  wire  regs_523_io_reset; // @[RegFile.scala 66:20:@49043.4]
  wire [63:0] regs_523_io_out; // @[RegFile.scala 66:20:@49043.4]
  wire  regs_523_io_enable; // @[RegFile.scala 66:20:@49043.4]
  wire  regs_524_clock; // @[RegFile.scala 66:20:@49057.4]
  wire  regs_524_reset; // @[RegFile.scala 66:20:@49057.4]
  wire [63:0] regs_524_io_in; // @[RegFile.scala 66:20:@49057.4]
  wire  regs_524_io_reset; // @[RegFile.scala 66:20:@49057.4]
  wire [63:0] regs_524_io_out; // @[RegFile.scala 66:20:@49057.4]
  wire  regs_524_io_enable; // @[RegFile.scala 66:20:@49057.4]
  wire  regs_525_clock; // @[RegFile.scala 66:20:@49071.4]
  wire  regs_525_reset; // @[RegFile.scala 66:20:@49071.4]
  wire [63:0] regs_525_io_in; // @[RegFile.scala 66:20:@49071.4]
  wire  regs_525_io_reset; // @[RegFile.scala 66:20:@49071.4]
  wire [63:0] regs_525_io_out; // @[RegFile.scala 66:20:@49071.4]
  wire  regs_525_io_enable; // @[RegFile.scala 66:20:@49071.4]
  wire  regs_526_clock; // @[RegFile.scala 66:20:@49085.4]
  wire  regs_526_reset; // @[RegFile.scala 66:20:@49085.4]
  wire [63:0] regs_526_io_in; // @[RegFile.scala 66:20:@49085.4]
  wire  regs_526_io_reset; // @[RegFile.scala 66:20:@49085.4]
  wire [63:0] regs_526_io_out; // @[RegFile.scala 66:20:@49085.4]
  wire  regs_526_io_enable; // @[RegFile.scala 66:20:@49085.4]
  wire  regs_527_clock; // @[RegFile.scala 66:20:@49099.4]
  wire  regs_527_reset; // @[RegFile.scala 66:20:@49099.4]
  wire [63:0] regs_527_io_in; // @[RegFile.scala 66:20:@49099.4]
  wire  regs_527_io_reset; // @[RegFile.scala 66:20:@49099.4]
  wire [63:0] regs_527_io_out; // @[RegFile.scala 66:20:@49099.4]
  wire  regs_527_io_enable; // @[RegFile.scala 66:20:@49099.4]
  wire  regs_528_clock; // @[RegFile.scala 66:20:@49113.4]
  wire  regs_528_reset; // @[RegFile.scala 66:20:@49113.4]
  wire [63:0] regs_528_io_in; // @[RegFile.scala 66:20:@49113.4]
  wire  regs_528_io_reset; // @[RegFile.scala 66:20:@49113.4]
  wire [63:0] regs_528_io_out; // @[RegFile.scala 66:20:@49113.4]
  wire  regs_528_io_enable; // @[RegFile.scala 66:20:@49113.4]
  wire  regs_529_clock; // @[RegFile.scala 66:20:@49127.4]
  wire  regs_529_reset; // @[RegFile.scala 66:20:@49127.4]
  wire [63:0] regs_529_io_in; // @[RegFile.scala 66:20:@49127.4]
  wire  regs_529_io_reset; // @[RegFile.scala 66:20:@49127.4]
  wire [63:0] regs_529_io_out; // @[RegFile.scala 66:20:@49127.4]
  wire  regs_529_io_enable; // @[RegFile.scala 66:20:@49127.4]
  wire  regs_530_clock; // @[RegFile.scala 66:20:@49141.4]
  wire  regs_530_reset; // @[RegFile.scala 66:20:@49141.4]
  wire [63:0] regs_530_io_in; // @[RegFile.scala 66:20:@49141.4]
  wire  regs_530_io_reset; // @[RegFile.scala 66:20:@49141.4]
  wire [63:0] regs_530_io_out; // @[RegFile.scala 66:20:@49141.4]
  wire  regs_530_io_enable; // @[RegFile.scala 66:20:@49141.4]
  wire  regs_531_clock; // @[RegFile.scala 66:20:@49155.4]
  wire  regs_531_reset; // @[RegFile.scala 66:20:@49155.4]
  wire [63:0] regs_531_io_in; // @[RegFile.scala 66:20:@49155.4]
  wire  regs_531_io_reset; // @[RegFile.scala 66:20:@49155.4]
  wire [63:0] regs_531_io_out; // @[RegFile.scala 66:20:@49155.4]
  wire  regs_531_io_enable; // @[RegFile.scala 66:20:@49155.4]
  wire  regs_532_clock; // @[RegFile.scala 66:20:@49169.4]
  wire  regs_532_reset; // @[RegFile.scala 66:20:@49169.4]
  wire [63:0] regs_532_io_in; // @[RegFile.scala 66:20:@49169.4]
  wire  regs_532_io_reset; // @[RegFile.scala 66:20:@49169.4]
  wire [63:0] regs_532_io_out; // @[RegFile.scala 66:20:@49169.4]
  wire  regs_532_io_enable; // @[RegFile.scala 66:20:@49169.4]
  wire  regs_533_clock; // @[RegFile.scala 66:20:@49183.4]
  wire  regs_533_reset; // @[RegFile.scala 66:20:@49183.4]
  wire [63:0] regs_533_io_in; // @[RegFile.scala 66:20:@49183.4]
  wire  regs_533_io_reset; // @[RegFile.scala 66:20:@49183.4]
  wire [63:0] regs_533_io_out; // @[RegFile.scala 66:20:@49183.4]
  wire  regs_533_io_enable; // @[RegFile.scala 66:20:@49183.4]
  wire [63:0] rport_io_ins_0; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_1; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_2; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_3; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_4; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_5; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_6; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_7; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_8; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_9; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_10; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_11; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_12; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_13; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_14; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_15; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_16; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_17; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_18; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_19; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_20; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_21; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_22; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_23; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_24; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_25; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_26; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_27; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_28; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_29; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_30; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_31; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_32; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_33; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_34; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_35; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_36; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_37; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_38; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_39; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_40; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_41; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_42; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_43; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_44; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_45; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_46; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_47; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_48; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_49; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_50; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_51; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_52; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_53; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_54; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_55; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_56; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_57; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_58; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_59; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_60; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_61; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_62; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_63; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_64; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_65; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_66; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_67; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_68; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_69; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_70; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_71; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_72; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_73; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_74; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_75; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_76; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_77; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_78; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_79; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_80; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_81; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_82; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_83; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_84; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_85; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_86; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_87; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_88; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_89; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_90; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_91; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_92; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_93; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_94; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_95; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_96; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_97; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_98; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_99; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_100; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_101; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_102; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_103; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_104; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_105; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_106; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_107; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_108; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_109; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_110; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_111; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_112; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_113; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_114; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_115; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_116; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_117; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_118; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_119; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_120; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_121; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_122; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_123; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_124; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_125; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_126; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_127; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_128; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_129; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_130; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_131; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_132; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_133; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_134; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_135; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_136; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_137; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_138; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_139; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_140; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_141; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_142; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_143; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_144; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_145; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_146; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_147; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_148; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_149; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_150; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_151; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_152; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_153; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_154; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_155; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_156; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_157; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_158; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_159; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_160; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_161; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_162; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_163; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_164; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_165; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_166; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_167; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_168; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_169; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_170; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_171; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_172; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_173; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_174; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_175; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_176; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_177; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_178; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_179; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_180; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_181; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_182; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_183; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_184; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_185; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_186; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_187; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_188; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_189; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_190; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_191; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_192; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_193; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_194; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_195; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_196; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_197; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_198; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_199; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_200; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_201; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_202; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_203; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_204; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_205; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_206; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_207; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_208; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_209; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_210; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_211; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_212; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_213; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_214; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_215; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_216; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_217; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_218; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_219; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_220; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_221; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_222; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_223; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_224; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_225; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_226; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_227; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_228; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_229; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_230; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_231; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_232; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_233; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_234; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_235; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_236; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_237; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_238; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_239; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_240; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_241; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_242; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_243; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_244; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_245; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_246; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_247; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_248; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_249; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_250; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_251; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_252; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_253; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_254; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_255; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_256; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_257; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_258; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_259; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_260; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_261; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_262; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_263; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_264; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_265; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_266; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_267; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_268; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_269; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_270; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_271; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_272; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_273; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_274; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_275; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_276; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_277; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_278; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_279; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_280; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_281; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_282; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_283; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_284; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_285; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_286; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_287; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_288; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_289; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_290; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_291; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_292; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_293; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_294; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_295; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_296; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_297; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_298; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_299; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_300; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_301; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_302; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_303; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_304; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_305; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_306; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_307; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_308; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_309; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_310; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_311; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_312; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_313; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_314; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_315; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_316; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_317; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_318; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_319; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_320; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_321; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_322; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_323; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_324; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_325; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_326; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_327; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_328; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_329; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_330; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_331; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_332; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_333; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_334; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_335; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_336; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_337; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_338; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_339; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_340; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_341; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_342; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_343; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_344; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_345; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_346; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_347; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_348; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_349; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_350; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_351; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_352; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_353; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_354; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_355; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_356; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_357; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_358; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_359; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_360; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_361; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_362; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_363; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_364; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_365; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_366; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_367; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_368; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_369; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_370; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_371; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_372; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_373; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_374; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_375; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_376; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_377; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_378; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_379; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_380; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_381; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_382; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_383; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_384; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_385; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_386; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_387; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_388; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_389; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_390; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_391; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_392; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_393; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_394; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_395; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_396; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_397; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_398; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_399; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_400; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_401; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_402; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_403; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_404; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_405; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_406; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_407; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_408; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_409; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_410; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_411; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_412; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_413; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_414; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_415; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_416; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_417; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_418; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_419; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_420; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_421; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_422; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_423; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_424; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_425; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_426; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_427; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_428; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_429; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_430; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_431; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_432; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_433; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_434; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_435; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_436; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_437; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_438; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_439; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_440; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_441; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_442; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_443; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_444; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_445; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_446; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_447; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_448; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_449; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_450; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_451; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_452; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_453; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_454; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_455; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_456; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_457; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_458; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_459; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_460; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_461; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_462; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_463; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_464; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_465; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_466; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_467; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_468; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_469; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_470; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_471; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_472; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_473; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_474; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_475; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_476; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_477; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_478; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_479; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_480; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_481; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_482; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_483; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_484; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_485; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_486; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_487; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_488; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_489; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_490; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_491; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_492; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_493; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_494; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_495; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_496; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_497; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_498; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_499; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_500; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_501; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_502; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_503; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_504; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_505; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_506; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_507; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_508; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_509; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_510; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_511; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_512; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_513; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_514; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_515; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_516; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_517; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_518; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_519; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_520; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_521; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_522; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_523; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_524; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_525; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_526; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_527; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_528; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_529; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_530; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_531; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_532; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_ins_533; // @[RegFile.scala 95:21:@49197.4]
  wire [9:0] rport_io_sel; // @[RegFile.scala 95:21:@49197.4]
  wire [63:0] rport_io_out; // @[RegFile.scala 95:21:@49197.4]
  wire  _T_3262; // @[RegFile.scala 80:42:@41723.4]
  wire  _T_3268; // @[RegFile.scala 68:46:@41735.4]
  wire  _T_3269; // @[RegFile.scala 68:34:@41736.4]
  wire  _T_3282; // @[RegFile.scala 80:42:@41754.4]
  wire  _T_3288; // @[RegFile.scala 74:80:@41766.4]
  wire  _T_3289; // @[RegFile.scala 74:68:@41767.4]
  wire  _T_3295; // @[RegFile.scala 74:80:@41780.4]
  wire  _T_3296; // @[RegFile.scala 74:68:@41781.4]
  wire  _T_3302; // @[RegFile.scala 74:80:@41794.4]
  wire  _T_3303; // @[RegFile.scala 74:68:@41795.4]
  wire  _T_3309; // @[RegFile.scala 74:80:@41808.4]
  wire  _T_3310; // @[RegFile.scala 74:68:@41809.4]
  wire  _T_3316; // @[RegFile.scala 74:80:@41822.4]
  wire  _T_3317; // @[RegFile.scala 74:68:@41823.4]
  wire  _T_3323; // @[RegFile.scala 74:80:@41836.4]
  wire  _T_3324; // @[RegFile.scala 74:68:@41837.4]
  wire  _T_3330; // @[RegFile.scala 74:80:@41850.4]
  wire  _T_3331; // @[RegFile.scala 74:68:@41851.4]
  wire  _T_3337; // @[RegFile.scala 74:80:@41864.4]
  wire  _T_3338; // @[RegFile.scala 74:68:@41865.4]
  wire  _T_3344; // @[RegFile.scala 74:80:@41878.4]
  wire  _T_3345; // @[RegFile.scala 74:68:@41879.4]
  wire  _T_3351; // @[RegFile.scala 74:80:@41892.4]
  wire  _T_3352; // @[RegFile.scala 74:68:@41893.4]
  wire  _T_3358; // @[RegFile.scala 74:80:@41906.4]
  wire  _T_3359; // @[RegFile.scala 74:68:@41907.4]
  wire  _T_3365; // @[RegFile.scala 74:80:@41920.4]
  wire  _T_3366; // @[RegFile.scala 74:68:@41921.4]
  wire  _T_3372; // @[RegFile.scala 74:80:@41934.4]
  wire  _T_3373; // @[RegFile.scala 74:68:@41935.4]
  wire  _T_3379; // @[RegFile.scala 74:80:@41948.4]
  wire  _T_3380; // @[RegFile.scala 74:68:@41949.4]
  wire  _T_3386; // @[RegFile.scala 74:80:@41962.4]
  wire  _T_3387; // @[RegFile.scala 74:68:@41963.4]
  wire  _T_3393; // @[RegFile.scala 74:80:@41976.4]
  wire  _T_3394; // @[RegFile.scala 74:68:@41977.4]
  wire  _T_3400; // @[RegFile.scala 74:80:@41990.4]
  wire  _T_3401; // @[RegFile.scala 74:68:@41991.4]
  wire  _T_3407; // @[RegFile.scala 74:80:@42004.4]
  wire  _T_3408; // @[RegFile.scala 74:68:@42005.4]
  wire  _T_3414; // @[RegFile.scala 74:80:@42018.4]
  wire  _T_3415; // @[RegFile.scala 74:68:@42019.4]
  wire  _T_3421; // @[RegFile.scala 74:80:@42032.4]
  wire  _T_3422; // @[RegFile.scala 74:68:@42033.4]
  wire  _T_3428; // @[RegFile.scala 74:80:@42046.4]
  wire  _T_3429; // @[RegFile.scala 74:68:@42047.4]
  wire  _T_3435; // @[RegFile.scala 74:80:@42060.4]
  wire  _T_3436; // @[RegFile.scala 74:68:@42061.4]
  wire  _T_3442; // @[RegFile.scala 74:80:@42074.4]
  wire  _T_3443; // @[RegFile.scala 74:68:@42075.4]
  wire  _T_3449; // @[RegFile.scala 74:80:@42088.4]
  wire  _T_3450; // @[RegFile.scala 74:68:@42089.4]
  wire  _T_3456; // @[RegFile.scala 74:80:@42102.4]
  wire  _T_3457; // @[RegFile.scala 74:68:@42103.4]
  wire  _T_3463; // @[RegFile.scala 74:80:@42116.4]
  wire  _T_3464; // @[RegFile.scala 74:68:@42117.4]
  wire  _T_3470; // @[RegFile.scala 74:80:@42130.4]
  wire  _T_3471; // @[RegFile.scala 74:68:@42131.4]
  wire  _T_3477; // @[RegFile.scala 74:80:@42144.4]
  wire  _T_3478; // @[RegFile.scala 74:68:@42145.4]
  wire  _T_3484; // @[RegFile.scala 74:80:@42158.4]
  wire  _T_3485; // @[RegFile.scala 74:68:@42159.4]
  wire  _T_3491; // @[RegFile.scala 74:80:@42172.4]
  wire  _T_3492; // @[RegFile.scala 74:68:@42173.4]
  wire  _T_3498; // @[RegFile.scala 74:80:@42186.4]
  wire  _T_3499; // @[RegFile.scala 74:68:@42187.4]
  wire  _T_3505; // @[RegFile.scala 74:80:@42200.4]
  wire  _T_3506; // @[RegFile.scala 74:68:@42201.4]
  FringeFF regs_0 ( // @[RegFile.scala 66:20:@41720.4]
    .clock(regs_0_clock),
    .reset(regs_0_reset),
    .io_in(regs_0_io_in),
    .io_reset(regs_0_io_reset),
    .io_out(regs_0_io_out),
    .io_enable(regs_0_io_enable)
  );
  FringeFF regs_1 ( // @[RegFile.scala 66:20:@41732.4]
    .clock(regs_1_clock),
    .reset(regs_1_reset),
    .io_in(regs_1_io_in),
    .io_reset(regs_1_io_reset),
    .io_out(regs_1_io_out),
    .io_enable(regs_1_io_enable)
  );
  FringeFF regs_2 ( // @[RegFile.scala 66:20:@41751.4]
    .clock(regs_2_clock),
    .reset(regs_2_reset),
    .io_in(regs_2_io_in),
    .io_reset(regs_2_io_reset),
    .io_out(regs_2_io_out),
    .io_enable(regs_2_io_enable)
  );
  FringeFF regs_3 ( // @[RegFile.scala 66:20:@41763.4]
    .clock(regs_3_clock),
    .reset(regs_3_reset),
    .io_in(regs_3_io_in),
    .io_reset(regs_3_io_reset),
    .io_out(regs_3_io_out),
    .io_enable(regs_3_io_enable)
  );
  FringeFF regs_4 ( // @[RegFile.scala 66:20:@41777.4]
    .clock(regs_4_clock),
    .reset(regs_4_reset),
    .io_in(regs_4_io_in),
    .io_reset(regs_4_io_reset),
    .io_out(regs_4_io_out),
    .io_enable(regs_4_io_enable)
  );
  FringeFF regs_5 ( // @[RegFile.scala 66:20:@41791.4]
    .clock(regs_5_clock),
    .reset(regs_5_reset),
    .io_in(regs_5_io_in),
    .io_reset(regs_5_io_reset),
    .io_out(regs_5_io_out),
    .io_enable(regs_5_io_enable)
  );
  FringeFF regs_6 ( // @[RegFile.scala 66:20:@41805.4]
    .clock(regs_6_clock),
    .reset(regs_6_reset),
    .io_in(regs_6_io_in),
    .io_reset(regs_6_io_reset),
    .io_out(regs_6_io_out),
    .io_enable(regs_6_io_enable)
  );
  FringeFF regs_7 ( // @[RegFile.scala 66:20:@41819.4]
    .clock(regs_7_clock),
    .reset(regs_7_reset),
    .io_in(regs_7_io_in),
    .io_reset(regs_7_io_reset),
    .io_out(regs_7_io_out),
    .io_enable(regs_7_io_enable)
  );
  FringeFF regs_8 ( // @[RegFile.scala 66:20:@41833.4]
    .clock(regs_8_clock),
    .reset(regs_8_reset),
    .io_in(regs_8_io_in),
    .io_reset(regs_8_io_reset),
    .io_out(regs_8_io_out),
    .io_enable(regs_8_io_enable)
  );
  FringeFF regs_9 ( // @[RegFile.scala 66:20:@41847.4]
    .clock(regs_9_clock),
    .reset(regs_9_reset),
    .io_in(regs_9_io_in),
    .io_reset(regs_9_io_reset),
    .io_out(regs_9_io_out),
    .io_enable(regs_9_io_enable)
  );
  FringeFF regs_10 ( // @[RegFile.scala 66:20:@41861.4]
    .clock(regs_10_clock),
    .reset(regs_10_reset),
    .io_in(regs_10_io_in),
    .io_reset(regs_10_io_reset),
    .io_out(regs_10_io_out),
    .io_enable(regs_10_io_enable)
  );
  FringeFF regs_11 ( // @[RegFile.scala 66:20:@41875.4]
    .clock(regs_11_clock),
    .reset(regs_11_reset),
    .io_in(regs_11_io_in),
    .io_reset(regs_11_io_reset),
    .io_out(regs_11_io_out),
    .io_enable(regs_11_io_enable)
  );
  FringeFF regs_12 ( // @[RegFile.scala 66:20:@41889.4]
    .clock(regs_12_clock),
    .reset(regs_12_reset),
    .io_in(regs_12_io_in),
    .io_reset(regs_12_io_reset),
    .io_out(regs_12_io_out),
    .io_enable(regs_12_io_enable)
  );
  FringeFF regs_13 ( // @[RegFile.scala 66:20:@41903.4]
    .clock(regs_13_clock),
    .reset(regs_13_reset),
    .io_in(regs_13_io_in),
    .io_reset(regs_13_io_reset),
    .io_out(regs_13_io_out),
    .io_enable(regs_13_io_enable)
  );
  FringeFF regs_14 ( // @[RegFile.scala 66:20:@41917.4]
    .clock(regs_14_clock),
    .reset(regs_14_reset),
    .io_in(regs_14_io_in),
    .io_reset(regs_14_io_reset),
    .io_out(regs_14_io_out),
    .io_enable(regs_14_io_enable)
  );
  FringeFF regs_15 ( // @[RegFile.scala 66:20:@41931.4]
    .clock(regs_15_clock),
    .reset(regs_15_reset),
    .io_in(regs_15_io_in),
    .io_reset(regs_15_io_reset),
    .io_out(regs_15_io_out),
    .io_enable(regs_15_io_enable)
  );
  FringeFF regs_16 ( // @[RegFile.scala 66:20:@41945.4]
    .clock(regs_16_clock),
    .reset(regs_16_reset),
    .io_in(regs_16_io_in),
    .io_reset(regs_16_io_reset),
    .io_out(regs_16_io_out),
    .io_enable(regs_16_io_enable)
  );
  FringeFF regs_17 ( // @[RegFile.scala 66:20:@41959.4]
    .clock(regs_17_clock),
    .reset(regs_17_reset),
    .io_in(regs_17_io_in),
    .io_reset(regs_17_io_reset),
    .io_out(regs_17_io_out),
    .io_enable(regs_17_io_enable)
  );
  FringeFF regs_18 ( // @[RegFile.scala 66:20:@41973.4]
    .clock(regs_18_clock),
    .reset(regs_18_reset),
    .io_in(regs_18_io_in),
    .io_reset(regs_18_io_reset),
    .io_out(regs_18_io_out),
    .io_enable(regs_18_io_enable)
  );
  FringeFF regs_19 ( // @[RegFile.scala 66:20:@41987.4]
    .clock(regs_19_clock),
    .reset(regs_19_reset),
    .io_in(regs_19_io_in),
    .io_reset(regs_19_io_reset),
    .io_out(regs_19_io_out),
    .io_enable(regs_19_io_enable)
  );
  FringeFF regs_20 ( // @[RegFile.scala 66:20:@42001.4]
    .clock(regs_20_clock),
    .reset(regs_20_reset),
    .io_in(regs_20_io_in),
    .io_reset(regs_20_io_reset),
    .io_out(regs_20_io_out),
    .io_enable(regs_20_io_enable)
  );
  FringeFF regs_21 ( // @[RegFile.scala 66:20:@42015.4]
    .clock(regs_21_clock),
    .reset(regs_21_reset),
    .io_in(regs_21_io_in),
    .io_reset(regs_21_io_reset),
    .io_out(regs_21_io_out),
    .io_enable(regs_21_io_enable)
  );
  FringeFF regs_22 ( // @[RegFile.scala 66:20:@42029.4]
    .clock(regs_22_clock),
    .reset(regs_22_reset),
    .io_in(regs_22_io_in),
    .io_reset(regs_22_io_reset),
    .io_out(regs_22_io_out),
    .io_enable(regs_22_io_enable)
  );
  FringeFF regs_23 ( // @[RegFile.scala 66:20:@42043.4]
    .clock(regs_23_clock),
    .reset(regs_23_reset),
    .io_in(regs_23_io_in),
    .io_reset(regs_23_io_reset),
    .io_out(regs_23_io_out),
    .io_enable(regs_23_io_enable)
  );
  FringeFF regs_24 ( // @[RegFile.scala 66:20:@42057.4]
    .clock(regs_24_clock),
    .reset(regs_24_reset),
    .io_in(regs_24_io_in),
    .io_reset(regs_24_io_reset),
    .io_out(regs_24_io_out),
    .io_enable(regs_24_io_enable)
  );
  FringeFF regs_25 ( // @[RegFile.scala 66:20:@42071.4]
    .clock(regs_25_clock),
    .reset(regs_25_reset),
    .io_in(regs_25_io_in),
    .io_reset(regs_25_io_reset),
    .io_out(regs_25_io_out),
    .io_enable(regs_25_io_enable)
  );
  FringeFF regs_26 ( // @[RegFile.scala 66:20:@42085.4]
    .clock(regs_26_clock),
    .reset(regs_26_reset),
    .io_in(regs_26_io_in),
    .io_reset(regs_26_io_reset),
    .io_out(regs_26_io_out),
    .io_enable(regs_26_io_enable)
  );
  FringeFF regs_27 ( // @[RegFile.scala 66:20:@42099.4]
    .clock(regs_27_clock),
    .reset(regs_27_reset),
    .io_in(regs_27_io_in),
    .io_reset(regs_27_io_reset),
    .io_out(regs_27_io_out),
    .io_enable(regs_27_io_enable)
  );
  FringeFF regs_28 ( // @[RegFile.scala 66:20:@42113.4]
    .clock(regs_28_clock),
    .reset(regs_28_reset),
    .io_in(regs_28_io_in),
    .io_reset(regs_28_io_reset),
    .io_out(regs_28_io_out),
    .io_enable(regs_28_io_enable)
  );
  FringeFF regs_29 ( // @[RegFile.scala 66:20:@42127.4]
    .clock(regs_29_clock),
    .reset(regs_29_reset),
    .io_in(regs_29_io_in),
    .io_reset(regs_29_io_reset),
    .io_out(regs_29_io_out),
    .io_enable(regs_29_io_enable)
  );
  FringeFF regs_30 ( // @[RegFile.scala 66:20:@42141.4]
    .clock(regs_30_clock),
    .reset(regs_30_reset),
    .io_in(regs_30_io_in),
    .io_reset(regs_30_io_reset),
    .io_out(regs_30_io_out),
    .io_enable(regs_30_io_enable)
  );
  FringeFF regs_31 ( // @[RegFile.scala 66:20:@42155.4]
    .clock(regs_31_clock),
    .reset(regs_31_reset),
    .io_in(regs_31_io_in),
    .io_reset(regs_31_io_reset),
    .io_out(regs_31_io_out),
    .io_enable(regs_31_io_enable)
  );
  FringeFF regs_32 ( // @[RegFile.scala 66:20:@42169.4]
    .clock(regs_32_clock),
    .reset(regs_32_reset),
    .io_in(regs_32_io_in),
    .io_reset(regs_32_io_reset),
    .io_out(regs_32_io_out),
    .io_enable(regs_32_io_enable)
  );
  FringeFF regs_33 ( // @[RegFile.scala 66:20:@42183.4]
    .clock(regs_33_clock),
    .reset(regs_33_reset),
    .io_in(regs_33_io_in),
    .io_reset(regs_33_io_reset),
    .io_out(regs_33_io_out),
    .io_enable(regs_33_io_enable)
  );
  FringeFF regs_34 ( // @[RegFile.scala 66:20:@42197.4]
    .clock(regs_34_clock),
    .reset(regs_34_reset),
    .io_in(regs_34_io_in),
    .io_reset(regs_34_io_reset),
    .io_out(regs_34_io_out),
    .io_enable(regs_34_io_enable)
  );
  FringeFF regs_35 ( // @[RegFile.scala 66:20:@42211.4]
    .clock(regs_35_clock),
    .reset(regs_35_reset),
    .io_in(regs_35_io_in),
    .io_reset(regs_35_io_reset),
    .io_out(regs_35_io_out),
    .io_enable(regs_35_io_enable)
  );
  FringeFF regs_36 ( // @[RegFile.scala 66:20:@42225.4]
    .clock(regs_36_clock),
    .reset(regs_36_reset),
    .io_in(regs_36_io_in),
    .io_reset(regs_36_io_reset),
    .io_out(regs_36_io_out),
    .io_enable(regs_36_io_enable)
  );
  FringeFF regs_37 ( // @[RegFile.scala 66:20:@42239.4]
    .clock(regs_37_clock),
    .reset(regs_37_reset),
    .io_in(regs_37_io_in),
    .io_reset(regs_37_io_reset),
    .io_out(regs_37_io_out),
    .io_enable(regs_37_io_enable)
  );
  FringeFF regs_38 ( // @[RegFile.scala 66:20:@42253.4]
    .clock(regs_38_clock),
    .reset(regs_38_reset),
    .io_in(regs_38_io_in),
    .io_reset(regs_38_io_reset),
    .io_out(regs_38_io_out),
    .io_enable(regs_38_io_enable)
  );
  FringeFF regs_39 ( // @[RegFile.scala 66:20:@42267.4]
    .clock(regs_39_clock),
    .reset(regs_39_reset),
    .io_in(regs_39_io_in),
    .io_reset(regs_39_io_reset),
    .io_out(regs_39_io_out),
    .io_enable(regs_39_io_enable)
  );
  FringeFF regs_40 ( // @[RegFile.scala 66:20:@42281.4]
    .clock(regs_40_clock),
    .reset(regs_40_reset),
    .io_in(regs_40_io_in),
    .io_reset(regs_40_io_reset),
    .io_out(regs_40_io_out),
    .io_enable(regs_40_io_enable)
  );
  FringeFF regs_41 ( // @[RegFile.scala 66:20:@42295.4]
    .clock(regs_41_clock),
    .reset(regs_41_reset),
    .io_in(regs_41_io_in),
    .io_reset(regs_41_io_reset),
    .io_out(regs_41_io_out),
    .io_enable(regs_41_io_enable)
  );
  FringeFF regs_42 ( // @[RegFile.scala 66:20:@42309.4]
    .clock(regs_42_clock),
    .reset(regs_42_reset),
    .io_in(regs_42_io_in),
    .io_reset(regs_42_io_reset),
    .io_out(regs_42_io_out),
    .io_enable(regs_42_io_enable)
  );
  FringeFF regs_43 ( // @[RegFile.scala 66:20:@42323.4]
    .clock(regs_43_clock),
    .reset(regs_43_reset),
    .io_in(regs_43_io_in),
    .io_reset(regs_43_io_reset),
    .io_out(regs_43_io_out),
    .io_enable(regs_43_io_enable)
  );
  FringeFF regs_44 ( // @[RegFile.scala 66:20:@42337.4]
    .clock(regs_44_clock),
    .reset(regs_44_reset),
    .io_in(regs_44_io_in),
    .io_reset(regs_44_io_reset),
    .io_out(regs_44_io_out),
    .io_enable(regs_44_io_enable)
  );
  FringeFF regs_45 ( // @[RegFile.scala 66:20:@42351.4]
    .clock(regs_45_clock),
    .reset(regs_45_reset),
    .io_in(regs_45_io_in),
    .io_reset(regs_45_io_reset),
    .io_out(regs_45_io_out),
    .io_enable(regs_45_io_enable)
  );
  FringeFF regs_46 ( // @[RegFile.scala 66:20:@42365.4]
    .clock(regs_46_clock),
    .reset(regs_46_reset),
    .io_in(regs_46_io_in),
    .io_reset(regs_46_io_reset),
    .io_out(regs_46_io_out),
    .io_enable(regs_46_io_enable)
  );
  FringeFF regs_47 ( // @[RegFile.scala 66:20:@42379.4]
    .clock(regs_47_clock),
    .reset(regs_47_reset),
    .io_in(regs_47_io_in),
    .io_reset(regs_47_io_reset),
    .io_out(regs_47_io_out),
    .io_enable(regs_47_io_enable)
  );
  FringeFF regs_48 ( // @[RegFile.scala 66:20:@42393.4]
    .clock(regs_48_clock),
    .reset(regs_48_reset),
    .io_in(regs_48_io_in),
    .io_reset(regs_48_io_reset),
    .io_out(regs_48_io_out),
    .io_enable(regs_48_io_enable)
  );
  FringeFF regs_49 ( // @[RegFile.scala 66:20:@42407.4]
    .clock(regs_49_clock),
    .reset(regs_49_reset),
    .io_in(regs_49_io_in),
    .io_reset(regs_49_io_reset),
    .io_out(regs_49_io_out),
    .io_enable(regs_49_io_enable)
  );
  FringeFF regs_50 ( // @[RegFile.scala 66:20:@42421.4]
    .clock(regs_50_clock),
    .reset(regs_50_reset),
    .io_in(regs_50_io_in),
    .io_reset(regs_50_io_reset),
    .io_out(regs_50_io_out),
    .io_enable(regs_50_io_enable)
  );
  FringeFF regs_51 ( // @[RegFile.scala 66:20:@42435.4]
    .clock(regs_51_clock),
    .reset(regs_51_reset),
    .io_in(regs_51_io_in),
    .io_reset(regs_51_io_reset),
    .io_out(regs_51_io_out),
    .io_enable(regs_51_io_enable)
  );
  FringeFF regs_52 ( // @[RegFile.scala 66:20:@42449.4]
    .clock(regs_52_clock),
    .reset(regs_52_reset),
    .io_in(regs_52_io_in),
    .io_reset(regs_52_io_reset),
    .io_out(regs_52_io_out),
    .io_enable(regs_52_io_enable)
  );
  FringeFF regs_53 ( // @[RegFile.scala 66:20:@42463.4]
    .clock(regs_53_clock),
    .reset(regs_53_reset),
    .io_in(regs_53_io_in),
    .io_reset(regs_53_io_reset),
    .io_out(regs_53_io_out),
    .io_enable(regs_53_io_enable)
  );
  FringeFF regs_54 ( // @[RegFile.scala 66:20:@42477.4]
    .clock(regs_54_clock),
    .reset(regs_54_reset),
    .io_in(regs_54_io_in),
    .io_reset(regs_54_io_reset),
    .io_out(regs_54_io_out),
    .io_enable(regs_54_io_enable)
  );
  FringeFF regs_55 ( // @[RegFile.scala 66:20:@42491.4]
    .clock(regs_55_clock),
    .reset(regs_55_reset),
    .io_in(regs_55_io_in),
    .io_reset(regs_55_io_reset),
    .io_out(regs_55_io_out),
    .io_enable(regs_55_io_enable)
  );
  FringeFF regs_56 ( // @[RegFile.scala 66:20:@42505.4]
    .clock(regs_56_clock),
    .reset(regs_56_reset),
    .io_in(regs_56_io_in),
    .io_reset(regs_56_io_reset),
    .io_out(regs_56_io_out),
    .io_enable(regs_56_io_enable)
  );
  FringeFF regs_57 ( // @[RegFile.scala 66:20:@42519.4]
    .clock(regs_57_clock),
    .reset(regs_57_reset),
    .io_in(regs_57_io_in),
    .io_reset(regs_57_io_reset),
    .io_out(regs_57_io_out),
    .io_enable(regs_57_io_enable)
  );
  FringeFF regs_58 ( // @[RegFile.scala 66:20:@42533.4]
    .clock(regs_58_clock),
    .reset(regs_58_reset),
    .io_in(regs_58_io_in),
    .io_reset(regs_58_io_reset),
    .io_out(regs_58_io_out),
    .io_enable(regs_58_io_enable)
  );
  FringeFF regs_59 ( // @[RegFile.scala 66:20:@42547.4]
    .clock(regs_59_clock),
    .reset(regs_59_reset),
    .io_in(regs_59_io_in),
    .io_reset(regs_59_io_reset),
    .io_out(regs_59_io_out),
    .io_enable(regs_59_io_enable)
  );
  FringeFF regs_60 ( // @[RegFile.scala 66:20:@42561.4]
    .clock(regs_60_clock),
    .reset(regs_60_reset),
    .io_in(regs_60_io_in),
    .io_reset(regs_60_io_reset),
    .io_out(regs_60_io_out),
    .io_enable(regs_60_io_enable)
  );
  FringeFF regs_61 ( // @[RegFile.scala 66:20:@42575.4]
    .clock(regs_61_clock),
    .reset(regs_61_reset),
    .io_in(regs_61_io_in),
    .io_reset(regs_61_io_reset),
    .io_out(regs_61_io_out),
    .io_enable(regs_61_io_enable)
  );
  FringeFF regs_62 ( // @[RegFile.scala 66:20:@42589.4]
    .clock(regs_62_clock),
    .reset(regs_62_reset),
    .io_in(regs_62_io_in),
    .io_reset(regs_62_io_reset),
    .io_out(regs_62_io_out),
    .io_enable(regs_62_io_enable)
  );
  FringeFF regs_63 ( // @[RegFile.scala 66:20:@42603.4]
    .clock(regs_63_clock),
    .reset(regs_63_reset),
    .io_in(regs_63_io_in),
    .io_reset(regs_63_io_reset),
    .io_out(regs_63_io_out),
    .io_enable(regs_63_io_enable)
  );
  FringeFF regs_64 ( // @[RegFile.scala 66:20:@42617.4]
    .clock(regs_64_clock),
    .reset(regs_64_reset),
    .io_in(regs_64_io_in),
    .io_reset(regs_64_io_reset),
    .io_out(regs_64_io_out),
    .io_enable(regs_64_io_enable)
  );
  FringeFF regs_65 ( // @[RegFile.scala 66:20:@42631.4]
    .clock(regs_65_clock),
    .reset(regs_65_reset),
    .io_in(regs_65_io_in),
    .io_reset(regs_65_io_reset),
    .io_out(regs_65_io_out),
    .io_enable(regs_65_io_enable)
  );
  FringeFF regs_66 ( // @[RegFile.scala 66:20:@42645.4]
    .clock(regs_66_clock),
    .reset(regs_66_reset),
    .io_in(regs_66_io_in),
    .io_reset(regs_66_io_reset),
    .io_out(regs_66_io_out),
    .io_enable(regs_66_io_enable)
  );
  FringeFF regs_67 ( // @[RegFile.scala 66:20:@42659.4]
    .clock(regs_67_clock),
    .reset(regs_67_reset),
    .io_in(regs_67_io_in),
    .io_reset(regs_67_io_reset),
    .io_out(regs_67_io_out),
    .io_enable(regs_67_io_enable)
  );
  FringeFF regs_68 ( // @[RegFile.scala 66:20:@42673.4]
    .clock(regs_68_clock),
    .reset(regs_68_reset),
    .io_in(regs_68_io_in),
    .io_reset(regs_68_io_reset),
    .io_out(regs_68_io_out),
    .io_enable(regs_68_io_enable)
  );
  FringeFF regs_69 ( // @[RegFile.scala 66:20:@42687.4]
    .clock(regs_69_clock),
    .reset(regs_69_reset),
    .io_in(regs_69_io_in),
    .io_reset(regs_69_io_reset),
    .io_out(regs_69_io_out),
    .io_enable(regs_69_io_enable)
  );
  FringeFF regs_70 ( // @[RegFile.scala 66:20:@42701.4]
    .clock(regs_70_clock),
    .reset(regs_70_reset),
    .io_in(regs_70_io_in),
    .io_reset(regs_70_io_reset),
    .io_out(regs_70_io_out),
    .io_enable(regs_70_io_enable)
  );
  FringeFF regs_71 ( // @[RegFile.scala 66:20:@42715.4]
    .clock(regs_71_clock),
    .reset(regs_71_reset),
    .io_in(regs_71_io_in),
    .io_reset(regs_71_io_reset),
    .io_out(regs_71_io_out),
    .io_enable(regs_71_io_enable)
  );
  FringeFF regs_72 ( // @[RegFile.scala 66:20:@42729.4]
    .clock(regs_72_clock),
    .reset(regs_72_reset),
    .io_in(regs_72_io_in),
    .io_reset(regs_72_io_reset),
    .io_out(regs_72_io_out),
    .io_enable(regs_72_io_enable)
  );
  FringeFF regs_73 ( // @[RegFile.scala 66:20:@42743.4]
    .clock(regs_73_clock),
    .reset(regs_73_reset),
    .io_in(regs_73_io_in),
    .io_reset(regs_73_io_reset),
    .io_out(regs_73_io_out),
    .io_enable(regs_73_io_enable)
  );
  FringeFF regs_74 ( // @[RegFile.scala 66:20:@42757.4]
    .clock(regs_74_clock),
    .reset(regs_74_reset),
    .io_in(regs_74_io_in),
    .io_reset(regs_74_io_reset),
    .io_out(regs_74_io_out),
    .io_enable(regs_74_io_enable)
  );
  FringeFF regs_75 ( // @[RegFile.scala 66:20:@42771.4]
    .clock(regs_75_clock),
    .reset(regs_75_reset),
    .io_in(regs_75_io_in),
    .io_reset(regs_75_io_reset),
    .io_out(regs_75_io_out),
    .io_enable(regs_75_io_enable)
  );
  FringeFF regs_76 ( // @[RegFile.scala 66:20:@42785.4]
    .clock(regs_76_clock),
    .reset(regs_76_reset),
    .io_in(regs_76_io_in),
    .io_reset(regs_76_io_reset),
    .io_out(regs_76_io_out),
    .io_enable(regs_76_io_enable)
  );
  FringeFF regs_77 ( // @[RegFile.scala 66:20:@42799.4]
    .clock(regs_77_clock),
    .reset(regs_77_reset),
    .io_in(regs_77_io_in),
    .io_reset(regs_77_io_reset),
    .io_out(regs_77_io_out),
    .io_enable(regs_77_io_enable)
  );
  FringeFF regs_78 ( // @[RegFile.scala 66:20:@42813.4]
    .clock(regs_78_clock),
    .reset(regs_78_reset),
    .io_in(regs_78_io_in),
    .io_reset(regs_78_io_reset),
    .io_out(regs_78_io_out),
    .io_enable(regs_78_io_enable)
  );
  FringeFF regs_79 ( // @[RegFile.scala 66:20:@42827.4]
    .clock(regs_79_clock),
    .reset(regs_79_reset),
    .io_in(regs_79_io_in),
    .io_reset(regs_79_io_reset),
    .io_out(regs_79_io_out),
    .io_enable(regs_79_io_enable)
  );
  FringeFF regs_80 ( // @[RegFile.scala 66:20:@42841.4]
    .clock(regs_80_clock),
    .reset(regs_80_reset),
    .io_in(regs_80_io_in),
    .io_reset(regs_80_io_reset),
    .io_out(regs_80_io_out),
    .io_enable(regs_80_io_enable)
  );
  FringeFF regs_81 ( // @[RegFile.scala 66:20:@42855.4]
    .clock(regs_81_clock),
    .reset(regs_81_reset),
    .io_in(regs_81_io_in),
    .io_reset(regs_81_io_reset),
    .io_out(regs_81_io_out),
    .io_enable(regs_81_io_enable)
  );
  FringeFF regs_82 ( // @[RegFile.scala 66:20:@42869.4]
    .clock(regs_82_clock),
    .reset(regs_82_reset),
    .io_in(regs_82_io_in),
    .io_reset(regs_82_io_reset),
    .io_out(regs_82_io_out),
    .io_enable(regs_82_io_enable)
  );
  FringeFF regs_83 ( // @[RegFile.scala 66:20:@42883.4]
    .clock(regs_83_clock),
    .reset(regs_83_reset),
    .io_in(regs_83_io_in),
    .io_reset(regs_83_io_reset),
    .io_out(regs_83_io_out),
    .io_enable(regs_83_io_enable)
  );
  FringeFF regs_84 ( // @[RegFile.scala 66:20:@42897.4]
    .clock(regs_84_clock),
    .reset(regs_84_reset),
    .io_in(regs_84_io_in),
    .io_reset(regs_84_io_reset),
    .io_out(regs_84_io_out),
    .io_enable(regs_84_io_enable)
  );
  FringeFF regs_85 ( // @[RegFile.scala 66:20:@42911.4]
    .clock(regs_85_clock),
    .reset(regs_85_reset),
    .io_in(regs_85_io_in),
    .io_reset(regs_85_io_reset),
    .io_out(regs_85_io_out),
    .io_enable(regs_85_io_enable)
  );
  FringeFF regs_86 ( // @[RegFile.scala 66:20:@42925.4]
    .clock(regs_86_clock),
    .reset(regs_86_reset),
    .io_in(regs_86_io_in),
    .io_reset(regs_86_io_reset),
    .io_out(regs_86_io_out),
    .io_enable(regs_86_io_enable)
  );
  FringeFF regs_87 ( // @[RegFile.scala 66:20:@42939.4]
    .clock(regs_87_clock),
    .reset(regs_87_reset),
    .io_in(regs_87_io_in),
    .io_reset(regs_87_io_reset),
    .io_out(regs_87_io_out),
    .io_enable(regs_87_io_enable)
  );
  FringeFF regs_88 ( // @[RegFile.scala 66:20:@42953.4]
    .clock(regs_88_clock),
    .reset(regs_88_reset),
    .io_in(regs_88_io_in),
    .io_reset(regs_88_io_reset),
    .io_out(regs_88_io_out),
    .io_enable(regs_88_io_enable)
  );
  FringeFF regs_89 ( // @[RegFile.scala 66:20:@42967.4]
    .clock(regs_89_clock),
    .reset(regs_89_reset),
    .io_in(regs_89_io_in),
    .io_reset(regs_89_io_reset),
    .io_out(regs_89_io_out),
    .io_enable(regs_89_io_enable)
  );
  FringeFF regs_90 ( // @[RegFile.scala 66:20:@42981.4]
    .clock(regs_90_clock),
    .reset(regs_90_reset),
    .io_in(regs_90_io_in),
    .io_reset(regs_90_io_reset),
    .io_out(regs_90_io_out),
    .io_enable(regs_90_io_enable)
  );
  FringeFF regs_91 ( // @[RegFile.scala 66:20:@42995.4]
    .clock(regs_91_clock),
    .reset(regs_91_reset),
    .io_in(regs_91_io_in),
    .io_reset(regs_91_io_reset),
    .io_out(regs_91_io_out),
    .io_enable(regs_91_io_enable)
  );
  FringeFF regs_92 ( // @[RegFile.scala 66:20:@43009.4]
    .clock(regs_92_clock),
    .reset(regs_92_reset),
    .io_in(regs_92_io_in),
    .io_reset(regs_92_io_reset),
    .io_out(regs_92_io_out),
    .io_enable(regs_92_io_enable)
  );
  FringeFF regs_93 ( // @[RegFile.scala 66:20:@43023.4]
    .clock(regs_93_clock),
    .reset(regs_93_reset),
    .io_in(regs_93_io_in),
    .io_reset(regs_93_io_reset),
    .io_out(regs_93_io_out),
    .io_enable(regs_93_io_enable)
  );
  FringeFF regs_94 ( // @[RegFile.scala 66:20:@43037.4]
    .clock(regs_94_clock),
    .reset(regs_94_reset),
    .io_in(regs_94_io_in),
    .io_reset(regs_94_io_reset),
    .io_out(regs_94_io_out),
    .io_enable(regs_94_io_enable)
  );
  FringeFF regs_95 ( // @[RegFile.scala 66:20:@43051.4]
    .clock(regs_95_clock),
    .reset(regs_95_reset),
    .io_in(regs_95_io_in),
    .io_reset(regs_95_io_reset),
    .io_out(regs_95_io_out),
    .io_enable(regs_95_io_enable)
  );
  FringeFF regs_96 ( // @[RegFile.scala 66:20:@43065.4]
    .clock(regs_96_clock),
    .reset(regs_96_reset),
    .io_in(regs_96_io_in),
    .io_reset(regs_96_io_reset),
    .io_out(regs_96_io_out),
    .io_enable(regs_96_io_enable)
  );
  FringeFF regs_97 ( // @[RegFile.scala 66:20:@43079.4]
    .clock(regs_97_clock),
    .reset(regs_97_reset),
    .io_in(regs_97_io_in),
    .io_reset(regs_97_io_reset),
    .io_out(regs_97_io_out),
    .io_enable(regs_97_io_enable)
  );
  FringeFF regs_98 ( // @[RegFile.scala 66:20:@43093.4]
    .clock(regs_98_clock),
    .reset(regs_98_reset),
    .io_in(regs_98_io_in),
    .io_reset(regs_98_io_reset),
    .io_out(regs_98_io_out),
    .io_enable(regs_98_io_enable)
  );
  FringeFF regs_99 ( // @[RegFile.scala 66:20:@43107.4]
    .clock(regs_99_clock),
    .reset(regs_99_reset),
    .io_in(regs_99_io_in),
    .io_reset(regs_99_io_reset),
    .io_out(regs_99_io_out),
    .io_enable(regs_99_io_enable)
  );
  FringeFF regs_100 ( // @[RegFile.scala 66:20:@43121.4]
    .clock(regs_100_clock),
    .reset(regs_100_reset),
    .io_in(regs_100_io_in),
    .io_reset(regs_100_io_reset),
    .io_out(regs_100_io_out),
    .io_enable(regs_100_io_enable)
  );
  FringeFF regs_101 ( // @[RegFile.scala 66:20:@43135.4]
    .clock(regs_101_clock),
    .reset(regs_101_reset),
    .io_in(regs_101_io_in),
    .io_reset(regs_101_io_reset),
    .io_out(regs_101_io_out),
    .io_enable(regs_101_io_enable)
  );
  FringeFF regs_102 ( // @[RegFile.scala 66:20:@43149.4]
    .clock(regs_102_clock),
    .reset(regs_102_reset),
    .io_in(regs_102_io_in),
    .io_reset(regs_102_io_reset),
    .io_out(regs_102_io_out),
    .io_enable(regs_102_io_enable)
  );
  FringeFF regs_103 ( // @[RegFile.scala 66:20:@43163.4]
    .clock(regs_103_clock),
    .reset(regs_103_reset),
    .io_in(regs_103_io_in),
    .io_reset(regs_103_io_reset),
    .io_out(regs_103_io_out),
    .io_enable(regs_103_io_enable)
  );
  FringeFF regs_104 ( // @[RegFile.scala 66:20:@43177.4]
    .clock(regs_104_clock),
    .reset(regs_104_reset),
    .io_in(regs_104_io_in),
    .io_reset(regs_104_io_reset),
    .io_out(regs_104_io_out),
    .io_enable(regs_104_io_enable)
  );
  FringeFF regs_105 ( // @[RegFile.scala 66:20:@43191.4]
    .clock(regs_105_clock),
    .reset(regs_105_reset),
    .io_in(regs_105_io_in),
    .io_reset(regs_105_io_reset),
    .io_out(regs_105_io_out),
    .io_enable(regs_105_io_enable)
  );
  FringeFF regs_106 ( // @[RegFile.scala 66:20:@43205.4]
    .clock(regs_106_clock),
    .reset(regs_106_reset),
    .io_in(regs_106_io_in),
    .io_reset(regs_106_io_reset),
    .io_out(regs_106_io_out),
    .io_enable(regs_106_io_enable)
  );
  FringeFF regs_107 ( // @[RegFile.scala 66:20:@43219.4]
    .clock(regs_107_clock),
    .reset(regs_107_reset),
    .io_in(regs_107_io_in),
    .io_reset(regs_107_io_reset),
    .io_out(regs_107_io_out),
    .io_enable(regs_107_io_enable)
  );
  FringeFF regs_108 ( // @[RegFile.scala 66:20:@43233.4]
    .clock(regs_108_clock),
    .reset(regs_108_reset),
    .io_in(regs_108_io_in),
    .io_reset(regs_108_io_reset),
    .io_out(regs_108_io_out),
    .io_enable(regs_108_io_enable)
  );
  FringeFF regs_109 ( // @[RegFile.scala 66:20:@43247.4]
    .clock(regs_109_clock),
    .reset(regs_109_reset),
    .io_in(regs_109_io_in),
    .io_reset(regs_109_io_reset),
    .io_out(regs_109_io_out),
    .io_enable(regs_109_io_enable)
  );
  FringeFF regs_110 ( // @[RegFile.scala 66:20:@43261.4]
    .clock(regs_110_clock),
    .reset(regs_110_reset),
    .io_in(regs_110_io_in),
    .io_reset(regs_110_io_reset),
    .io_out(regs_110_io_out),
    .io_enable(regs_110_io_enable)
  );
  FringeFF regs_111 ( // @[RegFile.scala 66:20:@43275.4]
    .clock(regs_111_clock),
    .reset(regs_111_reset),
    .io_in(regs_111_io_in),
    .io_reset(regs_111_io_reset),
    .io_out(regs_111_io_out),
    .io_enable(regs_111_io_enable)
  );
  FringeFF regs_112 ( // @[RegFile.scala 66:20:@43289.4]
    .clock(regs_112_clock),
    .reset(regs_112_reset),
    .io_in(regs_112_io_in),
    .io_reset(regs_112_io_reset),
    .io_out(regs_112_io_out),
    .io_enable(regs_112_io_enable)
  );
  FringeFF regs_113 ( // @[RegFile.scala 66:20:@43303.4]
    .clock(regs_113_clock),
    .reset(regs_113_reset),
    .io_in(regs_113_io_in),
    .io_reset(regs_113_io_reset),
    .io_out(regs_113_io_out),
    .io_enable(regs_113_io_enable)
  );
  FringeFF regs_114 ( // @[RegFile.scala 66:20:@43317.4]
    .clock(regs_114_clock),
    .reset(regs_114_reset),
    .io_in(regs_114_io_in),
    .io_reset(regs_114_io_reset),
    .io_out(regs_114_io_out),
    .io_enable(regs_114_io_enable)
  );
  FringeFF regs_115 ( // @[RegFile.scala 66:20:@43331.4]
    .clock(regs_115_clock),
    .reset(regs_115_reset),
    .io_in(regs_115_io_in),
    .io_reset(regs_115_io_reset),
    .io_out(regs_115_io_out),
    .io_enable(regs_115_io_enable)
  );
  FringeFF regs_116 ( // @[RegFile.scala 66:20:@43345.4]
    .clock(regs_116_clock),
    .reset(regs_116_reset),
    .io_in(regs_116_io_in),
    .io_reset(regs_116_io_reset),
    .io_out(regs_116_io_out),
    .io_enable(regs_116_io_enable)
  );
  FringeFF regs_117 ( // @[RegFile.scala 66:20:@43359.4]
    .clock(regs_117_clock),
    .reset(regs_117_reset),
    .io_in(regs_117_io_in),
    .io_reset(regs_117_io_reset),
    .io_out(regs_117_io_out),
    .io_enable(regs_117_io_enable)
  );
  FringeFF regs_118 ( // @[RegFile.scala 66:20:@43373.4]
    .clock(regs_118_clock),
    .reset(regs_118_reset),
    .io_in(regs_118_io_in),
    .io_reset(regs_118_io_reset),
    .io_out(regs_118_io_out),
    .io_enable(regs_118_io_enable)
  );
  FringeFF regs_119 ( // @[RegFile.scala 66:20:@43387.4]
    .clock(regs_119_clock),
    .reset(regs_119_reset),
    .io_in(regs_119_io_in),
    .io_reset(regs_119_io_reset),
    .io_out(regs_119_io_out),
    .io_enable(regs_119_io_enable)
  );
  FringeFF regs_120 ( // @[RegFile.scala 66:20:@43401.4]
    .clock(regs_120_clock),
    .reset(regs_120_reset),
    .io_in(regs_120_io_in),
    .io_reset(regs_120_io_reset),
    .io_out(regs_120_io_out),
    .io_enable(regs_120_io_enable)
  );
  FringeFF regs_121 ( // @[RegFile.scala 66:20:@43415.4]
    .clock(regs_121_clock),
    .reset(regs_121_reset),
    .io_in(regs_121_io_in),
    .io_reset(regs_121_io_reset),
    .io_out(regs_121_io_out),
    .io_enable(regs_121_io_enable)
  );
  FringeFF regs_122 ( // @[RegFile.scala 66:20:@43429.4]
    .clock(regs_122_clock),
    .reset(regs_122_reset),
    .io_in(regs_122_io_in),
    .io_reset(regs_122_io_reset),
    .io_out(regs_122_io_out),
    .io_enable(regs_122_io_enable)
  );
  FringeFF regs_123 ( // @[RegFile.scala 66:20:@43443.4]
    .clock(regs_123_clock),
    .reset(regs_123_reset),
    .io_in(regs_123_io_in),
    .io_reset(regs_123_io_reset),
    .io_out(regs_123_io_out),
    .io_enable(regs_123_io_enable)
  );
  FringeFF regs_124 ( // @[RegFile.scala 66:20:@43457.4]
    .clock(regs_124_clock),
    .reset(regs_124_reset),
    .io_in(regs_124_io_in),
    .io_reset(regs_124_io_reset),
    .io_out(regs_124_io_out),
    .io_enable(regs_124_io_enable)
  );
  FringeFF regs_125 ( // @[RegFile.scala 66:20:@43471.4]
    .clock(regs_125_clock),
    .reset(regs_125_reset),
    .io_in(regs_125_io_in),
    .io_reset(regs_125_io_reset),
    .io_out(regs_125_io_out),
    .io_enable(regs_125_io_enable)
  );
  FringeFF regs_126 ( // @[RegFile.scala 66:20:@43485.4]
    .clock(regs_126_clock),
    .reset(regs_126_reset),
    .io_in(regs_126_io_in),
    .io_reset(regs_126_io_reset),
    .io_out(regs_126_io_out),
    .io_enable(regs_126_io_enable)
  );
  FringeFF regs_127 ( // @[RegFile.scala 66:20:@43499.4]
    .clock(regs_127_clock),
    .reset(regs_127_reset),
    .io_in(regs_127_io_in),
    .io_reset(regs_127_io_reset),
    .io_out(regs_127_io_out),
    .io_enable(regs_127_io_enable)
  );
  FringeFF regs_128 ( // @[RegFile.scala 66:20:@43513.4]
    .clock(regs_128_clock),
    .reset(regs_128_reset),
    .io_in(regs_128_io_in),
    .io_reset(regs_128_io_reset),
    .io_out(regs_128_io_out),
    .io_enable(regs_128_io_enable)
  );
  FringeFF regs_129 ( // @[RegFile.scala 66:20:@43527.4]
    .clock(regs_129_clock),
    .reset(regs_129_reset),
    .io_in(regs_129_io_in),
    .io_reset(regs_129_io_reset),
    .io_out(regs_129_io_out),
    .io_enable(regs_129_io_enable)
  );
  FringeFF regs_130 ( // @[RegFile.scala 66:20:@43541.4]
    .clock(regs_130_clock),
    .reset(regs_130_reset),
    .io_in(regs_130_io_in),
    .io_reset(regs_130_io_reset),
    .io_out(regs_130_io_out),
    .io_enable(regs_130_io_enable)
  );
  FringeFF regs_131 ( // @[RegFile.scala 66:20:@43555.4]
    .clock(regs_131_clock),
    .reset(regs_131_reset),
    .io_in(regs_131_io_in),
    .io_reset(regs_131_io_reset),
    .io_out(regs_131_io_out),
    .io_enable(regs_131_io_enable)
  );
  FringeFF regs_132 ( // @[RegFile.scala 66:20:@43569.4]
    .clock(regs_132_clock),
    .reset(regs_132_reset),
    .io_in(regs_132_io_in),
    .io_reset(regs_132_io_reset),
    .io_out(regs_132_io_out),
    .io_enable(regs_132_io_enable)
  );
  FringeFF regs_133 ( // @[RegFile.scala 66:20:@43583.4]
    .clock(regs_133_clock),
    .reset(regs_133_reset),
    .io_in(regs_133_io_in),
    .io_reset(regs_133_io_reset),
    .io_out(regs_133_io_out),
    .io_enable(regs_133_io_enable)
  );
  FringeFF regs_134 ( // @[RegFile.scala 66:20:@43597.4]
    .clock(regs_134_clock),
    .reset(regs_134_reset),
    .io_in(regs_134_io_in),
    .io_reset(regs_134_io_reset),
    .io_out(regs_134_io_out),
    .io_enable(regs_134_io_enable)
  );
  FringeFF regs_135 ( // @[RegFile.scala 66:20:@43611.4]
    .clock(regs_135_clock),
    .reset(regs_135_reset),
    .io_in(regs_135_io_in),
    .io_reset(regs_135_io_reset),
    .io_out(regs_135_io_out),
    .io_enable(regs_135_io_enable)
  );
  FringeFF regs_136 ( // @[RegFile.scala 66:20:@43625.4]
    .clock(regs_136_clock),
    .reset(regs_136_reset),
    .io_in(regs_136_io_in),
    .io_reset(regs_136_io_reset),
    .io_out(regs_136_io_out),
    .io_enable(regs_136_io_enable)
  );
  FringeFF regs_137 ( // @[RegFile.scala 66:20:@43639.4]
    .clock(regs_137_clock),
    .reset(regs_137_reset),
    .io_in(regs_137_io_in),
    .io_reset(regs_137_io_reset),
    .io_out(regs_137_io_out),
    .io_enable(regs_137_io_enable)
  );
  FringeFF regs_138 ( // @[RegFile.scala 66:20:@43653.4]
    .clock(regs_138_clock),
    .reset(regs_138_reset),
    .io_in(regs_138_io_in),
    .io_reset(regs_138_io_reset),
    .io_out(regs_138_io_out),
    .io_enable(regs_138_io_enable)
  );
  FringeFF regs_139 ( // @[RegFile.scala 66:20:@43667.4]
    .clock(regs_139_clock),
    .reset(regs_139_reset),
    .io_in(regs_139_io_in),
    .io_reset(regs_139_io_reset),
    .io_out(regs_139_io_out),
    .io_enable(regs_139_io_enable)
  );
  FringeFF regs_140 ( // @[RegFile.scala 66:20:@43681.4]
    .clock(regs_140_clock),
    .reset(regs_140_reset),
    .io_in(regs_140_io_in),
    .io_reset(regs_140_io_reset),
    .io_out(regs_140_io_out),
    .io_enable(regs_140_io_enable)
  );
  FringeFF regs_141 ( // @[RegFile.scala 66:20:@43695.4]
    .clock(regs_141_clock),
    .reset(regs_141_reset),
    .io_in(regs_141_io_in),
    .io_reset(regs_141_io_reset),
    .io_out(regs_141_io_out),
    .io_enable(regs_141_io_enable)
  );
  FringeFF regs_142 ( // @[RegFile.scala 66:20:@43709.4]
    .clock(regs_142_clock),
    .reset(regs_142_reset),
    .io_in(regs_142_io_in),
    .io_reset(regs_142_io_reset),
    .io_out(regs_142_io_out),
    .io_enable(regs_142_io_enable)
  );
  FringeFF regs_143 ( // @[RegFile.scala 66:20:@43723.4]
    .clock(regs_143_clock),
    .reset(regs_143_reset),
    .io_in(regs_143_io_in),
    .io_reset(regs_143_io_reset),
    .io_out(regs_143_io_out),
    .io_enable(regs_143_io_enable)
  );
  FringeFF regs_144 ( // @[RegFile.scala 66:20:@43737.4]
    .clock(regs_144_clock),
    .reset(regs_144_reset),
    .io_in(regs_144_io_in),
    .io_reset(regs_144_io_reset),
    .io_out(regs_144_io_out),
    .io_enable(regs_144_io_enable)
  );
  FringeFF regs_145 ( // @[RegFile.scala 66:20:@43751.4]
    .clock(regs_145_clock),
    .reset(regs_145_reset),
    .io_in(regs_145_io_in),
    .io_reset(regs_145_io_reset),
    .io_out(regs_145_io_out),
    .io_enable(regs_145_io_enable)
  );
  FringeFF regs_146 ( // @[RegFile.scala 66:20:@43765.4]
    .clock(regs_146_clock),
    .reset(regs_146_reset),
    .io_in(regs_146_io_in),
    .io_reset(regs_146_io_reset),
    .io_out(regs_146_io_out),
    .io_enable(regs_146_io_enable)
  );
  FringeFF regs_147 ( // @[RegFile.scala 66:20:@43779.4]
    .clock(regs_147_clock),
    .reset(regs_147_reset),
    .io_in(regs_147_io_in),
    .io_reset(regs_147_io_reset),
    .io_out(regs_147_io_out),
    .io_enable(regs_147_io_enable)
  );
  FringeFF regs_148 ( // @[RegFile.scala 66:20:@43793.4]
    .clock(regs_148_clock),
    .reset(regs_148_reset),
    .io_in(regs_148_io_in),
    .io_reset(regs_148_io_reset),
    .io_out(regs_148_io_out),
    .io_enable(regs_148_io_enable)
  );
  FringeFF regs_149 ( // @[RegFile.scala 66:20:@43807.4]
    .clock(regs_149_clock),
    .reset(regs_149_reset),
    .io_in(regs_149_io_in),
    .io_reset(regs_149_io_reset),
    .io_out(regs_149_io_out),
    .io_enable(regs_149_io_enable)
  );
  FringeFF regs_150 ( // @[RegFile.scala 66:20:@43821.4]
    .clock(regs_150_clock),
    .reset(regs_150_reset),
    .io_in(regs_150_io_in),
    .io_reset(regs_150_io_reset),
    .io_out(regs_150_io_out),
    .io_enable(regs_150_io_enable)
  );
  FringeFF regs_151 ( // @[RegFile.scala 66:20:@43835.4]
    .clock(regs_151_clock),
    .reset(regs_151_reset),
    .io_in(regs_151_io_in),
    .io_reset(regs_151_io_reset),
    .io_out(regs_151_io_out),
    .io_enable(regs_151_io_enable)
  );
  FringeFF regs_152 ( // @[RegFile.scala 66:20:@43849.4]
    .clock(regs_152_clock),
    .reset(regs_152_reset),
    .io_in(regs_152_io_in),
    .io_reset(regs_152_io_reset),
    .io_out(regs_152_io_out),
    .io_enable(regs_152_io_enable)
  );
  FringeFF regs_153 ( // @[RegFile.scala 66:20:@43863.4]
    .clock(regs_153_clock),
    .reset(regs_153_reset),
    .io_in(regs_153_io_in),
    .io_reset(regs_153_io_reset),
    .io_out(regs_153_io_out),
    .io_enable(regs_153_io_enable)
  );
  FringeFF regs_154 ( // @[RegFile.scala 66:20:@43877.4]
    .clock(regs_154_clock),
    .reset(regs_154_reset),
    .io_in(regs_154_io_in),
    .io_reset(regs_154_io_reset),
    .io_out(regs_154_io_out),
    .io_enable(regs_154_io_enable)
  );
  FringeFF regs_155 ( // @[RegFile.scala 66:20:@43891.4]
    .clock(regs_155_clock),
    .reset(regs_155_reset),
    .io_in(regs_155_io_in),
    .io_reset(regs_155_io_reset),
    .io_out(regs_155_io_out),
    .io_enable(regs_155_io_enable)
  );
  FringeFF regs_156 ( // @[RegFile.scala 66:20:@43905.4]
    .clock(regs_156_clock),
    .reset(regs_156_reset),
    .io_in(regs_156_io_in),
    .io_reset(regs_156_io_reset),
    .io_out(regs_156_io_out),
    .io_enable(regs_156_io_enable)
  );
  FringeFF regs_157 ( // @[RegFile.scala 66:20:@43919.4]
    .clock(regs_157_clock),
    .reset(regs_157_reset),
    .io_in(regs_157_io_in),
    .io_reset(regs_157_io_reset),
    .io_out(regs_157_io_out),
    .io_enable(regs_157_io_enable)
  );
  FringeFF regs_158 ( // @[RegFile.scala 66:20:@43933.4]
    .clock(regs_158_clock),
    .reset(regs_158_reset),
    .io_in(regs_158_io_in),
    .io_reset(regs_158_io_reset),
    .io_out(regs_158_io_out),
    .io_enable(regs_158_io_enable)
  );
  FringeFF regs_159 ( // @[RegFile.scala 66:20:@43947.4]
    .clock(regs_159_clock),
    .reset(regs_159_reset),
    .io_in(regs_159_io_in),
    .io_reset(regs_159_io_reset),
    .io_out(regs_159_io_out),
    .io_enable(regs_159_io_enable)
  );
  FringeFF regs_160 ( // @[RegFile.scala 66:20:@43961.4]
    .clock(regs_160_clock),
    .reset(regs_160_reset),
    .io_in(regs_160_io_in),
    .io_reset(regs_160_io_reset),
    .io_out(regs_160_io_out),
    .io_enable(regs_160_io_enable)
  );
  FringeFF regs_161 ( // @[RegFile.scala 66:20:@43975.4]
    .clock(regs_161_clock),
    .reset(regs_161_reset),
    .io_in(regs_161_io_in),
    .io_reset(regs_161_io_reset),
    .io_out(regs_161_io_out),
    .io_enable(regs_161_io_enable)
  );
  FringeFF regs_162 ( // @[RegFile.scala 66:20:@43989.4]
    .clock(regs_162_clock),
    .reset(regs_162_reset),
    .io_in(regs_162_io_in),
    .io_reset(regs_162_io_reset),
    .io_out(regs_162_io_out),
    .io_enable(regs_162_io_enable)
  );
  FringeFF regs_163 ( // @[RegFile.scala 66:20:@44003.4]
    .clock(regs_163_clock),
    .reset(regs_163_reset),
    .io_in(regs_163_io_in),
    .io_reset(regs_163_io_reset),
    .io_out(regs_163_io_out),
    .io_enable(regs_163_io_enable)
  );
  FringeFF regs_164 ( // @[RegFile.scala 66:20:@44017.4]
    .clock(regs_164_clock),
    .reset(regs_164_reset),
    .io_in(regs_164_io_in),
    .io_reset(regs_164_io_reset),
    .io_out(regs_164_io_out),
    .io_enable(regs_164_io_enable)
  );
  FringeFF regs_165 ( // @[RegFile.scala 66:20:@44031.4]
    .clock(regs_165_clock),
    .reset(regs_165_reset),
    .io_in(regs_165_io_in),
    .io_reset(regs_165_io_reset),
    .io_out(regs_165_io_out),
    .io_enable(regs_165_io_enable)
  );
  FringeFF regs_166 ( // @[RegFile.scala 66:20:@44045.4]
    .clock(regs_166_clock),
    .reset(regs_166_reset),
    .io_in(regs_166_io_in),
    .io_reset(regs_166_io_reset),
    .io_out(regs_166_io_out),
    .io_enable(regs_166_io_enable)
  );
  FringeFF regs_167 ( // @[RegFile.scala 66:20:@44059.4]
    .clock(regs_167_clock),
    .reset(regs_167_reset),
    .io_in(regs_167_io_in),
    .io_reset(regs_167_io_reset),
    .io_out(regs_167_io_out),
    .io_enable(regs_167_io_enable)
  );
  FringeFF regs_168 ( // @[RegFile.scala 66:20:@44073.4]
    .clock(regs_168_clock),
    .reset(regs_168_reset),
    .io_in(regs_168_io_in),
    .io_reset(regs_168_io_reset),
    .io_out(regs_168_io_out),
    .io_enable(regs_168_io_enable)
  );
  FringeFF regs_169 ( // @[RegFile.scala 66:20:@44087.4]
    .clock(regs_169_clock),
    .reset(regs_169_reset),
    .io_in(regs_169_io_in),
    .io_reset(regs_169_io_reset),
    .io_out(regs_169_io_out),
    .io_enable(regs_169_io_enable)
  );
  FringeFF regs_170 ( // @[RegFile.scala 66:20:@44101.4]
    .clock(regs_170_clock),
    .reset(regs_170_reset),
    .io_in(regs_170_io_in),
    .io_reset(regs_170_io_reset),
    .io_out(regs_170_io_out),
    .io_enable(regs_170_io_enable)
  );
  FringeFF regs_171 ( // @[RegFile.scala 66:20:@44115.4]
    .clock(regs_171_clock),
    .reset(regs_171_reset),
    .io_in(regs_171_io_in),
    .io_reset(regs_171_io_reset),
    .io_out(regs_171_io_out),
    .io_enable(regs_171_io_enable)
  );
  FringeFF regs_172 ( // @[RegFile.scala 66:20:@44129.4]
    .clock(regs_172_clock),
    .reset(regs_172_reset),
    .io_in(regs_172_io_in),
    .io_reset(regs_172_io_reset),
    .io_out(regs_172_io_out),
    .io_enable(regs_172_io_enable)
  );
  FringeFF regs_173 ( // @[RegFile.scala 66:20:@44143.4]
    .clock(regs_173_clock),
    .reset(regs_173_reset),
    .io_in(regs_173_io_in),
    .io_reset(regs_173_io_reset),
    .io_out(regs_173_io_out),
    .io_enable(regs_173_io_enable)
  );
  FringeFF regs_174 ( // @[RegFile.scala 66:20:@44157.4]
    .clock(regs_174_clock),
    .reset(regs_174_reset),
    .io_in(regs_174_io_in),
    .io_reset(regs_174_io_reset),
    .io_out(regs_174_io_out),
    .io_enable(regs_174_io_enable)
  );
  FringeFF regs_175 ( // @[RegFile.scala 66:20:@44171.4]
    .clock(regs_175_clock),
    .reset(regs_175_reset),
    .io_in(regs_175_io_in),
    .io_reset(regs_175_io_reset),
    .io_out(regs_175_io_out),
    .io_enable(regs_175_io_enable)
  );
  FringeFF regs_176 ( // @[RegFile.scala 66:20:@44185.4]
    .clock(regs_176_clock),
    .reset(regs_176_reset),
    .io_in(regs_176_io_in),
    .io_reset(regs_176_io_reset),
    .io_out(regs_176_io_out),
    .io_enable(regs_176_io_enable)
  );
  FringeFF regs_177 ( // @[RegFile.scala 66:20:@44199.4]
    .clock(regs_177_clock),
    .reset(regs_177_reset),
    .io_in(regs_177_io_in),
    .io_reset(regs_177_io_reset),
    .io_out(regs_177_io_out),
    .io_enable(regs_177_io_enable)
  );
  FringeFF regs_178 ( // @[RegFile.scala 66:20:@44213.4]
    .clock(regs_178_clock),
    .reset(regs_178_reset),
    .io_in(regs_178_io_in),
    .io_reset(regs_178_io_reset),
    .io_out(regs_178_io_out),
    .io_enable(regs_178_io_enable)
  );
  FringeFF regs_179 ( // @[RegFile.scala 66:20:@44227.4]
    .clock(regs_179_clock),
    .reset(regs_179_reset),
    .io_in(regs_179_io_in),
    .io_reset(regs_179_io_reset),
    .io_out(regs_179_io_out),
    .io_enable(regs_179_io_enable)
  );
  FringeFF regs_180 ( // @[RegFile.scala 66:20:@44241.4]
    .clock(regs_180_clock),
    .reset(regs_180_reset),
    .io_in(regs_180_io_in),
    .io_reset(regs_180_io_reset),
    .io_out(regs_180_io_out),
    .io_enable(regs_180_io_enable)
  );
  FringeFF regs_181 ( // @[RegFile.scala 66:20:@44255.4]
    .clock(regs_181_clock),
    .reset(regs_181_reset),
    .io_in(regs_181_io_in),
    .io_reset(regs_181_io_reset),
    .io_out(regs_181_io_out),
    .io_enable(regs_181_io_enable)
  );
  FringeFF regs_182 ( // @[RegFile.scala 66:20:@44269.4]
    .clock(regs_182_clock),
    .reset(regs_182_reset),
    .io_in(regs_182_io_in),
    .io_reset(regs_182_io_reset),
    .io_out(regs_182_io_out),
    .io_enable(regs_182_io_enable)
  );
  FringeFF regs_183 ( // @[RegFile.scala 66:20:@44283.4]
    .clock(regs_183_clock),
    .reset(regs_183_reset),
    .io_in(regs_183_io_in),
    .io_reset(regs_183_io_reset),
    .io_out(regs_183_io_out),
    .io_enable(regs_183_io_enable)
  );
  FringeFF regs_184 ( // @[RegFile.scala 66:20:@44297.4]
    .clock(regs_184_clock),
    .reset(regs_184_reset),
    .io_in(regs_184_io_in),
    .io_reset(regs_184_io_reset),
    .io_out(regs_184_io_out),
    .io_enable(regs_184_io_enable)
  );
  FringeFF regs_185 ( // @[RegFile.scala 66:20:@44311.4]
    .clock(regs_185_clock),
    .reset(regs_185_reset),
    .io_in(regs_185_io_in),
    .io_reset(regs_185_io_reset),
    .io_out(regs_185_io_out),
    .io_enable(regs_185_io_enable)
  );
  FringeFF regs_186 ( // @[RegFile.scala 66:20:@44325.4]
    .clock(regs_186_clock),
    .reset(regs_186_reset),
    .io_in(regs_186_io_in),
    .io_reset(regs_186_io_reset),
    .io_out(regs_186_io_out),
    .io_enable(regs_186_io_enable)
  );
  FringeFF regs_187 ( // @[RegFile.scala 66:20:@44339.4]
    .clock(regs_187_clock),
    .reset(regs_187_reset),
    .io_in(regs_187_io_in),
    .io_reset(regs_187_io_reset),
    .io_out(regs_187_io_out),
    .io_enable(regs_187_io_enable)
  );
  FringeFF regs_188 ( // @[RegFile.scala 66:20:@44353.4]
    .clock(regs_188_clock),
    .reset(regs_188_reset),
    .io_in(regs_188_io_in),
    .io_reset(regs_188_io_reset),
    .io_out(regs_188_io_out),
    .io_enable(regs_188_io_enable)
  );
  FringeFF regs_189 ( // @[RegFile.scala 66:20:@44367.4]
    .clock(regs_189_clock),
    .reset(regs_189_reset),
    .io_in(regs_189_io_in),
    .io_reset(regs_189_io_reset),
    .io_out(regs_189_io_out),
    .io_enable(regs_189_io_enable)
  );
  FringeFF regs_190 ( // @[RegFile.scala 66:20:@44381.4]
    .clock(regs_190_clock),
    .reset(regs_190_reset),
    .io_in(regs_190_io_in),
    .io_reset(regs_190_io_reset),
    .io_out(regs_190_io_out),
    .io_enable(regs_190_io_enable)
  );
  FringeFF regs_191 ( // @[RegFile.scala 66:20:@44395.4]
    .clock(regs_191_clock),
    .reset(regs_191_reset),
    .io_in(regs_191_io_in),
    .io_reset(regs_191_io_reset),
    .io_out(regs_191_io_out),
    .io_enable(regs_191_io_enable)
  );
  FringeFF regs_192 ( // @[RegFile.scala 66:20:@44409.4]
    .clock(regs_192_clock),
    .reset(regs_192_reset),
    .io_in(regs_192_io_in),
    .io_reset(regs_192_io_reset),
    .io_out(regs_192_io_out),
    .io_enable(regs_192_io_enable)
  );
  FringeFF regs_193 ( // @[RegFile.scala 66:20:@44423.4]
    .clock(regs_193_clock),
    .reset(regs_193_reset),
    .io_in(regs_193_io_in),
    .io_reset(regs_193_io_reset),
    .io_out(regs_193_io_out),
    .io_enable(regs_193_io_enable)
  );
  FringeFF regs_194 ( // @[RegFile.scala 66:20:@44437.4]
    .clock(regs_194_clock),
    .reset(regs_194_reset),
    .io_in(regs_194_io_in),
    .io_reset(regs_194_io_reset),
    .io_out(regs_194_io_out),
    .io_enable(regs_194_io_enable)
  );
  FringeFF regs_195 ( // @[RegFile.scala 66:20:@44451.4]
    .clock(regs_195_clock),
    .reset(regs_195_reset),
    .io_in(regs_195_io_in),
    .io_reset(regs_195_io_reset),
    .io_out(regs_195_io_out),
    .io_enable(regs_195_io_enable)
  );
  FringeFF regs_196 ( // @[RegFile.scala 66:20:@44465.4]
    .clock(regs_196_clock),
    .reset(regs_196_reset),
    .io_in(regs_196_io_in),
    .io_reset(regs_196_io_reset),
    .io_out(regs_196_io_out),
    .io_enable(regs_196_io_enable)
  );
  FringeFF regs_197 ( // @[RegFile.scala 66:20:@44479.4]
    .clock(regs_197_clock),
    .reset(regs_197_reset),
    .io_in(regs_197_io_in),
    .io_reset(regs_197_io_reset),
    .io_out(regs_197_io_out),
    .io_enable(regs_197_io_enable)
  );
  FringeFF regs_198 ( // @[RegFile.scala 66:20:@44493.4]
    .clock(regs_198_clock),
    .reset(regs_198_reset),
    .io_in(regs_198_io_in),
    .io_reset(regs_198_io_reset),
    .io_out(regs_198_io_out),
    .io_enable(regs_198_io_enable)
  );
  FringeFF regs_199 ( // @[RegFile.scala 66:20:@44507.4]
    .clock(regs_199_clock),
    .reset(regs_199_reset),
    .io_in(regs_199_io_in),
    .io_reset(regs_199_io_reset),
    .io_out(regs_199_io_out),
    .io_enable(regs_199_io_enable)
  );
  FringeFF regs_200 ( // @[RegFile.scala 66:20:@44521.4]
    .clock(regs_200_clock),
    .reset(regs_200_reset),
    .io_in(regs_200_io_in),
    .io_reset(regs_200_io_reset),
    .io_out(regs_200_io_out),
    .io_enable(regs_200_io_enable)
  );
  FringeFF regs_201 ( // @[RegFile.scala 66:20:@44535.4]
    .clock(regs_201_clock),
    .reset(regs_201_reset),
    .io_in(regs_201_io_in),
    .io_reset(regs_201_io_reset),
    .io_out(regs_201_io_out),
    .io_enable(regs_201_io_enable)
  );
  FringeFF regs_202 ( // @[RegFile.scala 66:20:@44549.4]
    .clock(regs_202_clock),
    .reset(regs_202_reset),
    .io_in(regs_202_io_in),
    .io_reset(regs_202_io_reset),
    .io_out(regs_202_io_out),
    .io_enable(regs_202_io_enable)
  );
  FringeFF regs_203 ( // @[RegFile.scala 66:20:@44563.4]
    .clock(regs_203_clock),
    .reset(regs_203_reset),
    .io_in(regs_203_io_in),
    .io_reset(regs_203_io_reset),
    .io_out(regs_203_io_out),
    .io_enable(regs_203_io_enable)
  );
  FringeFF regs_204 ( // @[RegFile.scala 66:20:@44577.4]
    .clock(regs_204_clock),
    .reset(regs_204_reset),
    .io_in(regs_204_io_in),
    .io_reset(regs_204_io_reset),
    .io_out(regs_204_io_out),
    .io_enable(regs_204_io_enable)
  );
  FringeFF regs_205 ( // @[RegFile.scala 66:20:@44591.4]
    .clock(regs_205_clock),
    .reset(regs_205_reset),
    .io_in(regs_205_io_in),
    .io_reset(regs_205_io_reset),
    .io_out(regs_205_io_out),
    .io_enable(regs_205_io_enable)
  );
  FringeFF regs_206 ( // @[RegFile.scala 66:20:@44605.4]
    .clock(regs_206_clock),
    .reset(regs_206_reset),
    .io_in(regs_206_io_in),
    .io_reset(regs_206_io_reset),
    .io_out(regs_206_io_out),
    .io_enable(regs_206_io_enable)
  );
  FringeFF regs_207 ( // @[RegFile.scala 66:20:@44619.4]
    .clock(regs_207_clock),
    .reset(regs_207_reset),
    .io_in(regs_207_io_in),
    .io_reset(regs_207_io_reset),
    .io_out(regs_207_io_out),
    .io_enable(regs_207_io_enable)
  );
  FringeFF regs_208 ( // @[RegFile.scala 66:20:@44633.4]
    .clock(regs_208_clock),
    .reset(regs_208_reset),
    .io_in(regs_208_io_in),
    .io_reset(regs_208_io_reset),
    .io_out(regs_208_io_out),
    .io_enable(regs_208_io_enable)
  );
  FringeFF regs_209 ( // @[RegFile.scala 66:20:@44647.4]
    .clock(regs_209_clock),
    .reset(regs_209_reset),
    .io_in(regs_209_io_in),
    .io_reset(regs_209_io_reset),
    .io_out(regs_209_io_out),
    .io_enable(regs_209_io_enable)
  );
  FringeFF regs_210 ( // @[RegFile.scala 66:20:@44661.4]
    .clock(regs_210_clock),
    .reset(regs_210_reset),
    .io_in(regs_210_io_in),
    .io_reset(regs_210_io_reset),
    .io_out(regs_210_io_out),
    .io_enable(regs_210_io_enable)
  );
  FringeFF regs_211 ( // @[RegFile.scala 66:20:@44675.4]
    .clock(regs_211_clock),
    .reset(regs_211_reset),
    .io_in(regs_211_io_in),
    .io_reset(regs_211_io_reset),
    .io_out(regs_211_io_out),
    .io_enable(regs_211_io_enable)
  );
  FringeFF regs_212 ( // @[RegFile.scala 66:20:@44689.4]
    .clock(regs_212_clock),
    .reset(regs_212_reset),
    .io_in(regs_212_io_in),
    .io_reset(regs_212_io_reset),
    .io_out(regs_212_io_out),
    .io_enable(regs_212_io_enable)
  );
  FringeFF regs_213 ( // @[RegFile.scala 66:20:@44703.4]
    .clock(regs_213_clock),
    .reset(regs_213_reset),
    .io_in(regs_213_io_in),
    .io_reset(regs_213_io_reset),
    .io_out(regs_213_io_out),
    .io_enable(regs_213_io_enable)
  );
  FringeFF regs_214 ( // @[RegFile.scala 66:20:@44717.4]
    .clock(regs_214_clock),
    .reset(regs_214_reset),
    .io_in(regs_214_io_in),
    .io_reset(regs_214_io_reset),
    .io_out(regs_214_io_out),
    .io_enable(regs_214_io_enable)
  );
  FringeFF regs_215 ( // @[RegFile.scala 66:20:@44731.4]
    .clock(regs_215_clock),
    .reset(regs_215_reset),
    .io_in(regs_215_io_in),
    .io_reset(regs_215_io_reset),
    .io_out(regs_215_io_out),
    .io_enable(regs_215_io_enable)
  );
  FringeFF regs_216 ( // @[RegFile.scala 66:20:@44745.4]
    .clock(regs_216_clock),
    .reset(regs_216_reset),
    .io_in(regs_216_io_in),
    .io_reset(regs_216_io_reset),
    .io_out(regs_216_io_out),
    .io_enable(regs_216_io_enable)
  );
  FringeFF regs_217 ( // @[RegFile.scala 66:20:@44759.4]
    .clock(regs_217_clock),
    .reset(regs_217_reset),
    .io_in(regs_217_io_in),
    .io_reset(regs_217_io_reset),
    .io_out(regs_217_io_out),
    .io_enable(regs_217_io_enable)
  );
  FringeFF regs_218 ( // @[RegFile.scala 66:20:@44773.4]
    .clock(regs_218_clock),
    .reset(regs_218_reset),
    .io_in(regs_218_io_in),
    .io_reset(regs_218_io_reset),
    .io_out(regs_218_io_out),
    .io_enable(regs_218_io_enable)
  );
  FringeFF regs_219 ( // @[RegFile.scala 66:20:@44787.4]
    .clock(regs_219_clock),
    .reset(regs_219_reset),
    .io_in(regs_219_io_in),
    .io_reset(regs_219_io_reset),
    .io_out(regs_219_io_out),
    .io_enable(regs_219_io_enable)
  );
  FringeFF regs_220 ( // @[RegFile.scala 66:20:@44801.4]
    .clock(regs_220_clock),
    .reset(regs_220_reset),
    .io_in(regs_220_io_in),
    .io_reset(regs_220_io_reset),
    .io_out(regs_220_io_out),
    .io_enable(regs_220_io_enable)
  );
  FringeFF regs_221 ( // @[RegFile.scala 66:20:@44815.4]
    .clock(regs_221_clock),
    .reset(regs_221_reset),
    .io_in(regs_221_io_in),
    .io_reset(regs_221_io_reset),
    .io_out(regs_221_io_out),
    .io_enable(regs_221_io_enable)
  );
  FringeFF regs_222 ( // @[RegFile.scala 66:20:@44829.4]
    .clock(regs_222_clock),
    .reset(regs_222_reset),
    .io_in(regs_222_io_in),
    .io_reset(regs_222_io_reset),
    .io_out(regs_222_io_out),
    .io_enable(regs_222_io_enable)
  );
  FringeFF regs_223 ( // @[RegFile.scala 66:20:@44843.4]
    .clock(regs_223_clock),
    .reset(regs_223_reset),
    .io_in(regs_223_io_in),
    .io_reset(regs_223_io_reset),
    .io_out(regs_223_io_out),
    .io_enable(regs_223_io_enable)
  );
  FringeFF regs_224 ( // @[RegFile.scala 66:20:@44857.4]
    .clock(regs_224_clock),
    .reset(regs_224_reset),
    .io_in(regs_224_io_in),
    .io_reset(regs_224_io_reset),
    .io_out(regs_224_io_out),
    .io_enable(regs_224_io_enable)
  );
  FringeFF regs_225 ( // @[RegFile.scala 66:20:@44871.4]
    .clock(regs_225_clock),
    .reset(regs_225_reset),
    .io_in(regs_225_io_in),
    .io_reset(regs_225_io_reset),
    .io_out(regs_225_io_out),
    .io_enable(regs_225_io_enable)
  );
  FringeFF regs_226 ( // @[RegFile.scala 66:20:@44885.4]
    .clock(regs_226_clock),
    .reset(regs_226_reset),
    .io_in(regs_226_io_in),
    .io_reset(regs_226_io_reset),
    .io_out(regs_226_io_out),
    .io_enable(regs_226_io_enable)
  );
  FringeFF regs_227 ( // @[RegFile.scala 66:20:@44899.4]
    .clock(regs_227_clock),
    .reset(regs_227_reset),
    .io_in(regs_227_io_in),
    .io_reset(regs_227_io_reset),
    .io_out(regs_227_io_out),
    .io_enable(regs_227_io_enable)
  );
  FringeFF regs_228 ( // @[RegFile.scala 66:20:@44913.4]
    .clock(regs_228_clock),
    .reset(regs_228_reset),
    .io_in(regs_228_io_in),
    .io_reset(regs_228_io_reset),
    .io_out(regs_228_io_out),
    .io_enable(regs_228_io_enable)
  );
  FringeFF regs_229 ( // @[RegFile.scala 66:20:@44927.4]
    .clock(regs_229_clock),
    .reset(regs_229_reset),
    .io_in(regs_229_io_in),
    .io_reset(regs_229_io_reset),
    .io_out(regs_229_io_out),
    .io_enable(regs_229_io_enable)
  );
  FringeFF regs_230 ( // @[RegFile.scala 66:20:@44941.4]
    .clock(regs_230_clock),
    .reset(regs_230_reset),
    .io_in(regs_230_io_in),
    .io_reset(regs_230_io_reset),
    .io_out(regs_230_io_out),
    .io_enable(regs_230_io_enable)
  );
  FringeFF regs_231 ( // @[RegFile.scala 66:20:@44955.4]
    .clock(regs_231_clock),
    .reset(regs_231_reset),
    .io_in(regs_231_io_in),
    .io_reset(regs_231_io_reset),
    .io_out(regs_231_io_out),
    .io_enable(regs_231_io_enable)
  );
  FringeFF regs_232 ( // @[RegFile.scala 66:20:@44969.4]
    .clock(regs_232_clock),
    .reset(regs_232_reset),
    .io_in(regs_232_io_in),
    .io_reset(regs_232_io_reset),
    .io_out(regs_232_io_out),
    .io_enable(regs_232_io_enable)
  );
  FringeFF regs_233 ( // @[RegFile.scala 66:20:@44983.4]
    .clock(regs_233_clock),
    .reset(regs_233_reset),
    .io_in(regs_233_io_in),
    .io_reset(regs_233_io_reset),
    .io_out(regs_233_io_out),
    .io_enable(regs_233_io_enable)
  );
  FringeFF regs_234 ( // @[RegFile.scala 66:20:@44997.4]
    .clock(regs_234_clock),
    .reset(regs_234_reset),
    .io_in(regs_234_io_in),
    .io_reset(regs_234_io_reset),
    .io_out(regs_234_io_out),
    .io_enable(regs_234_io_enable)
  );
  FringeFF regs_235 ( // @[RegFile.scala 66:20:@45011.4]
    .clock(regs_235_clock),
    .reset(regs_235_reset),
    .io_in(regs_235_io_in),
    .io_reset(regs_235_io_reset),
    .io_out(regs_235_io_out),
    .io_enable(regs_235_io_enable)
  );
  FringeFF regs_236 ( // @[RegFile.scala 66:20:@45025.4]
    .clock(regs_236_clock),
    .reset(regs_236_reset),
    .io_in(regs_236_io_in),
    .io_reset(regs_236_io_reset),
    .io_out(regs_236_io_out),
    .io_enable(regs_236_io_enable)
  );
  FringeFF regs_237 ( // @[RegFile.scala 66:20:@45039.4]
    .clock(regs_237_clock),
    .reset(regs_237_reset),
    .io_in(regs_237_io_in),
    .io_reset(regs_237_io_reset),
    .io_out(regs_237_io_out),
    .io_enable(regs_237_io_enable)
  );
  FringeFF regs_238 ( // @[RegFile.scala 66:20:@45053.4]
    .clock(regs_238_clock),
    .reset(regs_238_reset),
    .io_in(regs_238_io_in),
    .io_reset(regs_238_io_reset),
    .io_out(regs_238_io_out),
    .io_enable(regs_238_io_enable)
  );
  FringeFF regs_239 ( // @[RegFile.scala 66:20:@45067.4]
    .clock(regs_239_clock),
    .reset(regs_239_reset),
    .io_in(regs_239_io_in),
    .io_reset(regs_239_io_reset),
    .io_out(regs_239_io_out),
    .io_enable(regs_239_io_enable)
  );
  FringeFF regs_240 ( // @[RegFile.scala 66:20:@45081.4]
    .clock(regs_240_clock),
    .reset(regs_240_reset),
    .io_in(regs_240_io_in),
    .io_reset(regs_240_io_reset),
    .io_out(regs_240_io_out),
    .io_enable(regs_240_io_enable)
  );
  FringeFF regs_241 ( // @[RegFile.scala 66:20:@45095.4]
    .clock(regs_241_clock),
    .reset(regs_241_reset),
    .io_in(regs_241_io_in),
    .io_reset(regs_241_io_reset),
    .io_out(regs_241_io_out),
    .io_enable(regs_241_io_enable)
  );
  FringeFF regs_242 ( // @[RegFile.scala 66:20:@45109.4]
    .clock(regs_242_clock),
    .reset(regs_242_reset),
    .io_in(regs_242_io_in),
    .io_reset(regs_242_io_reset),
    .io_out(regs_242_io_out),
    .io_enable(regs_242_io_enable)
  );
  FringeFF regs_243 ( // @[RegFile.scala 66:20:@45123.4]
    .clock(regs_243_clock),
    .reset(regs_243_reset),
    .io_in(regs_243_io_in),
    .io_reset(regs_243_io_reset),
    .io_out(regs_243_io_out),
    .io_enable(regs_243_io_enable)
  );
  FringeFF regs_244 ( // @[RegFile.scala 66:20:@45137.4]
    .clock(regs_244_clock),
    .reset(regs_244_reset),
    .io_in(regs_244_io_in),
    .io_reset(regs_244_io_reset),
    .io_out(regs_244_io_out),
    .io_enable(regs_244_io_enable)
  );
  FringeFF regs_245 ( // @[RegFile.scala 66:20:@45151.4]
    .clock(regs_245_clock),
    .reset(regs_245_reset),
    .io_in(regs_245_io_in),
    .io_reset(regs_245_io_reset),
    .io_out(regs_245_io_out),
    .io_enable(regs_245_io_enable)
  );
  FringeFF regs_246 ( // @[RegFile.scala 66:20:@45165.4]
    .clock(regs_246_clock),
    .reset(regs_246_reset),
    .io_in(regs_246_io_in),
    .io_reset(regs_246_io_reset),
    .io_out(regs_246_io_out),
    .io_enable(regs_246_io_enable)
  );
  FringeFF regs_247 ( // @[RegFile.scala 66:20:@45179.4]
    .clock(regs_247_clock),
    .reset(regs_247_reset),
    .io_in(regs_247_io_in),
    .io_reset(regs_247_io_reset),
    .io_out(regs_247_io_out),
    .io_enable(regs_247_io_enable)
  );
  FringeFF regs_248 ( // @[RegFile.scala 66:20:@45193.4]
    .clock(regs_248_clock),
    .reset(regs_248_reset),
    .io_in(regs_248_io_in),
    .io_reset(regs_248_io_reset),
    .io_out(regs_248_io_out),
    .io_enable(regs_248_io_enable)
  );
  FringeFF regs_249 ( // @[RegFile.scala 66:20:@45207.4]
    .clock(regs_249_clock),
    .reset(regs_249_reset),
    .io_in(regs_249_io_in),
    .io_reset(regs_249_io_reset),
    .io_out(regs_249_io_out),
    .io_enable(regs_249_io_enable)
  );
  FringeFF regs_250 ( // @[RegFile.scala 66:20:@45221.4]
    .clock(regs_250_clock),
    .reset(regs_250_reset),
    .io_in(regs_250_io_in),
    .io_reset(regs_250_io_reset),
    .io_out(regs_250_io_out),
    .io_enable(regs_250_io_enable)
  );
  FringeFF regs_251 ( // @[RegFile.scala 66:20:@45235.4]
    .clock(regs_251_clock),
    .reset(regs_251_reset),
    .io_in(regs_251_io_in),
    .io_reset(regs_251_io_reset),
    .io_out(regs_251_io_out),
    .io_enable(regs_251_io_enable)
  );
  FringeFF regs_252 ( // @[RegFile.scala 66:20:@45249.4]
    .clock(regs_252_clock),
    .reset(regs_252_reset),
    .io_in(regs_252_io_in),
    .io_reset(regs_252_io_reset),
    .io_out(regs_252_io_out),
    .io_enable(regs_252_io_enable)
  );
  FringeFF regs_253 ( // @[RegFile.scala 66:20:@45263.4]
    .clock(regs_253_clock),
    .reset(regs_253_reset),
    .io_in(regs_253_io_in),
    .io_reset(regs_253_io_reset),
    .io_out(regs_253_io_out),
    .io_enable(regs_253_io_enable)
  );
  FringeFF regs_254 ( // @[RegFile.scala 66:20:@45277.4]
    .clock(regs_254_clock),
    .reset(regs_254_reset),
    .io_in(regs_254_io_in),
    .io_reset(regs_254_io_reset),
    .io_out(regs_254_io_out),
    .io_enable(regs_254_io_enable)
  );
  FringeFF regs_255 ( // @[RegFile.scala 66:20:@45291.4]
    .clock(regs_255_clock),
    .reset(regs_255_reset),
    .io_in(regs_255_io_in),
    .io_reset(regs_255_io_reset),
    .io_out(regs_255_io_out),
    .io_enable(regs_255_io_enable)
  );
  FringeFF regs_256 ( // @[RegFile.scala 66:20:@45305.4]
    .clock(regs_256_clock),
    .reset(regs_256_reset),
    .io_in(regs_256_io_in),
    .io_reset(regs_256_io_reset),
    .io_out(regs_256_io_out),
    .io_enable(regs_256_io_enable)
  );
  FringeFF regs_257 ( // @[RegFile.scala 66:20:@45319.4]
    .clock(regs_257_clock),
    .reset(regs_257_reset),
    .io_in(regs_257_io_in),
    .io_reset(regs_257_io_reset),
    .io_out(regs_257_io_out),
    .io_enable(regs_257_io_enable)
  );
  FringeFF regs_258 ( // @[RegFile.scala 66:20:@45333.4]
    .clock(regs_258_clock),
    .reset(regs_258_reset),
    .io_in(regs_258_io_in),
    .io_reset(regs_258_io_reset),
    .io_out(regs_258_io_out),
    .io_enable(regs_258_io_enable)
  );
  FringeFF regs_259 ( // @[RegFile.scala 66:20:@45347.4]
    .clock(regs_259_clock),
    .reset(regs_259_reset),
    .io_in(regs_259_io_in),
    .io_reset(regs_259_io_reset),
    .io_out(regs_259_io_out),
    .io_enable(regs_259_io_enable)
  );
  FringeFF regs_260 ( // @[RegFile.scala 66:20:@45361.4]
    .clock(regs_260_clock),
    .reset(regs_260_reset),
    .io_in(regs_260_io_in),
    .io_reset(regs_260_io_reset),
    .io_out(regs_260_io_out),
    .io_enable(regs_260_io_enable)
  );
  FringeFF regs_261 ( // @[RegFile.scala 66:20:@45375.4]
    .clock(regs_261_clock),
    .reset(regs_261_reset),
    .io_in(regs_261_io_in),
    .io_reset(regs_261_io_reset),
    .io_out(regs_261_io_out),
    .io_enable(regs_261_io_enable)
  );
  FringeFF regs_262 ( // @[RegFile.scala 66:20:@45389.4]
    .clock(regs_262_clock),
    .reset(regs_262_reset),
    .io_in(regs_262_io_in),
    .io_reset(regs_262_io_reset),
    .io_out(regs_262_io_out),
    .io_enable(regs_262_io_enable)
  );
  FringeFF regs_263 ( // @[RegFile.scala 66:20:@45403.4]
    .clock(regs_263_clock),
    .reset(regs_263_reset),
    .io_in(regs_263_io_in),
    .io_reset(regs_263_io_reset),
    .io_out(regs_263_io_out),
    .io_enable(regs_263_io_enable)
  );
  FringeFF regs_264 ( // @[RegFile.scala 66:20:@45417.4]
    .clock(regs_264_clock),
    .reset(regs_264_reset),
    .io_in(regs_264_io_in),
    .io_reset(regs_264_io_reset),
    .io_out(regs_264_io_out),
    .io_enable(regs_264_io_enable)
  );
  FringeFF regs_265 ( // @[RegFile.scala 66:20:@45431.4]
    .clock(regs_265_clock),
    .reset(regs_265_reset),
    .io_in(regs_265_io_in),
    .io_reset(regs_265_io_reset),
    .io_out(regs_265_io_out),
    .io_enable(regs_265_io_enable)
  );
  FringeFF regs_266 ( // @[RegFile.scala 66:20:@45445.4]
    .clock(regs_266_clock),
    .reset(regs_266_reset),
    .io_in(regs_266_io_in),
    .io_reset(regs_266_io_reset),
    .io_out(regs_266_io_out),
    .io_enable(regs_266_io_enable)
  );
  FringeFF regs_267 ( // @[RegFile.scala 66:20:@45459.4]
    .clock(regs_267_clock),
    .reset(regs_267_reset),
    .io_in(regs_267_io_in),
    .io_reset(regs_267_io_reset),
    .io_out(regs_267_io_out),
    .io_enable(regs_267_io_enable)
  );
  FringeFF regs_268 ( // @[RegFile.scala 66:20:@45473.4]
    .clock(regs_268_clock),
    .reset(regs_268_reset),
    .io_in(regs_268_io_in),
    .io_reset(regs_268_io_reset),
    .io_out(regs_268_io_out),
    .io_enable(regs_268_io_enable)
  );
  FringeFF regs_269 ( // @[RegFile.scala 66:20:@45487.4]
    .clock(regs_269_clock),
    .reset(regs_269_reset),
    .io_in(regs_269_io_in),
    .io_reset(regs_269_io_reset),
    .io_out(regs_269_io_out),
    .io_enable(regs_269_io_enable)
  );
  FringeFF regs_270 ( // @[RegFile.scala 66:20:@45501.4]
    .clock(regs_270_clock),
    .reset(regs_270_reset),
    .io_in(regs_270_io_in),
    .io_reset(regs_270_io_reset),
    .io_out(regs_270_io_out),
    .io_enable(regs_270_io_enable)
  );
  FringeFF regs_271 ( // @[RegFile.scala 66:20:@45515.4]
    .clock(regs_271_clock),
    .reset(regs_271_reset),
    .io_in(regs_271_io_in),
    .io_reset(regs_271_io_reset),
    .io_out(regs_271_io_out),
    .io_enable(regs_271_io_enable)
  );
  FringeFF regs_272 ( // @[RegFile.scala 66:20:@45529.4]
    .clock(regs_272_clock),
    .reset(regs_272_reset),
    .io_in(regs_272_io_in),
    .io_reset(regs_272_io_reset),
    .io_out(regs_272_io_out),
    .io_enable(regs_272_io_enable)
  );
  FringeFF regs_273 ( // @[RegFile.scala 66:20:@45543.4]
    .clock(regs_273_clock),
    .reset(regs_273_reset),
    .io_in(regs_273_io_in),
    .io_reset(regs_273_io_reset),
    .io_out(regs_273_io_out),
    .io_enable(regs_273_io_enable)
  );
  FringeFF regs_274 ( // @[RegFile.scala 66:20:@45557.4]
    .clock(regs_274_clock),
    .reset(regs_274_reset),
    .io_in(regs_274_io_in),
    .io_reset(regs_274_io_reset),
    .io_out(regs_274_io_out),
    .io_enable(regs_274_io_enable)
  );
  FringeFF regs_275 ( // @[RegFile.scala 66:20:@45571.4]
    .clock(regs_275_clock),
    .reset(regs_275_reset),
    .io_in(regs_275_io_in),
    .io_reset(regs_275_io_reset),
    .io_out(regs_275_io_out),
    .io_enable(regs_275_io_enable)
  );
  FringeFF regs_276 ( // @[RegFile.scala 66:20:@45585.4]
    .clock(regs_276_clock),
    .reset(regs_276_reset),
    .io_in(regs_276_io_in),
    .io_reset(regs_276_io_reset),
    .io_out(regs_276_io_out),
    .io_enable(regs_276_io_enable)
  );
  FringeFF regs_277 ( // @[RegFile.scala 66:20:@45599.4]
    .clock(regs_277_clock),
    .reset(regs_277_reset),
    .io_in(regs_277_io_in),
    .io_reset(regs_277_io_reset),
    .io_out(regs_277_io_out),
    .io_enable(regs_277_io_enable)
  );
  FringeFF regs_278 ( // @[RegFile.scala 66:20:@45613.4]
    .clock(regs_278_clock),
    .reset(regs_278_reset),
    .io_in(regs_278_io_in),
    .io_reset(regs_278_io_reset),
    .io_out(regs_278_io_out),
    .io_enable(regs_278_io_enable)
  );
  FringeFF regs_279 ( // @[RegFile.scala 66:20:@45627.4]
    .clock(regs_279_clock),
    .reset(regs_279_reset),
    .io_in(regs_279_io_in),
    .io_reset(regs_279_io_reset),
    .io_out(regs_279_io_out),
    .io_enable(regs_279_io_enable)
  );
  FringeFF regs_280 ( // @[RegFile.scala 66:20:@45641.4]
    .clock(regs_280_clock),
    .reset(regs_280_reset),
    .io_in(regs_280_io_in),
    .io_reset(regs_280_io_reset),
    .io_out(regs_280_io_out),
    .io_enable(regs_280_io_enable)
  );
  FringeFF regs_281 ( // @[RegFile.scala 66:20:@45655.4]
    .clock(regs_281_clock),
    .reset(regs_281_reset),
    .io_in(regs_281_io_in),
    .io_reset(regs_281_io_reset),
    .io_out(regs_281_io_out),
    .io_enable(regs_281_io_enable)
  );
  FringeFF regs_282 ( // @[RegFile.scala 66:20:@45669.4]
    .clock(regs_282_clock),
    .reset(regs_282_reset),
    .io_in(regs_282_io_in),
    .io_reset(regs_282_io_reset),
    .io_out(regs_282_io_out),
    .io_enable(regs_282_io_enable)
  );
  FringeFF regs_283 ( // @[RegFile.scala 66:20:@45683.4]
    .clock(regs_283_clock),
    .reset(regs_283_reset),
    .io_in(regs_283_io_in),
    .io_reset(regs_283_io_reset),
    .io_out(regs_283_io_out),
    .io_enable(regs_283_io_enable)
  );
  FringeFF regs_284 ( // @[RegFile.scala 66:20:@45697.4]
    .clock(regs_284_clock),
    .reset(regs_284_reset),
    .io_in(regs_284_io_in),
    .io_reset(regs_284_io_reset),
    .io_out(regs_284_io_out),
    .io_enable(regs_284_io_enable)
  );
  FringeFF regs_285 ( // @[RegFile.scala 66:20:@45711.4]
    .clock(regs_285_clock),
    .reset(regs_285_reset),
    .io_in(regs_285_io_in),
    .io_reset(regs_285_io_reset),
    .io_out(regs_285_io_out),
    .io_enable(regs_285_io_enable)
  );
  FringeFF regs_286 ( // @[RegFile.scala 66:20:@45725.4]
    .clock(regs_286_clock),
    .reset(regs_286_reset),
    .io_in(regs_286_io_in),
    .io_reset(regs_286_io_reset),
    .io_out(regs_286_io_out),
    .io_enable(regs_286_io_enable)
  );
  FringeFF regs_287 ( // @[RegFile.scala 66:20:@45739.4]
    .clock(regs_287_clock),
    .reset(regs_287_reset),
    .io_in(regs_287_io_in),
    .io_reset(regs_287_io_reset),
    .io_out(regs_287_io_out),
    .io_enable(regs_287_io_enable)
  );
  FringeFF regs_288 ( // @[RegFile.scala 66:20:@45753.4]
    .clock(regs_288_clock),
    .reset(regs_288_reset),
    .io_in(regs_288_io_in),
    .io_reset(regs_288_io_reset),
    .io_out(regs_288_io_out),
    .io_enable(regs_288_io_enable)
  );
  FringeFF regs_289 ( // @[RegFile.scala 66:20:@45767.4]
    .clock(regs_289_clock),
    .reset(regs_289_reset),
    .io_in(regs_289_io_in),
    .io_reset(regs_289_io_reset),
    .io_out(regs_289_io_out),
    .io_enable(regs_289_io_enable)
  );
  FringeFF regs_290 ( // @[RegFile.scala 66:20:@45781.4]
    .clock(regs_290_clock),
    .reset(regs_290_reset),
    .io_in(regs_290_io_in),
    .io_reset(regs_290_io_reset),
    .io_out(regs_290_io_out),
    .io_enable(regs_290_io_enable)
  );
  FringeFF regs_291 ( // @[RegFile.scala 66:20:@45795.4]
    .clock(regs_291_clock),
    .reset(regs_291_reset),
    .io_in(regs_291_io_in),
    .io_reset(regs_291_io_reset),
    .io_out(regs_291_io_out),
    .io_enable(regs_291_io_enable)
  );
  FringeFF regs_292 ( // @[RegFile.scala 66:20:@45809.4]
    .clock(regs_292_clock),
    .reset(regs_292_reset),
    .io_in(regs_292_io_in),
    .io_reset(regs_292_io_reset),
    .io_out(regs_292_io_out),
    .io_enable(regs_292_io_enable)
  );
  FringeFF regs_293 ( // @[RegFile.scala 66:20:@45823.4]
    .clock(regs_293_clock),
    .reset(regs_293_reset),
    .io_in(regs_293_io_in),
    .io_reset(regs_293_io_reset),
    .io_out(regs_293_io_out),
    .io_enable(regs_293_io_enable)
  );
  FringeFF regs_294 ( // @[RegFile.scala 66:20:@45837.4]
    .clock(regs_294_clock),
    .reset(regs_294_reset),
    .io_in(regs_294_io_in),
    .io_reset(regs_294_io_reset),
    .io_out(regs_294_io_out),
    .io_enable(regs_294_io_enable)
  );
  FringeFF regs_295 ( // @[RegFile.scala 66:20:@45851.4]
    .clock(regs_295_clock),
    .reset(regs_295_reset),
    .io_in(regs_295_io_in),
    .io_reset(regs_295_io_reset),
    .io_out(regs_295_io_out),
    .io_enable(regs_295_io_enable)
  );
  FringeFF regs_296 ( // @[RegFile.scala 66:20:@45865.4]
    .clock(regs_296_clock),
    .reset(regs_296_reset),
    .io_in(regs_296_io_in),
    .io_reset(regs_296_io_reset),
    .io_out(regs_296_io_out),
    .io_enable(regs_296_io_enable)
  );
  FringeFF regs_297 ( // @[RegFile.scala 66:20:@45879.4]
    .clock(regs_297_clock),
    .reset(regs_297_reset),
    .io_in(regs_297_io_in),
    .io_reset(regs_297_io_reset),
    .io_out(regs_297_io_out),
    .io_enable(regs_297_io_enable)
  );
  FringeFF regs_298 ( // @[RegFile.scala 66:20:@45893.4]
    .clock(regs_298_clock),
    .reset(regs_298_reset),
    .io_in(regs_298_io_in),
    .io_reset(regs_298_io_reset),
    .io_out(regs_298_io_out),
    .io_enable(regs_298_io_enable)
  );
  FringeFF regs_299 ( // @[RegFile.scala 66:20:@45907.4]
    .clock(regs_299_clock),
    .reset(regs_299_reset),
    .io_in(regs_299_io_in),
    .io_reset(regs_299_io_reset),
    .io_out(regs_299_io_out),
    .io_enable(regs_299_io_enable)
  );
  FringeFF regs_300 ( // @[RegFile.scala 66:20:@45921.4]
    .clock(regs_300_clock),
    .reset(regs_300_reset),
    .io_in(regs_300_io_in),
    .io_reset(regs_300_io_reset),
    .io_out(regs_300_io_out),
    .io_enable(regs_300_io_enable)
  );
  FringeFF regs_301 ( // @[RegFile.scala 66:20:@45935.4]
    .clock(regs_301_clock),
    .reset(regs_301_reset),
    .io_in(regs_301_io_in),
    .io_reset(regs_301_io_reset),
    .io_out(regs_301_io_out),
    .io_enable(regs_301_io_enable)
  );
  FringeFF regs_302 ( // @[RegFile.scala 66:20:@45949.4]
    .clock(regs_302_clock),
    .reset(regs_302_reset),
    .io_in(regs_302_io_in),
    .io_reset(regs_302_io_reset),
    .io_out(regs_302_io_out),
    .io_enable(regs_302_io_enable)
  );
  FringeFF regs_303 ( // @[RegFile.scala 66:20:@45963.4]
    .clock(regs_303_clock),
    .reset(regs_303_reset),
    .io_in(regs_303_io_in),
    .io_reset(regs_303_io_reset),
    .io_out(regs_303_io_out),
    .io_enable(regs_303_io_enable)
  );
  FringeFF regs_304 ( // @[RegFile.scala 66:20:@45977.4]
    .clock(regs_304_clock),
    .reset(regs_304_reset),
    .io_in(regs_304_io_in),
    .io_reset(regs_304_io_reset),
    .io_out(regs_304_io_out),
    .io_enable(regs_304_io_enable)
  );
  FringeFF regs_305 ( // @[RegFile.scala 66:20:@45991.4]
    .clock(regs_305_clock),
    .reset(regs_305_reset),
    .io_in(regs_305_io_in),
    .io_reset(regs_305_io_reset),
    .io_out(regs_305_io_out),
    .io_enable(regs_305_io_enable)
  );
  FringeFF regs_306 ( // @[RegFile.scala 66:20:@46005.4]
    .clock(regs_306_clock),
    .reset(regs_306_reset),
    .io_in(regs_306_io_in),
    .io_reset(regs_306_io_reset),
    .io_out(regs_306_io_out),
    .io_enable(regs_306_io_enable)
  );
  FringeFF regs_307 ( // @[RegFile.scala 66:20:@46019.4]
    .clock(regs_307_clock),
    .reset(regs_307_reset),
    .io_in(regs_307_io_in),
    .io_reset(regs_307_io_reset),
    .io_out(regs_307_io_out),
    .io_enable(regs_307_io_enable)
  );
  FringeFF regs_308 ( // @[RegFile.scala 66:20:@46033.4]
    .clock(regs_308_clock),
    .reset(regs_308_reset),
    .io_in(regs_308_io_in),
    .io_reset(regs_308_io_reset),
    .io_out(regs_308_io_out),
    .io_enable(regs_308_io_enable)
  );
  FringeFF regs_309 ( // @[RegFile.scala 66:20:@46047.4]
    .clock(regs_309_clock),
    .reset(regs_309_reset),
    .io_in(regs_309_io_in),
    .io_reset(regs_309_io_reset),
    .io_out(regs_309_io_out),
    .io_enable(regs_309_io_enable)
  );
  FringeFF regs_310 ( // @[RegFile.scala 66:20:@46061.4]
    .clock(regs_310_clock),
    .reset(regs_310_reset),
    .io_in(regs_310_io_in),
    .io_reset(regs_310_io_reset),
    .io_out(regs_310_io_out),
    .io_enable(regs_310_io_enable)
  );
  FringeFF regs_311 ( // @[RegFile.scala 66:20:@46075.4]
    .clock(regs_311_clock),
    .reset(regs_311_reset),
    .io_in(regs_311_io_in),
    .io_reset(regs_311_io_reset),
    .io_out(regs_311_io_out),
    .io_enable(regs_311_io_enable)
  );
  FringeFF regs_312 ( // @[RegFile.scala 66:20:@46089.4]
    .clock(regs_312_clock),
    .reset(regs_312_reset),
    .io_in(regs_312_io_in),
    .io_reset(regs_312_io_reset),
    .io_out(regs_312_io_out),
    .io_enable(regs_312_io_enable)
  );
  FringeFF regs_313 ( // @[RegFile.scala 66:20:@46103.4]
    .clock(regs_313_clock),
    .reset(regs_313_reset),
    .io_in(regs_313_io_in),
    .io_reset(regs_313_io_reset),
    .io_out(regs_313_io_out),
    .io_enable(regs_313_io_enable)
  );
  FringeFF regs_314 ( // @[RegFile.scala 66:20:@46117.4]
    .clock(regs_314_clock),
    .reset(regs_314_reset),
    .io_in(regs_314_io_in),
    .io_reset(regs_314_io_reset),
    .io_out(regs_314_io_out),
    .io_enable(regs_314_io_enable)
  );
  FringeFF regs_315 ( // @[RegFile.scala 66:20:@46131.4]
    .clock(regs_315_clock),
    .reset(regs_315_reset),
    .io_in(regs_315_io_in),
    .io_reset(regs_315_io_reset),
    .io_out(regs_315_io_out),
    .io_enable(regs_315_io_enable)
  );
  FringeFF regs_316 ( // @[RegFile.scala 66:20:@46145.4]
    .clock(regs_316_clock),
    .reset(regs_316_reset),
    .io_in(regs_316_io_in),
    .io_reset(regs_316_io_reset),
    .io_out(regs_316_io_out),
    .io_enable(regs_316_io_enable)
  );
  FringeFF regs_317 ( // @[RegFile.scala 66:20:@46159.4]
    .clock(regs_317_clock),
    .reset(regs_317_reset),
    .io_in(regs_317_io_in),
    .io_reset(regs_317_io_reset),
    .io_out(regs_317_io_out),
    .io_enable(regs_317_io_enable)
  );
  FringeFF regs_318 ( // @[RegFile.scala 66:20:@46173.4]
    .clock(regs_318_clock),
    .reset(regs_318_reset),
    .io_in(regs_318_io_in),
    .io_reset(regs_318_io_reset),
    .io_out(regs_318_io_out),
    .io_enable(regs_318_io_enable)
  );
  FringeFF regs_319 ( // @[RegFile.scala 66:20:@46187.4]
    .clock(regs_319_clock),
    .reset(regs_319_reset),
    .io_in(regs_319_io_in),
    .io_reset(regs_319_io_reset),
    .io_out(regs_319_io_out),
    .io_enable(regs_319_io_enable)
  );
  FringeFF regs_320 ( // @[RegFile.scala 66:20:@46201.4]
    .clock(regs_320_clock),
    .reset(regs_320_reset),
    .io_in(regs_320_io_in),
    .io_reset(regs_320_io_reset),
    .io_out(regs_320_io_out),
    .io_enable(regs_320_io_enable)
  );
  FringeFF regs_321 ( // @[RegFile.scala 66:20:@46215.4]
    .clock(regs_321_clock),
    .reset(regs_321_reset),
    .io_in(regs_321_io_in),
    .io_reset(regs_321_io_reset),
    .io_out(regs_321_io_out),
    .io_enable(regs_321_io_enable)
  );
  FringeFF regs_322 ( // @[RegFile.scala 66:20:@46229.4]
    .clock(regs_322_clock),
    .reset(regs_322_reset),
    .io_in(regs_322_io_in),
    .io_reset(regs_322_io_reset),
    .io_out(regs_322_io_out),
    .io_enable(regs_322_io_enable)
  );
  FringeFF regs_323 ( // @[RegFile.scala 66:20:@46243.4]
    .clock(regs_323_clock),
    .reset(regs_323_reset),
    .io_in(regs_323_io_in),
    .io_reset(regs_323_io_reset),
    .io_out(regs_323_io_out),
    .io_enable(regs_323_io_enable)
  );
  FringeFF regs_324 ( // @[RegFile.scala 66:20:@46257.4]
    .clock(regs_324_clock),
    .reset(regs_324_reset),
    .io_in(regs_324_io_in),
    .io_reset(regs_324_io_reset),
    .io_out(regs_324_io_out),
    .io_enable(regs_324_io_enable)
  );
  FringeFF regs_325 ( // @[RegFile.scala 66:20:@46271.4]
    .clock(regs_325_clock),
    .reset(regs_325_reset),
    .io_in(regs_325_io_in),
    .io_reset(regs_325_io_reset),
    .io_out(regs_325_io_out),
    .io_enable(regs_325_io_enable)
  );
  FringeFF regs_326 ( // @[RegFile.scala 66:20:@46285.4]
    .clock(regs_326_clock),
    .reset(regs_326_reset),
    .io_in(regs_326_io_in),
    .io_reset(regs_326_io_reset),
    .io_out(regs_326_io_out),
    .io_enable(regs_326_io_enable)
  );
  FringeFF regs_327 ( // @[RegFile.scala 66:20:@46299.4]
    .clock(regs_327_clock),
    .reset(regs_327_reset),
    .io_in(regs_327_io_in),
    .io_reset(regs_327_io_reset),
    .io_out(regs_327_io_out),
    .io_enable(regs_327_io_enable)
  );
  FringeFF regs_328 ( // @[RegFile.scala 66:20:@46313.4]
    .clock(regs_328_clock),
    .reset(regs_328_reset),
    .io_in(regs_328_io_in),
    .io_reset(regs_328_io_reset),
    .io_out(regs_328_io_out),
    .io_enable(regs_328_io_enable)
  );
  FringeFF regs_329 ( // @[RegFile.scala 66:20:@46327.4]
    .clock(regs_329_clock),
    .reset(regs_329_reset),
    .io_in(regs_329_io_in),
    .io_reset(regs_329_io_reset),
    .io_out(regs_329_io_out),
    .io_enable(regs_329_io_enable)
  );
  FringeFF regs_330 ( // @[RegFile.scala 66:20:@46341.4]
    .clock(regs_330_clock),
    .reset(regs_330_reset),
    .io_in(regs_330_io_in),
    .io_reset(regs_330_io_reset),
    .io_out(regs_330_io_out),
    .io_enable(regs_330_io_enable)
  );
  FringeFF regs_331 ( // @[RegFile.scala 66:20:@46355.4]
    .clock(regs_331_clock),
    .reset(regs_331_reset),
    .io_in(regs_331_io_in),
    .io_reset(regs_331_io_reset),
    .io_out(regs_331_io_out),
    .io_enable(regs_331_io_enable)
  );
  FringeFF regs_332 ( // @[RegFile.scala 66:20:@46369.4]
    .clock(regs_332_clock),
    .reset(regs_332_reset),
    .io_in(regs_332_io_in),
    .io_reset(regs_332_io_reset),
    .io_out(regs_332_io_out),
    .io_enable(regs_332_io_enable)
  );
  FringeFF regs_333 ( // @[RegFile.scala 66:20:@46383.4]
    .clock(regs_333_clock),
    .reset(regs_333_reset),
    .io_in(regs_333_io_in),
    .io_reset(regs_333_io_reset),
    .io_out(regs_333_io_out),
    .io_enable(regs_333_io_enable)
  );
  FringeFF regs_334 ( // @[RegFile.scala 66:20:@46397.4]
    .clock(regs_334_clock),
    .reset(regs_334_reset),
    .io_in(regs_334_io_in),
    .io_reset(regs_334_io_reset),
    .io_out(regs_334_io_out),
    .io_enable(regs_334_io_enable)
  );
  FringeFF regs_335 ( // @[RegFile.scala 66:20:@46411.4]
    .clock(regs_335_clock),
    .reset(regs_335_reset),
    .io_in(regs_335_io_in),
    .io_reset(regs_335_io_reset),
    .io_out(regs_335_io_out),
    .io_enable(regs_335_io_enable)
  );
  FringeFF regs_336 ( // @[RegFile.scala 66:20:@46425.4]
    .clock(regs_336_clock),
    .reset(regs_336_reset),
    .io_in(regs_336_io_in),
    .io_reset(regs_336_io_reset),
    .io_out(regs_336_io_out),
    .io_enable(regs_336_io_enable)
  );
  FringeFF regs_337 ( // @[RegFile.scala 66:20:@46439.4]
    .clock(regs_337_clock),
    .reset(regs_337_reset),
    .io_in(regs_337_io_in),
    .io_reset(regs_337_io_reset),
    .io_out(regs_337_io_out),
    .io_enable(regs_337_io_enable)
  );
  FringeFF regs_338 ( // @[RegFile.scala 66:20:@46453.4]
    .clock(regs_338_clock),
    .reset(regs_338_reset),
    .io_in(regs_338_io_in),
    .io_reset(regs_338_io_reset),
    .io_out(regs_338_io_out),
    .io_enable(regs_338_io_enable)
  );
  FringeFF regs_339 ( // @[RegFile.scala 66:20:@46467.4]
    .clock(regs_339_clock),
    .reset(regs_339_reset),
    .io_in(regs_339_io_in),
    .io_reset(regs_339_io_reset),
    .io_out(regs_339_io_out),
    .io_enable(regs_339_io_enable)
  );
  FringeFF regs_340 ( // @[RegFile.scala 66:20:@46481.4]
    .clock(regs_340_clock),
    .reset(regs_340_reset),
    .io_in(regs_340_io_in),
    .io_reset(regs_340_io_reset),
    .io_out(regs_340_io_out),
    .io_enable(regs_340_io_enable)
  );
  FringeFF regs_341 ( // @[RegFile.scala 66:20:@46495.4]
    .clock(regs_341_clock),
    .reset(regs_341_reset),
    .io_in(regs_341_io_in),
    .io_reset(regs_341_io_reset),
    .io_out(regs_341_io_out),
    .io_enable(regs_341_io_enable)
  );
  FringeFF regs_342 ( // @[RegFile.scala 66:20:@46509.4]
    .clock(regs_342_clock),
    .reset(regs_342_reset),
    .io_in(regs_342_io_in),
    .io_reset(regs_342_io_reset),
    .io_out(regs_342_io_out),
    .io_enable(regs_342_io_enable)
  );
  FringeFF regs_343 ( // @[RegFile.scala 66:20:@46523.4]
    .clock(regs_343_clock),
    .reset(regs_343_reset),
    .io_in(regs_343_io_in),
    .io_reset(regs_343_io_reset),
    .io_out(regs_343_io_out),
    .io_enable(regs_343_io_enable)
  );
  FringeFF regs_344 ( // @[RegFile.scala 66:20:@46537.4]
    .clock(regs_344_clock),
    .reset(regs_344_reset),
    .io_in(regs_344_io_in),
    .io_reset(regs_344_io_reset),
    .io_out(regs_344_io_out),
    .io_enable(regs_344_io_enable)
  );
  FringeFF regs_345 ( // @[RegFile.scala 66:20:@46551.4]
    .clock(regs_345_clock),
    .reset(regs_345_reset),
    .io_in(regs_345_io_in),
    .io_reset(regs_345_io_reset),
    .io_out(regs_345_io_out),
    .io_enable(regs_345_io_enable)
  );
  FringeFF regs_346 ( // @[RegFile.scala 66:20:@46565.4]
    .clock(regs_346_clock),
    .reset(regs_346_reset),
    .io_in(regs_346_io_in),
    .io_reset(regs_346_io_reset),
    .io_out(regs_346_io_out),
    .io_enable(regs_346_io_enable)
  );
  FringeFF regs_347 ( // @[RegFile.scala 66:20:@46579.4]
    .clock(regs_347_clock),
    .reset(regs_347_reset),
    .io_in(regs_347_io_in),
    .io_reset(regs_347_io_reset),
    .io_out(regs_347_io_out),
    .io_enable(regs_347_io_enable)
  );
  FringeFF regs_348 ( // @[RegFile.scala 66:20:@46593.4]
    .clock(regs_348_clock),
    .reset(regs_348_reset),
    .io_in(regs_348_io_in),
    .io_reset(regs_348_io_reset),
    .io_out(regs_348_io_out),
    .io_enable(regs_348_io_enable)
  );
  FringeFF regs_349 ( // @[RegFile.scala 66:20:@46607.4]
    .clock(regs_349_clock),
    .reset(regs_349_reset),
    .io_in(regs_349_io_in),
    .io_reset(regs_349_io_reset),
    .io_out(regs_349_io_out),
    .io_enable(regs_349_io_enable)
  );
  FringeFF regs_350 ( // @[RegFile.scala 66:20:@46621.4]
    .clock(regs_350_clock),
    .reset(regs_350_reset),
    .io_in(regs_350_io_in),
    .io_reset(regs_350_io_reset),
    .io_out(regs_350_io_out),
    .io_enable(regs_350_io_enable)
  );
  FringeFF regs_351 ( // @[RegFile.scala 66:20:@46635.4]
    .clock(regs_351_clock),
    .reset(regs_351_reset),
    .io_in(regs_351_io_in),
    .io_reset(regs_351_io_reset),
    .io_out(regs_351_io_out),
    .io_enable(regs_351_io_enable)
  );
  FringeFF regs_352 ( // @[RegFile.scala 66:20:@46649.4]
    .clock(regs_352_clock),
    .reset(regs_352_reset),
    .io_in(regs_352_io_in),
    .io_reset(regs_352_io_reset),
    .io_out(regs_352_io_out),
    .io_enable(regs_352_io_enable)
  );
  FringeFF regs_353 ( // @[RegFile.scala 66:20:@46663.4]
    .clock(regs_353_clock),
    .reset(regs_353_reset),
    .io_in(regs_353_io_in),
    .io_reset(regs_353_io_reset),
    .io_out(regs_353_io_out),
    .io_enable(regs_353_io_enable)
  );
  FringeFF regs_354 ( // @[RegFile.scala 66:20:@46677.4]
    .clock(regs_354_clock),
    .reset(regs_354_reset),
    .io_in(regs_354_io_in),
    .io_reset(regs_354_io_reset),
    .io_out(regs_354_io_out),
    .io_enable(regs_354_io_enable)
  );
  FringeFF regs_355 ( // @[RegFile.scala 66:20:@46691.4]
    .clock(regs_355_clock),
    .reset(regs_355_reset),
    .io_in(regs_355_io_in),
    .io_reset(regs_355_io_reset),
    .io_out(regs_355_io_out),
    .io_enable(regs_355_io_enable)
  );
  FringeFF regs_356 ( // @[RegFile.scala 66:20:@46705.4]
    .clock(regs_356_clock),
    .reset(regs_356_reset),
    .io_in(regs_356_io_in),
    .io_reset(regs_356_io_reset),
    .io_out(regs_356_io_out),
    .io_enable(regs_356_io_enable)
  );
  FringeFF regs_357 ( // @[RegFile.scala 66:20:@46719.4]
    .clock(regs_357_clock),
    .reset(regs_357_reset),
    .io_in(regs_357_io_in),
    .io_reset(regs_357_io_reset),
    .io_out(regs_357_io_out),
    .io_enable(regs_357_io_enable)
  );
  FringeFF regs_358 ( // @[RegFile.scala 66:20:@46733.4]
    .clock(regs_358_clock),
    .reset(regs_358_reset),
    .io_in(regs_358_io_in),
    .io_reset(regs_358_io_reset),
    .io_out(regs_358_io_out),
    .io_enable(regs_358_io_enable)
  );
  FringeFF regs_359 ( // @[RegFile.scala 66:20:@46747.4]
    .clock(regs_359_clock),
    .reset(regs_359_reset),
    .io_in(regs_359_io_in),
    .io_reset(regs_359_io_reset),
    .io_out(regs_359_io_out),
    .io_enable(regs_359_io_enable)
  );
  FringeFF regs_360 ( // @[RegFile.scala 66:20:@46761.4]
    .clock(regs_360_clock),
    .reset(regs_360_reset),
    .io_in(regs_360_io_in),
    .io_reset(regs_360_io_reset),
    .io_out(regs_360_io_out),
    .io_enable(regs_360_io_enable)
  );
  FringeFF regs_361 ( // @[RegFile.scala 66:20:@46775.4]
    .clock(regs_361_clock),
    .reset(regs_361_reset),
    .io_in(regs_361_io_in),
    .io_reset(regs_361_io_reset),
    .io_out(regs_361_io_out),
    .io_enable(regs_361_io_enable)
  );
  FringeFF regs_362 ( // @[RegFile.scala 66:20:@46789.4]
    .clock(regs_362_clock),
    .reset(regs_362_reset),
    .io_in(regs_362_io_in),
    .io_reset(regs_362_io_reset),
    .io_out(regs_362_io_out),
    .io_enable(regs_362_io_enable)
  );
  FringeFF regs_363 ( // @[RegFile.scala 66:20:@46803.4]
    .clock(regs_363_clock),
    .reset(regs_363_reset),
    .io_in(regs_363_io_in),
    .io_reset(regs_363_io_reset),
    .io_out(regs_363_io_out),
    .io_enable(regs_363_io_enable)
  );
  FringeFF regs_364 ( // @[RegFile.scala 66:20:@46817.4]
    .clock(regs_364_clock),
    .reset(regs_364_reset),
    .io_in(regs_364_io_in),
    .io_reset(regs_364_io_reset),
    .io_out(regs_364_io_out),
    .io_enable(regs_364_io_enable)
  );
  FringeFF regs_365 ( // @[RegFile.scala 66:20:@46831.4]
    .clock(regs_365_clock),
    .reset(regs_365_reset),
    .io_in(regs_365_io_in),
    .io_reset(regs_365_io_reset),
    .io_out(regs_365_io_out),
    .io_enable(regs_365_io_enable)
  );
  FringeFF regs_366 ( // @[RegFile.scala 66:20:@46845.4]
    .clock(regs_366_clock),
    .reset(regs_366_reset),
    .io_in(regs_366_io_in),
    .io_reset(regs_366_io_reset),
    .io_out(regs_366_io_out),
    .io_enable(regs_366_io_enable)
  );
  FringeFF regs_367 ( // @[RegFile.scala 66:20:@46859.4]
    .clock(regs_367_clock),
    .reset(regs_367_reset),
    .io_in(regs_367_io_in),
    .io_reset(regs_367_io_reset),
    .io_out(regs_367_io_out),
    .io_enable(regs_367_io_enable)
  );
  FringeFF regs_368 ( // @[RegFile.scala 66:20:@46873.4]
    .clock(regs_368_clock),
    .reset(regs_368_reset),
    .io_in(regs_368_io_in),
    .io_reset(regs_368_io_reset),
    .io_out(regs_368_io_out),
    .io_enable(regs_368_io_enable)
  );
  FringeFF regs_369 ( // @[RegFile.scala 66:20:@46887.4]
    .clock(regs_369_clock),
    .reset(regs_369_reset),
    .io_in(regs_369_io_in),
    .io_reset(regs_369_io_reset),
    .io_out(regs_369_io_out),
    .io_enable(regs_369_io_enable)
  );
  FringeFF regs_370 ( // @[RegFile.scala 66:20:@46901.4]
    .clock(regs_370_clock),
    .reset(regs_370_reset),
    .io_in(regs_370_io_in),
    .io_reset(regs_370_io_reset),
    .io_out(regs_370_io_out),
    .io_enable(regs_370_io_enable)
  );
  FringeFF regs_371 ( // @[RegFile.scala 66:20:@46915.4]
    .clock(regs_371_clock),
    .reset(regs_371_reset),
    .io_in(regs_371_io_in),
    .io_reset(regs_371_io_reset),
    .io_out(regs_371_io_out),
    .io_enable(regs_371_io_enable)
  );
  FringeFF regs_372 ( // @[RegFile.scala 66:20:@46929.4]
    .clock(regs_372_clock),
    .reset(regs_372_reset),
    .io_in(regs_372_io_in),
    .io_reset(regs_372_io_reset),
    .io_out(regs_372_io_out),
    .io_enable(regs_372_io_enable)
  );
  FringeFF regs_373 ( // @[RegFile.scala 66:20:@46943.4]
    .clock(regs_373_clock),
    .reset(regs_373_reset),
    .io_in(regs_373_io_in),
    .io_reset(regs_373_io_reset),
    .io_out(regs_373_io_out),
    .io_enable(regs_373_io_enable)
  );
  FringeFF regs_374 ( // @[RegFile.scala 66:20:@46957.4]
    .clock(regs_374_clock),
    .reset(regs_374_reset),
    .io_in(regs_374_io_in),
    .io_reset(regs_374_io_reset),
    .io_out(regs_374_io_out),
    .io_enable(regs_374_io_enable)
  );
  FringeFF regs_375 ( // @[RegFile.scala 66:20:@46971.4]
    .clock(regs_375_clock),
    .reset(regs_375_reset),
    .io_in(regs_375_io_in),
    .io_reset(regs_375_io_reset),
    .io_out(regs_375_io_out),
    .io_enable(regs_375_io_enable)
  );
  FringeFF regs_376 ( // @[RegFile.scala 66:20:@46985.4]
    .clock(regs_376_clock),
    .reset(regs_376_reset),
    .io_in(regs_376_io_in),
    .io_reset(regs_376_io_reset),
    .io_out(regs_376_io_out),
    .io_enable(regs_376_io_enable)
  );
  FringeFF regs_377 ( // @[RegFile.scala 66:20:@46999.4]
    .clock(regs_377_clock),
    .reset(regs_377_reset),
    .io_in(regs_377_io_in),
    .io_reset(regs_377_io_reset),
    .io_out(regs_377_io_out),
    .io_enable(regs_377_io_enable)
  );
  FringeFF regs_378 ( // @[RegFile.scala 66:20:@47013.4]
    .clock(regs_378_clock),
    .reset(regs_378_reset),
    .io_in(regs_378_io_in),
    .io_reset(regs_378_io_reset),
    .io_out(regs_378_io_out),
    .io_enable(regs_378_io_enable)
  );
  FringeFF regs_379 ( // @[RegFile.scala 66:20:@47027.4]
    .clock(regs_379_clock),
    .reset(regs_379_reset),
    .io_in(regs_379_io_in),
    .io_reset(regs_379_io_reset),
    .io_out(regs_379_io_out),
    .io_enable(regs_379_io_enable)
  );
  FringeFF regs_380 ( // @[RegFile.scala 66:20:@47041.4]
    .clock(regs_380_clock),
    .reset(regs_380_reset),
    .io_in(regs_380_io_in),
    .io_reset(regs_380_io_reset),
    .io_out(regs_380_io_out),
    .io_enable(regs_380_io_enable)
  );
  FringeFF regs_381 ( // @[RegFile.scala 66:20:@47055.4]
    .clock(regs_381_clock),
    .reset(regs_381_reset),
    .io_in(regs_381_io_in),
    .io_reset(regs_381_io_reset),
    .io_out(regs_381_io_out),
    .io_enable(regs_381_io_enable)
  );
  FringeFF regs_382 ( // @[RegFile.scala 66:20:@47069.4]
    .clock(regs_382_clock),
    .reset(regs_382_reset),
    .io_in(regs_382_io_in),
    .io_reset(regs_382_io_reset),
    .io_out(regs_382_io_out),
    .io_enable(regs_382_io_enable)
  );
  FringeFF regs_383 ( // @[RegFile.scala 66:20:@47083.4]
    .clock(regs_383_clock),
    .reset(regs_383_reset),
    .io_in(regs_383_io_in),
    .io_reset(regs_383_io_reset),
    .io_out(regs_383_io_out),
    .io_enable(regs_383_io_enable)
  );
  FringeFF regs_384 ( // @[RegFile.scala 66:20:@47097.4]
    .clock(regs_384_clock),
    .reset(regs_384_reset),
    .io_in(regs_384_io_in),
    .io_reset(regs_384_io_reset),
    .io_out(regs_384_io_out),
    .io_enable(regs_384_io_enable)
  );
  FringeFF regs_385 ( // @[RegFile.scala 66:20:@47111.4]
    .clock(regs_385_clock),
    .reset(regs_385_reset),
    .io_in(regs_385_io_in),
    .io_reset(regs_385_io_reset),
    .io_out(regs_385_io_out),
    .io_enable(regs_385_io_enable)
  );
  FringeFF regs_386 ( // @[RegFile.scala 66:20:@47125.4]
    .clock(regs_386_clock),
    .reset(regs_386_reset),
    .io_in(regs_386_io_in),
    .io_reset(regs_386_io_reset),
    .io_out(regs_386_io_out),
    .io_enable(regs_386_io_enable)
  );
  FringeFF regs_387 ( // @[RegFile.scala 66:20:@47139.4]
    .clock(regs_387_clock),
    .reset(regs_387_reset),
    .io_in(regs_387_io_in),
    .io_reset(regs_387_io_reset),
    .io_out(regs_387_io_out),
    .io_enable(regs_387_io_enable)
  );
  FringeFF regs_388 ( // @[RegFile.scala 66:20:@47153.4]
    .clock(regs_388_clock),
    .reset(regs_388_reset),
    .io_in(regs_388_io_in),
    .io_reset(regs_388_io_reset),
    .io_out(regs_388_io_out),
    .io_enable(regs_388_io_enable)
  );
  FringeFF regs_389 ( // @[RegFile.scala 66:20:@47167.4]
    .clock(regs_389_clock),
    .reset(regs_389_reset),
    .io_in(regs_389_io_in),
    .io_reset(regs_389_io_reset),
    .io_out(regs_389_io_out),
    .io_enable(regs_389_io_enable)
  );
  FringeFF regs_390 ( // @[RegFile.scala 66:20:@47181.4]
    .clock(regs_390_clock),
    .reset(regs_390_reset),
    .io_in(regs_390_io_in),
    .io_reset(regs_390_io_reset),
    .io_out(regs_390_io_out),
    .io_enable(regs_390_io_enable)
  );
  FringeFF regs_391 ( // @[RegFile.scala 66:20:@47195.4]
    .clock(regs_391_clock),
    .reset(regs_391_reset),
    .io_in(regs_391_io_in),
    .io_reset(regs_391_io_reset),
    .io_out(regs_391_io_out),
    .io_enable(regs_391_io_enable)
  );
  FringeFF regs_392 ( // @[RegFile.scala 66:20:@47209.4]
    .clock(regs_392_clock),
    .reset(regs_392_reset),
    .io_in(regs_392_io_in),
    .io_reset(regs_392_io_reset),
    .io_out(regs_392_io_out),
    .io_enable(regs_392_io_enable)
  );
  FringeFF regs_393 ( // @[RegFile.scala 66:20:@47223.4]
    .clock(regs_393_clock),
    .reset(regs_393_reset),
    .io_in(regs_393_io_in),
    .io_reset(regs_393_io_reset),
    .io_out(regs_393_io_out),
    .io_enable(regs_393_io_enable)
  );
  FringeFF regs_394 ( // @[RegFile.scala 66:20:@47237.4]
    .clock(regs_394_clock),
    .reset(regs_394_reset),
    .io_in(regs_394_io_in),
    .io_reset(regs_394_io_reset),
    .io_out(regs_394_io_out),
    .io_enable(regs_394_io_enable)
  );
  FringeFF regs_395 ( // @[RegFile.scala 66:20:@47251.4]
    .clock(regs_395_clock),
    .reset(regs_395_reset),
    .io_in(regs_395_io_in),
    .io_reset(regs_395_io_reset),
    .io_out(regs_395_io_out),
    .io_enable(regs_395_io_enable)
  );
  FringeFF regs_396 ( // @[RegFile.scala 66:20:@47265.4]
    .clock(regs_396_clock),
    .reset(regs_396_reset),
    .io_in(regs_396_io_in),
    .io_reset(regs_396_io_reset),
    .io_out(regs_396_io_out),
    .io_enable(regs_396_io_enable)
  );
  FringeFF regs_397 ( // @[RegFile.scala 66:20:@47279.4]
    .clock(regs_397_clock),
    .reset(regs_397_reset),
    .io_in(regs_397_io_in),
    .io_reset(regs_397_io_reset),
    .io_out(regs_397_io_out),
    .io_enable(regs_397_io_enable)
  );
  FringeFF regs_398 ( // @[RegFile.scala 66:20:@47293.4]
    .clock(regs_398_clock),
    .reset(regs_398_reset),
    .io_in(regs_398_io_in),
    .io_reset(regs_398_io_reset),
    .io_out(regs_398_io_out),
    .io_enable(regs_398_io_enable)
  );
  FringeFF regs_399 ( // @[RegFile.scala 66:20:@47307.4]
    .clock(regs_399_clock),
    .reset(regs_399_reset),
    .io_in(regs_399_io_in),
    .io_reset(regs_399_io_reset),
    .io_out(regs_399_io_out),
    .io_enable(regs_399_io_enable)
  );
  FringeFF regs_400 ( // @[RegFile.scala 66:20:@47321.4]
    .clock(regs_400_clock),
    .reset(regs_400_reset),
    .io_in(regs_400_io_in),
    .io_reset(regs_400_io_reset),
    .io_out(regs_400_io_out),
    .io_enable(regs_400_io_enable)
  );
  FringeFF regs_401 ( // @[RegFile.scala 66:20:@47335.4]
    .clock(regs_401_clock),
    .reset(regs_401_reset),
    .io_in(regs_401_io_in),
    .io_reset(regs_401_io_reset),
    .io_out(regs_401_io_out),
    .io_enable(regs_401_io_enable)
  );
  FringeFF regs_402 ( // @[RegFile.scala 66:20:@47349.4]
    .clock(regs_402_clock),
    .reset(regs_402_reset),
    .io_in(regs_402_io_in),
    .io_reset(regs_402_io_reset),
    .io_out(regs_402_io_out),
    .io_enable(regs_402_io_enable)
  );
  FringeFF regs_403 ( // @[RegFile.scala 66:20:@47363.4]
    .clock(regs_403_clock),
    .reset(regs_403_reset),
    .io_in(regs_403_io_in),
    .io_reset(regs_403_io_reset),
    .io_out(regs_403_io_out),
    .io_enable(regs_403_io_enable)
  );
  FringeFF regs_404 ( // @[RegFile.scala 66:20:@47377.4]
    .clock(regs_404_clock),
    .reset(regs_404_reset),
    .io_in(regs_404_io_in),
    .io_reset(regs_404_io_reset),
    .io_out(regs_404_io_out),
    .io_enable(regs_404_io_enable)
  );
  FringeFF regs_405 ( // @[RegFile.scala 66:20:@47391.4]
    .clock(regs_405_clock),
    .reset(regs_405_reset),
    .io_in(regs_405_io_in),
    .io_reset(regs_405_io_reset),
    .io_out(regs_405_io_out),
    .io_enable(regs_405_io_enable)
  );
  FringeFF regs_406 ( // @[RegFile.scala 66:20:@47405.4]
    .clock(regs_406_clock),
    .reset(regs_406_reset),
    .io_in(regs_406_io_in),
    .io_reset(regs_406_io_reset),
    .io_out(regs_406_io_out),
    .io_enable(regs_406_io_enable)
  );
  FringeFF regs_407 ( // @[RegFile.scala 66:20:@47419.4]
    .clock(regs_407_clock),
    .reset(regs_407_reset),
    .io_in(regs_407_io_in),
    .io_reset(regs_407_io_reset),
    .io_out(regs_407_io_out),
    .io_enable(regs_407_io_enable)
  );
  FringeFF regs_408 ( // @[RegFile.scala 66:20:@47433.4]
    .clock(regs_408_clock),
    .reset(regs_408_reset),
    .io_in(regs_408_io_in),
    .io_reset(regs_408_io_reset),
    .io_out(regs_408_io_out),
    .io_enable(regs_408_io_enable)
  );
  FringeFF regs_409 ( // @[RegFile.scala 66:20:@47447.4]
    .clock(regs_409_clock),
    .reset(regs_409_reset),
    .io_in(regs_409_io_in),
    .io_reset(regs_409_io_reset),
    .io_out(regs_409_io_out),
    .io_enable(regs_409_io_enable)
  );
  FringeFF regs_410 ( // @[RegFile.scala 66:20:@47461.4]
    .clock(regs_410_clock),
    .reset(regs_410_reset),
    .io_in(regs_410_io_in),
    .io_reset(regs_410_io_reset),
    .io_out(regs_410_io_out),
    .io_enable(regs_410_io_enable)
  );
  FringeFF regs_411 ( // @[RegFile.scala 66:20:@47475.4]
    .clock(regs_411_clock),
    .reset(regs_411_reset),
    .io_in(regs_411_io_in),
    .io_reset(regs_411_io_reset),
    .io_out(regs_411_io_out),
    .io_enable(regs_411_io_enable)
  );
  FringeFF regs_412 ( // @[RegFile.scala 66:20:@47489.4]
    .clock(regs_412_clock),
    .reset(regs_412_reset),
    .io_in(regs_412_io_in),
    .io_reset(regs_412_io_reset),
    .io_out(regs_412_io_out),
    .io_enable(regs_412_io_enable)
  );
  FringeFF regs_413 ( // @[RegFile.scala 66:20:@47503.4]
    .clock(regs_413_clock),
    .reset(regs_413_reset),
    .io_in(regs_413_io_in),
    .io_reset(regs_413_io_reset),
    .io_out(regs_413_io_out),
    .io_enable(regs_413_io_enable)
  );
  FringeFF regs_414 ( // @[RegFile.scala 66:20:@47517.4]
    .clock(regs_414_clock),
    .reset(regs_414_reset),
    .io_in(regs_414_io_in),
    .io_reset(regs_414_io_reset),
    .io_out(regs_414_io_out),
    .io_enable(regs_414_io_enable)
  );
  FringeFF regs_415 ( // @[RegFile.scala 66:20:@47531.4]
    .clock(regs_415_clock),
    .reset(regs_415_reset),
    .io_in(regs_415_io_in),
    .io_reset(regs_415_io_reset),
    .io_out(regs_415_io_out),
    .io_enable(regs_415_io_enable)
  );
  FringeFF regs_416 ( // @[RegFile.scala 66:20:@47545.4]
    .clock(regs_416_clock),
    .reset(regs_416_reset),
    .io_in(regs_416_io_in),
    .io_reset(regs_416_io_reset),
    .io_out(regs_416_io_out),
    .io_enable(regs_416_io_enable)
  );
  FringeFF regs_417 ( // @[RegFile.scala 66:20:@47559.4]
    .clock(regs_417_clock),
    .reset(regs_417_reset),
    .io_in(regs_417_io_in),
    .io_reset(regs_417_io_reset),
    .io_out(regs_417_io_out),
    .io_enable(regs_417_io_enable)
  );
  FringeFF regs_418 ( // @[RegFile.scala 66:20:@47573.4]
    .clock(regs_418_clock),
    .reset(regs_418_reset),
    .io_in(regs_418_io_in),
    .io_reset(regs_418_io_reset),
    .io_out(regs_418_io_out),
    .io_enable(regs_418_io_enable)
  );
  FringeFF regs_419 ( // @[RegFile.scala 66:20:@47587.4]
    .clock(regs_419_clock),
    .reset(regs_419_reset),
    .io_in(regs_419_io_in),
    .io_reset(regs_419_io_reset),
    .io_out(regs_419_io_out),
    .io_enable(regs_419_io_enable)
  );
  FringeFF regs_420 ( // @[RegFile.scala 66:20:@47601.4]
    .clock(regs_420_clock),
    .reset(regs_420_reset),
    .io_in(regs_420_io_in),
    .io_reset(regs_420_io_reset),
    .io_out(regs_420_io_out),
    .io_enable(regs_420_io_enable)
  );
  FringeFF regs_421 ( // @[RegFile.scala 66:20:@47615.4]
    .clock(regs_421_clock),
    .reset(regs_421_reset),
    .io_in(regs_421_io_in),
    .io_reset(regs_421_io_reset),
    .io_out(regs_421_io_out),
    .io_enable(regs_421_io_enable)
  );
  FringeFF regs_422 ( // @[RegFile.scala 66:20:@47629.4]
    .clock(regs_422_clock),
    .reset(regs_422_reset),
    .io_in(regs_422_io_in),
    .io_reset(regs_422_io_reset),
    .io_out(regs_422_io_out),
    .io_enable(regs_422_io_enable)
  );
  FringeFF regs_423 ( // @[RegFile.scala 66:20:@47643.4]
    .clock(regs_423_clock),
    .reset(regs_423_reset),
    .io_in(regs_423_io_in),
    .io_reset(regs_423_io_reset),
    .io_out(regs_423_io_out),
    .io_enable(regs_423_io_enable)
  );
  FringeFF regs_424 ( // @[RegFile.scala 66:20:@47657.4]
    .clock(regs_424_clock),
    .reset(regs_424_reset),
    .io_in(regs_424_io_in),
    .io_reset(regs_424_io_reset),
    .io_out(regs_424_io_out),
    .io_enable(regs_424_io_enable)
  );
  FringeFF regs_425 ( // @[RegFile.scala 66:20:@47671.4]
    .clock(regs_425_clock),
    .reset(regs_425_reset),
    .io_in(regs_425_io_in),
    .io_reset(regs_425_io_reset),
    .io_out(regs_425_io_out),
    .io_enable(regs_425_io_enable)
  );
  FringeFF regs_426 ( // @[RegFile.scala 66:20:@47685.4]
    .clock(regs_426_clock),
    .reset(regs_426_reset),
    .io_in(regs_426_io_in),
    .io_reset(regs_426_io_reset),
    .io_out(regs_426_io_out),
    .io_enable(regs_426_io_enable)
  );
  FringeFF regs_427 ( // @[RegFile.scala 66:20:@47699.4]
    .clock(regs_427_clock),
    .reset(regs_427_reset),
    .io_in(regs_427_io_in),
    .io_reset(regs_427_io_reset),
    .io_out(regs_427_io_out),
    .io_enable(regs_427_io_enable)
  );
  FringeFF regs_428 ( // @[RegFile.scala 66:20:@47713.4]
    .clock(regs_428_clock),
    .reset(regs_428_reset),
    .io_in(regs_428_io_in),
    .io_reset(regs_428_io_reset),
    .io_out(regs_428_io_out),
    .io_enable(regs_428_io_enable)
  );
  FringeFF regs_429 ( // @[RegFile.scala 66:20:@47727.4]
    .clock(regs_429_clock),
    .reset(regs_429_reset),
    .io_in(regs_429_io_in),
    .io_reset(regs_429_io_reset),
    .io_out(regs_429_io_out),
    .io_enable(regs_429_io_enable)
  );
  FringeFF regs_430 ( // @[RegFile.scala 66:20:@47741.4]
    .clock(regs_430_clock),
    .reset(regs_430_reset),
    .io_in(regs_430_io_in),
    .io_reset(regs_430_io_reset),
    .io_out(regs_430_io_out),
    .io_enable(regs_430_io_enable)
  );
  FringeFF regs_431 ( // @[RegFile.scala 66:20:@47755.4]
    .clock(regs_431_clock),
    .reset(regs_431_reset),
    .io_in(regs_431_io_in),
    .io_reset(regs_431_io_reset),
    .io_out(regs_431_io_out),
    .io_enable(regs_431_io_enable)
  );
  FringeFF regs_432 ( // @[RegFile.scala 66:20:@47769.4]
    .clock(regs_432_clock),
    .reset(regs_432_reset),
    .io_in(regs_432_io_in),
    .io_reset(regs_432_io_reset),
    .io_out(regs_432_io_out),
    .io_enable(regs_432_io_enable)
  );
  FringeFF regs_433 ( // @[RegFile.scala 66:20:@47783.4]
    .clock(regs_433_clock),
    .reset(regs_433_reset),
    .io_in(regs_433_io_in),
    .io_reset(regs_433_io_reset),
    .io_out(regs_433_io_out),
    .io_enable(regs_433_io_enable)
  );
  FringeFF regs_434 ( // @[RegFile.scala 66:20:@47797.4]
    .clock(regs_434_clock),
    .reset(regs_434_reset),
    .io_in(regs_434_io_in),
    .io_reset(regs_434_io_reset),
    .io_out(regs_434_io_out),
    .io_enable(regs_434_io_enable)
  );
  FringeFF regs_435 ( // @[RegFile.scala 66:20:@47811.4]
    .clock(regs_435_clock),
    .reset(regs_435_reset),
    .io_in(regs_435_io_in),
    .io_reset(regs_435_io_reset),
    .io_out(regs_435_io_out),
    .io_enable(regs_435_io_enable)
  );
  FringeFF regs_436 ( // @[RegFile.scala 66:20:@47825.4]
    .clock(regs_436_clock),
    .reset(regs_436_reset),
    .io_in(regs_436_io_in),
    .io_reset(regs_436_io_reset),
    .io_out(regs_436_io_out),
    .io_enable(regs_436_io_enable)
  );
  FringeFF regs_437 ( // @[RegFile.scala 66:20:@47839.4]
    .clock(regs_437_clock),
    .reset(regs_437_reset),
    .io_in(regs_437_io_in),
    .io_reset(regs_437_io_reset),
    .io_out(regs_437_io_out),
    .io_enable(regs_437_io_enable)
  );
  FringeFF regs_438 ( // @[RegFile.scala 66:20:@47853.4]
    .clock(regs_438_clock),
    .reset(regs_438_reset),
    .io_in(regs_438_io_in),
    .io_reset(regs_438_io_reset),
    .io_out(regs_438_io_out),
    .io_enable(regs_438_io_enable)
  );
  FringeFF regs_439 ( // @[RegFile.scala 66:20:@47867.4]
    .clock(regs_439_clock),
    .reset(regs_439_reset),
    .io_in(regs_439_io_in),
    .io_reset(regs_439_io_reset),
    .io_out(regs_439_io_out),
    .io_enable(regs_439_io_enable)
  );
  FringeFF regs_440 ( // @[RegFile.scala 66:20:@47881.4]
    .clock(regs_440_clock),
    .reset(regs_440_reset),
    .io_in(regs_440_io_in),
    .io_reset(regs_440_io_reset),
    .io_out(regs_440_io_out),
    .io_enable(regs_440_io_enable)
  );
  FringeFF regs_441 ( // @[RegFile.scala 66:20:@47895.4]
    .clock(regs_441_clock),
    .reset(regs_441_reset),
    .io_in(regs_441_io_in),
    .io_reset(regs_441_io_reset),
    .io_out(regs_441_io_out),
    .io_enable(regs_441_io_enable)
  );
  FringeFF regs_442 ( // @[RegFile.scala 66:20:@47909.4]
    .clock(regs_442_clock),
    .reset(regs_442_reset),
    .io_in(regs_442_io_in),
    .io_reset(regs_442_io_reset),
    .io_out(regs_442_io_out),
    .io_enable(regs_442_io_enable)
  );
  FringeFF regs_443 ( // @[RegFile.scala 66:20:@47923.4]
    .clock(regs_443_clock),
    .reset(regs_443_reset),
    .io_in(regs_443_io_in),
    .io_reset(regs_443_io_reset),
    .io_out(regs_443_io_out),
    .io_enable(regs_443_io_enable)
  );
  FringeFF regs_444 ( // @[RegFile.scala 66:20:@47937.4]
    .clock(regs_444_clock),
    .reset(regs_444_reset),
    .io_in(regs_444_io_in),
    .io_reset(regs_444_io_reset),
    .io_out(regs_444_io_out),
    .io_enable(regs_444_io_enable)
  );
  FringeFF regs_445 ( // @[RegFile.scala 66:20:@47951.4]
    .clock(regs_445_clock),
    .reset(regs_445_reset),
    .io_in(regs_445_io_in),
    .io_reset(regs_445_io_reset),
    .io_out(regs_445_io_out),
    .io_enable(regs_445_io_enable)
  );
  FringeFF regs_446 ( // @[RegFile.scala 66:20:@47965.4]
    .clock(regs_446_clock),
    .reset(regs_446_reset),
    .io_in(regs_446_io_in),
    .io_reset(regs_446_io_reset),
    .io_out(regs_446_io_out),
    .io_enable(regs_446_io_enable)
  );
  FringeFF regs_447 ( // @[RegFile.scala 66:20:@47979.4]
    .clock(regs_447_clock),
    .reset(regs_447_reset),
    .io_in(regs_447_io_in),
    .io_reset(regs_447_io_reset),
    .io_out(regs_447_io_out),
    .io_enable(regs_447_io_enable)
  );
  FringeFF regs_448 ( // @[RegFile.scala 66:20:@47993.4]
    .clock(regs_448_clock),
    .reset(regs_448_reset),
    .io_in(regs_448_io_in),
    .io_reset(regs_448_io_reset),
    .io_out(regs_448_io_out),
    .io_enable(regs_448_io_enable)
  );
  FringeFF regs_449 ( // @[RegFile.scala 66:20:@48007.4]
    .clock(regs_449_clock),
    .reset(regs_449_reset),
    .io_in(regs_449_io_in),
    .io_reset(regs_449_io_reset),
    .io_out(regs_449_io_out),
    .io_enable(regs_449_io_enable)
  );
  FringeFF regs_450 ( // @[RegFile.scala 66:20:@48021.4]
    .clock(regs_450_clock),
    .reset(regs_450_reset),
    .io_in(regs_450_io_in),
    .io_reset(regs_450_io_reset),
    .io_out(regs_450_io_out),
    .io_enable(regs_450_io_enable)
  );
  FringeFF regs_451 ( // @[RegFile.scala 66:20:@48035.4]
    .clock(regs_451_clock),
    .reset(regs_451_reset),
    .io_in(regs_451_io_in),
    .io_reset(regs_451_io_reset),
    .io_out(regs_451_io_out),
    .io_enable(regs_451_io_enable)
  );
  FringeFF regs_452 ( // @[RegFile.scala 66:20:@48049.4]
    .clock(regs_452_clock),
    .reset(regs_452_reset),
    .io_in(regs_452_io_in),
    .io_reset(regs_452_io_reset),
    .io_out(regs_452_io_out),
    .io_enable(regs_452_io_enable)
  );
  FringeFF regs_453 ( // @[RegFile.scala 66:20:@48063.4]
    .clock(regs_453_clock),
    .reset(regs_453_reset),
    .io_in(regs_453_io_in),
    .io_reset(regs_453_io_reset),
    .io_out(regs_453_io_out),
    .io_enable(regs_453_io_enable)
  );
  FringeFF regs_454 ( // @[RegFile.scala 66:20:@48077.4]
    .clock(regs_454_clock),
    .reset(regs_454_reset),
    .io_in(regs_454_io_in),
    .io_reset(regs_454_io_reset),
    .io_out(regs_454_io_out),
    .io_enable(regs_454_io_enable)
  );
  FringeFF regs_455 ( // @[RegFile.scala 66:20:@48091.4]
    .clock(regs_455_clock),
    .reset(regs_455_reset),
    .io_in(regs_455_io_in),
    .io_reset(regs_455_io_reset),
    .io_out(regs_455_io_out),
    .io_enable(regs_455_io_enable)
  );
  FringeFF regs_456 ( // @[RegFile.scala 66:20:@48105.4]
    .clock(regs_456_clock),
    .reset(regs_456_reset),
    .io_in(regs_456_io_in),
    .io_reset(regs_456_io_reset),
    .io_out(regs_456_io_out),
    .io_enable(regs_456_io_enable)
  );
  FringeFF regs_457 ( // @[RegFile.scala 66:20:@48119.4]
    .clock(regs_457_clock),
    .reset(regs_457_reset),
    .io_in(regs_457_io_in),
    .io_reset(regs_457_io_reset),
    .io_out(regs_457_io_out),
    .io_enable(regs_457_io_enable)
  );
  FringeFF regs_458 ( // @[RegFile.scala 66:20:@48133.4]
    .clock(regs_458_clock),
    .reset(regs_458_reset),
    .io_in(regs_458_io_in),
    .io_reset(regs_458_io_reset),
    .io_out(regs_458_io_out),
    .io_enable(regs_458_io_enable)
  );
  FringeFF regs_459 ( // @[RegFile.scala 66:20:@48147.4]
    .clock(regs_459_clock),
    .reset(regs_459_reset),
    .io_in(regs_459_io_in),
    .io_reset(regs_459_io_reset),
    .io_out(regs_459_io_out),
    .io_enable(regs_459_io_enable)
  );
  FringeFF regs_460 ( // @[RegFile.scala 66:20:@48161.4]
    .clock(regs_460_clock),
    .reset(regs_460_reset),
    .io_in(regs_460_io_in),
    .io_reset(regs_460_io_reset),
    .io_out(regs_460_io_out),
    .io_enable(regs_460_io_enable)
  );
  FringeFF regs_461 ( // @[RegFile.scala 66:20:@48175.4]
    .clock(regs_461_clock),
    .reset(regs_461_reset),
    .io_in(regs_461_io_in),
    .io_reset(regs_461_io_reset),
    .io_out(regs_461_io_out),
    .io_enable(regs_461_io_enable)
  );
  FringeFF regs_462 ( // @[RegFile.scala 66:20:@48189.4]
    .clock(regs_462_clock),
    .reset(regs_462_reset),
    .io_in(regs_462_io_in),
    .io_reset(regs_462_io_reset),
    .io_out(regs_462_io_out),
    .io_enable(regs_462_io_enable)
  );
  FringeFF regs_463 ( // @[RegFile.scala 66:20:@48203.4]
    .clock(regs_463_clock),
    .reset(regs_463_reset),
    .io_in(regs_463_io_in),
    .io_reset(regs_463_io_reset),
    .io_out(regs_463_io_out),
    .io_enable(regs_463_io_enable)
  );
  FringeFF regs_464 ( // @[RegFile.scala 66:20:@48217.4]
    .clock(regs_464_clock),
    .reset(regs_464_reset),
    .io_in(regs_464_io_in),
    .io_reset(regs_464_io_reset),
    .io_out(regs_464_io_out),
    .io_enable(regs_464_io_enable)
  );
  FringeFF regs_465 ( // @[RegFile.scala 66:20:@48231.4]
    .clock(regs_465_clock),
    .reset(regs_465_reset),
    .io_in(regs_465_io_in),
    .io_reset(regs_465_io_reset),
    .io_out(regs_465_io_out),
    .io_enable(regs_465_io_enable)
  );
  FringeFF regs_466 ( // @[RegFile.scala 66:20:@48245.4]
    .clock(regs_466_clock),
    .reset(regs_466_reset),
    .io_in(regs_466_io_in),
    .io_reset(regs_466_io_reset),
    .io_out(regs_466_io_out),
    .io_enable(regs_466_io_enable)
  );
  FringeFF regs_467 ( // @[RegFile.scala 66:20:@48259.4]
    .clock(regs_467_clock),
    .reset(regs_467_reset),
    .io_in(regs_467_io_in),
    .io_reset(regs_467_io_reset),
    .io_out(regs_467_io_out),
    .io_enable(regs_467_io_enable)
  );
  FringeFF regs_468 ( // @[RegFile.scala 66:20:@48273.4]
    .clock(regs_468_clock),
    .reset(regs_468_reset),
    .io_in(regs_468_io_in),
    .io_reset(regs_468_io_reset),
    .io_out(regs_468_io_out),
    .io_enable(regs_468_io_enable)
  );
  FringeFF regs_469 ( // @[RegFile.scala 66:20:@48287.4]
    .clock(regs_469_clock),
    .reset(regs_469_reset),
    .io_in(regs_469_io_in),
    .io_reset(regs_469_io_reset),
    .io_out(regs_469_io_out),
    .io_enable(regs_469_io_enable)
  );
  FringeFF regs_470 ( // @[RegFile.scala 66:20:@48301.4]
    .clock(regs_470_clock),
    .reset(regs_470_reset),
    .io_in(regs_470_io_in),
    .io_reset(regs_470_io_reset),
    .io_out(regs_470_io_out),
    .io_enable(regs_470_io_enable)
  );
  FringeFF regs_471 ( // @[RegFile.scala 66:20:@48315.4]
    .clock(regs_471_clock),
    .reset(regs_471_reset),
    .io_in(regs_471_io_in),
    .io_reset(regs_471_io_reset),
    .io_out(regs_471_io_out),
    .io_enable(regs_471_io_enable)
  );
  FringeFF regs_472 ( // @[RegFile.scala 66:20:@48329.4]
    .clock(regs_472_clock),
    .reset(regs_472_reset),
    .io_in(regs_472_io_in),
    .io_reset(regs_472_io_reset),
    .io_out(regs_472_io_out),
    .io_enable(regs_472_io_enable)
  );
  FringeFF regs_473 ( // @[RegFile.scala 66:20:@48343.4]
    .clock(regs_473_clock),
    .reset(regs_473_reset),
    .io_in(regs_473_io_in),
    .io_reset(regs_473_io_reset),
    .io_out(regs_473_io_out),
    .io_enable(regs_473_io_enable)
  );
  FringeFF regs_474 ( // @[RegFile.scala 66:20:@48357.4]
    .clock(regs_474_clock),
    .reset(regs_474_reset),
    .io_in(regs_474_io_in),
    .io_reset(regs_474_io_reset),
    .io_out(regs_474_io_out),
    .io_enable(regs_474_io_enable)
  );
  FringeFF regs_475 ( // @[RegFile.scala 66:20:@48371.4]
    .clock(regs_475_clock),
    .reset(regs_475_reset),
    .io_in(regs_475_io_in),
    .io_reset(regs_475_io_reset),
    .io_out(regs_475_io_out),
    .io_enable(regs_475_io_enable)
  );
  FringeFF regs_476 ( // @[RegFile.scala 66:20:@48385.4]
    .clock(regs_476_clock),
    .reset(regs_476_reset),
    .io_in(regs_476_io_in),
    .io_reset(regs_476_io_reset),
    .io_out(regs_476_io_out),
    .io_enable(regs_476_io_enable)
  );
  FringeFF regs_477 ( // @[RegFile.scala 66:20:@48399.4]
    .clock(regs_477_clock),
    .reset(regs_477_reset),
    .io_in(regs_477_io_in),
    .io_reset(regs_477_io_reset),
    .io_out(regs_477_io_out),
    .io_enable(regs_477_io_enable)
  );
  FringeFF regs_478 ( // @[RegFile.scala 66:20:@48413.4]
    .clock(regs_478_clock),
    .reset(regs_478_reset),
    .io_in(regs_478_io_in),
    .io_reset(regs_478_io_reset),
    .io_out(regs_478_io_out),
    .io_enable(regs_478_io_enable)
  );
  FringeFF regs_479 ( // @[RegFile.scala 66:20:@48427.4]
    .clock(regs_479_clock),
    .reset(regs_479_reset),
    .io_in(regs_479_io_in),
    .io_reset(regs_479_io_reset),
    .io_out(regs_479_io_out),
    .io_enable(regs_479_io_enable)
  );
  FringeFF regs_480 ( // @[RegFile.scala 66:20:@48441.4]
    .clock(regs_480_clock),
    .reset(regs_480_reset),
    .io_in(regs_480_io_in),
    .io_reset(regs_480_io_reset),
    .io_out(regs_480_io_out),
    .io_enable(regs_480_io_enable)
  );
  FringeFF regs_481 ( // @[RegFile.scala 66:20:@48455.4]
    .clock(regs_481_clock),
    .reset(regs_481_reset),
    .io_in(regs_481_io_in),
    .io_reset(regs_481_io_reset),
    .io_out(regs_481_io_out),
    .io_enable(regs_481_io_enable)
  );
  FringeFF regs_482 ( // @[RegFile.scala 66:20:@48469.4]
    .clock(regs_482_clock),
    .reset(regs_482_reset),
    .io_in(regs_482_io_in),
    .io_reset(regs_482_io_reset),
    .io_out(regs_482_io_out),
    .io_enable(regs_482_io_enable)
  );
  FringeFF regs_483 ( // @[RegFile.scala 66:20:@48483.4]
    .clock(regs_483_clock),
    .reset(regs_483_reset),
    .io_in(regs_483_io_in),
    .io_reset(regs_483_io_reset),
    .io_out(regs_483_io_out),
    .io_enable(regs_483_io_enable)
  );
  FringeFF regs_484 ( // @[RegFile.scala 66:20:@48497.4]
    .clock(regs_484_clock),
    .reset(regs_484_reset),
    .io_in(regs_484_io_in),
    .io_reset(regs_484_io_reset),
    .io_out(regs_484_io_out),
    .io_enable(regs_484_io_enable)
  );
  FringeFF regs_485 ( // @[RegFile.scala 66:20:@48511.4]
    .clock(regs_485_clock),
    .reset(regs_485_reset),
    .io_in(regs_485_io_in),
    .io_reset(regs_485_io_reset),
    .io_out(regs_485_io_out),
    .io_enable(regs_485_io_enable)
  );
  FringeFF regs_486 ( // @[RegFile.scala 66:20:@48525.4]
    .clock(regs_486_clock),
    .reset(regs_486_reset),
    .io_in(regs_486_io_in),
    .io_reset(regs_486_io_reset),
    .io_out(regs_486_io_out),
    .io_enable(regs_486_io_enable)
  );
  FringeFF regs_487 ( // @[RegFile.scala 66:20:@48539.4]
    .clock(regs_487_clock),
    .reset(regs_487_reset),
    .io_in(regs_487_io_in),
    .io_reset(regs_487_io_reset),
    .io_out(regs_487_io_out),
    .io_enable(regs_487_io_enable)
  );
  FringeFF regs_488 ( // @[RegFile.scala 66:20:@48553.4]
    .clock(regs_488_clock),
    .reset(regs_488_reset),
    .io_in(regs_488_io_in),
    .io_reset(regs_488_io_reset),
    .io_out(regs_488_io_out),
    .io_enable(regs_488_io_enable)
  );
  FringeFF regs_489 ( // @[RegFile.scala 66:20:@48567.4]
    .clock(regs_489_clock),
    .reset(regs_489_reset),
    .io_in(regs_489_io_in),
    .io_reset(regs_489_io_reset),
    .io_out(regs_489_io_out),
    .io_enable(regs_489_io_enable)
  );
  FringeFF regs_490 ( // @[RegFile.scala 66:20:@48581.4]
    .clock(regs_490_clock),
    .reset(regs_490_reset),
    .io_in(regs_490_io_in),
    .io_reset(regs_490_io_reset),
    .io_out(regs_490_io_out),
    .io_enable(regs_490_io_enable)
  );
  FringeFF regs_491 ( // @[RegFile.scala 66:20:@48595.4]
    .clock(regs_491_clock),
    .reset(regs_491_reset),
    .io_in(regs_491_io_in),
    .io_reset(regs_491_io_reset),
    .io_out(regs_491_io_out),
    .io_enable(regs_491_io_enable)
  );
  FringeFF regs_492 ( // @[RegFile.scala 66:20:@48609.4]
    .clock(regs_492_clock),
    .reset(regs_492_reset),
    .io_in(regs_492_io_in),
    .io_reset(regs_492_io_reset),
    .io_out(regs_492_io_out),
    .io_enable(regs_492_io_enable)
  );
  FringeFF regs_493 ( // @[RegFile.scala 66:20:@48623.4]
    .clock(regs_493_clock),
    .reset(regs_493_reset),
    .io_in(regs_493_io_in),
    .io_reset(regs_493_io_reset),
    .io_out(regs_493_io_out),
    .io_enable(regs_493_io_enable)
  );
  FringeFF regs_494 ( // @[RegFile.scala 66:20:@48637.4]
    .clock(regs_494_clock),
    .reset(regs_494_reset),
    .io_in(regs_494_io_in),
    .io_reset(regs_494_io_reset),
    .io_out(regs_494_io_out),
    .io_enable(regs_494_io_enable)
  );
  FringeFF regs_495 ( // @[RegFile.scala 66:20:@48651.4]
    .clock(regs_495_clock),
    .reset(regs_495_reset),
    .io_in(regs_495_io_in),
    .io_reset(regs_495_io_reset),
    .io_out(regs_495_io_out),
    .io_enable(regs_495_io_enable)
  );
  FringeFF regs_496 ( // @[RegFile.scala 66:20:@48665.4]
    .clock(regs_496_clock),
    .reset(regs_496_reset),
    .io_in(regs_496_io_in),
    .io_reset(regs_496_io_reset),
    .io_out(regs_496_io_out),
    .io_enable(regs_496_io_enable)
  );
  FringeFF regs_497 ( // @[RegFile.scala 66:20:@48679.4]
    .clock(regs_497_clock),
    .reset(regs_497_reset),
    .io_in(regs_497_io_in),
    .io_reset(regs_497_io_reset),
    .io_out(regs_497_io_out),
    .io_enable(regs_497_io_enable)
  );
  FringeFF regs_498 ( // @[RegFile.scala 66:20:@48693.4]
    .clock(regs_498_clock),
    .reset(regs_498_reset),
    .io_in(regs_498_io_in),
    .io_reset(regs_498_io_reset),
    .io_out(regs_498_io_out),
    .io_enable(regs_498_io_enable)
  );
  FringeFF regs_499 ( // @[RegFile.scala 66:20:@48707.4]
    .clock(regs_499_clock),
    .reset(regs_499_reset),
    .io_in(regs_499_io_in),
    .io_reset(regs_499_io_reset),
    .io_out(regs_499_io_out),
    .io_enable(regs_499_io_enable)
  );
  FringeFF regs_500 ( // @[RegFile.scala 66:20:@48721.4]
    .clock(regs_500_clock),
    .reset(regs_500_reset),
    .io_in(regs_500_io_in),
    .io_reset(regs_500_io_reset),
    .io_out(regs_500_io_out),
    .io_enable(regs_500_io_enable)
  );
  FringeFF regs_501 ( // @[RegFile.scala 66:20:@48735.4]
    .clock(regs_501_clock),
    .reset(regs_501_reset),
    .io_in(regs_501_io_in),
    .io_reset(regs_501_io_reset),
    .io_out(regs_501_io_out),
    .io_enable(regs_501_io_enable)
  );
  FringeFF regs_502 ( // @[RegFile.scala 66:20:@48749.4]
    .clock(regs_502_clock),
    .reset(regs_502_reset),
    .io_in(regs_502_io_in),
    .io_reset(regs_502_io_reset),
    .io_out(regs_502_io_out),
    .io_enable(regs_502_io_enable)
  );
  FringeFF regs_503 ( // @[RegFile.scala 66:20:@48763.4]
    .clock(regs_503_clock),
    .reset(regs_503_reset),
    .io_in(regs_503_io_in),
    .io_reset(regs_503_io_reset),
    .io_out(regs_503_io_out),
    .io_enable(regs_503_io_enable)
  );
  FringeFF regs_504 ( // @[RegFile.scala 66:20:@48777.4]
    .clock(regs_504_clock),
    .reset(regs_504_reset),
    .io_in(regs_504_io_in),
    .io_reset(regs_504_io_reset),
    .io_out(regs_504_io_out),
    .io_enable(regs_504_io_enable)
  );
  FringeFF regs_505 ( // @[RegFile.scala 66:20:@48791.4]
    .clock(regs_505_clock),
    .reset(regs_505_reset),
    .io_in(regs_505_io_in),
    .io_reset(regs_505_io_reset),
    .io_out(regs_505_io_out),
    .io_enable(regs_505_io_enable)
  );
  FringeFF regs_506 ( // @[RegFile.scala 66:20:@48805.4]
    .clock(regs_506_clock),
    .reset(regs_506_reset),
    .io_in(regs_506_io_in),
    .io_reset(regs_506_io_reset),
    .io_out(regs_506_io_out),
    .io_enable(regs_506_io_enable)
  );
  FringeFF regs_507 ( // @[RegFile.scala 66:20:@48819.4]
    .clock(regs_507_clock),
    .reset(regs_507_reset),
    .io_in(regs_507_io_in),
    .io_reset(regs_507_io_reset),
    .io_out(regs_507_io_out),
    .io_enable(regs_507_io_enable)
  );
  FringeFF regs_508 ( // @[RegFile.scala 66:20:@48833.4]
    .clock(regs_508_clock),
    .reset(regs_508_reset),
    .io_in(regs_508_io_in),
    .io_reset(regs_508_io_reset),
    .io_out(regs_508_io_out),
    .io_enable(regs_508_io_enable)
  );
  FringeFF regs_509 ( // @[RegFile.scala 66:20:@48847.4]
    .clock(regs_509_clock),
    .reset(regs_509_reset),
    .io_in(regs_509_io_in),
    .io_reset(regs_509_io_reset),
    .io_out(regs_509_io_out),
    .io_enable(regs_509_io_enable)
  );
  FringeFF regs_510 ( // @[RegFile.scala 66:20:@48861.4]
    .clock(regs_510_clock),
    .reset(regs_510_reset),
    .io_in(regs_510_io_in),
    .io_reset(regs_510_io_reset),
    .io_out(regs_510_io_out),
    .io_enable(regs_510_io_enable)
  );
  FringeFF regs_511 ( // @[RegFile.scala 66:20:@48875.4]
    .clock(regs_511_clock),
    .reset(regs_511_reset),
    .io_in(regs_511_io_in),
    .io_reset(regs_511_io_reset),
    .io_out(regs_511_io_out),
    .io_enable(regs_511_io_enable)
  );
  FringeFF regs_512 ( // @[RegFile.scala 66:20:@48889.4]
    .clock(regs_512_clock),
    .reset(regs_512_reset),
    .io_in(regs_512_io_in),
    .io_reset(regs_512_io_reset),
    .io_out(regs_512_io_out),
    .io_enable(regs_512_io_enable)
  );
  FringeFF regs_513 ( // @[RegFile.scala 66:20:@48903.4]
    .clock(regs_513_clock),
    .reset(regs_513_reset),
    .io_in(regs_513_io_in),
    .io_reset(regs_513_io_reset),
    .io_out(regs_513_io_out),
    .io_enable(regs_513_io_enable)
  );
  FringeFF regs_514 ( // @[RegFile.scala 66:20:@48917.4]
    .clock(regs_514_clock),
    .reset(regs_514_reset),
    .io_in(regs_514_io_in),
    .io_reset(regs_514_io_reset),
    .io_out(regs_514_io_out),
    .io_enable(regs_514_io_enable)
  );
  FringeFF regs_515 ( // @[RegFile.scala 66:20:@48931.4]
    .clock(regs_515_clock),
    .reset(regs_515_reset),
    .io_in(regs_515_io_in),
    .io_reset(regs_515_io_reset),
    .io_out(regs_515_io_out),
    .io_enable(regs_515_io_enable)
  );
  FringeFF regs_516 ( // @[RegFile.scala 66:20:@48945.4]
    .clock(regs_516_clock),
    .reset(regs_516_reset),
    .io_in(regs_516_io_in),
    .io_reset(regs_516_io_reset),
    .io_out(regs_516_io_out),
    .io_enable(regs_516_io_enable)
  );
  FringeFF regs_517 ( // @[RegFile.scala 66:20:@48959.4]
    .clock(regs_517_clock),
    .reset(regs_517_reset),
    .io_in(regs_517_io_in),
    .io_reset(regs_517_io_reset),
    .io_out(regs_517_io_out),
    .io_enable(regs_517_io_enable)
  );
  FringeFF regs_518 ( // @[RegFile.scala 66:20:@48973.4]
    .clock(regs_518_clock),
    .reset(regs_518_reset),
    .io_in(regs_518_io_in),
    .io_reset(regs_518_io_reset),
    .io_out(regs_518_io_out),
    .io_enable(regs_518_io_enable)
  );
  FringeFF regs_519 ( // @[RegFile.scala 66:20:@48987.4]
    .clock(regs_519_clock),
    .reset(regs_519_reset),
    .io_in(regs_519_io_in),
    .io_reset(regs_519_io_reset),
    .io_out(regs_519_io_out),
    .io_enable(regs_519_io_enable)
  );
  FringeFF regs_520 ( // @[RegFile.scala 66:20:@49001.4]
    .clock(regs_520_clock),
    .reset(regs_520_reset),
    .io_in(regs_520_io_in),
    .io_reset(regs_520_io_reset),
    .io_out(regs_520_io_out),
    .io_enable(regs_520_io_enable)
  );
  FringeFF regs_521 ( // @[RegFile.scala 66:20:@49015.4]
    .clock(regs_521_clock),
    .reset(regs_521_reset),
    .io_in(regs_521_io_in),
    .io_reset(regs_521_io_reset),
    .io_out(regs_521_io_out),
    .io_enable(regs_521_io_enable)
  );
  FringeFF regs_522 ( // @[RegFile.scala 66:20:@49029.4]
    .clock(regs_522_clock),
    .reset(regs_522_reset),
    .io_in(regs_522_io_in),
    .io_reset(regs_522_io_reset),
    .io_out(regs_522_io_out),
    .io_enable(regs_522_io_enable)
  );
  FringeFF regs_523 ( // @[RegFile.scala 66:20:@49043.4]
    .clock(regs_523_clock),
    .reset(regs_523_reset),
    .io_in(regs_523_io_in),
    .io_reset(regs_523_io_reset),
    .io_out(regs_523_io_out),
    .io_enable(regs_523_io_enable)
  );
  FringeFF regs_524 ( // @[RegFile.scala 66:20:@49057.4]
    .clock(regs_524_clock),
    .reset(regs_524_reset),
    .io_in(regs_524_io_in),
    .io_reset(regs_524_io_reset),
    .io_out(regs_524_io_out),
    .io_enable(regs_524_io_enable)
  );
  FringeFF regs_525 ( // @[RegFile.scala 66:20:@49071.4]
    .clock(regs_525_clock),
    .reset(regs_525_reset),
    .io_in(regs_525_io_in),
    .io_reset(regs_525_io_reset),
    .io_out(regs_525_io_out),
    .io_enable(regs_525_io_enable)
  );
  FringeFF regs_526 ( // @[RegFile.scala 66:20:@49085.4]
    .clock(regs_526_clock),
    .reset(regs_526_reset),
    .io_in(regs_526_io_in),
    .io_reset(regs_526_io_reset),
    .io_out(regs_526_io_out),
    .io_enable(regs_526_io_enable)
  );
  FringeFF regs_527 ( // @[RegFile.scala 66:20:@49099.4]
    .clock(regs_527_clock),
    .reset(regs_527_reset),
    .io_in(regs_527_io_in),
    .io_reset(regs_527_io_reset),
    .io_out(regs_527_io_out),
    .io_enable(regs_527_io_enable)
  );
  FringeFF regs_528 ( // @[RegFile.scala 66:20:@49113.4]
    .clock(regs_528_clock),
    .reset(regs_528_reset),
    .io_in(regs_528_io_in),
    .io_reset(regs_528_io_reset),
    .io_out(regs_528_io_out),
    .io_enable(regs_528_io_enable)
  );
  FringeFF regs_529 ( // @[RegFile.scala 66:20:@49127.4]
    .clock(regs_529_clock),
    .reset(regs_529_reset),
    .io_in(regs_529_io_in),
    .io_reset(regs_529_io_reset),
    .io_out(regs_529_io_out),
    .io_enable(regs_529_io_enable)
  );
  FringeFF regs_530 ( // @[RegFile.scala 66:20:@49141.4]
    .clock(regs_530_clock),
    .reset(regs_530_reset),
    .io_in(regs_530_io_in),
    .io_reset(regs_530_io_reset),
    .io_out(regs_530_io_out),
    .io_enable(regs_530_io_enable)
  );
  FringeFF regs_531 ( // @[RegFile.scala 66:20:@49155.4]
    .clock(regs_531_clock),
    .reset(regs_531_reset),
    .io_in(regs_531_io_in),
    .io_reset(regs_531_io_reset),
    .io_out(regs_531_io_out),
    .io_enable(regs_531_io_enable)
  );
  FringeFF regs_532 ( // @[RegFile.scala 66:20:@49169.4]
    .clock(regs_532_clock),
    .reset(regs_532_reset),
    .io_in(regs_532_io_in),
    .io_reset(regs_532_io_reset),
    .io_out(regs_532_io_out),
    .io_enable(regs_532_io_enable)
  );
  FringeFF regs_533 ( // @[RegFile.scala 66:20:@49183.4]
    .clock(regs_533_clock),
    .reset(regs_533_reset),
    .io_in(regs_533_io_in),
    .io_reset(regs_533_io_reset),
    .io_out(regs_533_io_out),
    .io_enable(regs_533_io_enable)
  );
  MuxN rport ( // @[RegFile.scala 95:21:@49197.4]
    .io_ins_0(rport_io_ins_0),
    .io_ins_1(rport_io_ins_1),
    .io_ins_2(rport_io_ins_2),
    .io_ins_3(rport_io_ins_3),
    .io_ins_4(rport_io_ins_4),
    .io_ins_5(rport_io_ins_5),
    .io_ins_6(rport_io_ins_6),
    .io_ins_7(rport_io_ins_7),
    .io_ins_8(rport_io_ins_8),
    .io_ins_9(rport_io_ins_9),
    .io_ins_10(rport_io_ins_10),
    .io_ins_11(rport_io_ins_11),
    .io_ins_12(rport_io_ins_12),
    .io_ins_13(rport_io_ins_13),
    .io_ins_14(rport_io_ins_14),
    .io_ins_15(rport_io_ins_15),
    .io_ins_16(rport_io_ins_16),
    .io_ins_17(rport_io_ins_17),
    .io_ins_18(rport_io_ins_18),
    .io_ins_19(rport_io_ins_19),
    .io_ins_20(rport_io_ins_20),
    .io_ins_21(rport_io_ins_21),
    .io_ins_22(rport_io_ins_22),
    .io_ins_23(rport_io_ins_23),
    .io_ins_24(rport_io_ins_24),
    .io_ins_25(rport_io_ins_25),
    .io_ins_26(rport_io_ins_26),
    .io_ins_27(rport_io_ins_27),
    .io_ins_28(rport_io_ins_28),
    .io_ins_29(rport_io_ins_29),
    .io_ins_30(rport_io_ins_30),
    .io_ins_31(rport_io_ins_31),
    .io_ins_32(rport_io_ins_32),
    .io_ins_33(rport_io_ins_33),
    .io_ins_34(rport_io_ins_34),
    .io_ins_35(rport_io_ins_35),
    .io_ins_36(rport_io_ins_36),
    .io_ins_37(rport_io_ins_37),
    .io_ins_38(rport_io_ins_38),
    .io_ins_39(rport_io_ins_39),
    .io_ins_40(rport_io_ins_40),
    .io_ins_41(rport_io_ins_41),
    .io_ins_42(rport_io_ins_42),
    .io_ins_43(rport_io_ins_43),
    .io_ins_44(rport_io_ins_44),
    .io_ins_45(rport_io_ins_45),
    .io_ins_46(rport_io_ins_46),
    .io_ins_47(rport_io_ins_47),
    .io_ins_48(rport_io_ins_48),
    .io_ins_49(rport_io_ins_49),
    .io_ins_50(rport_io_ins_50),
    .io_ins_51(rport_io_ins_51),
    .io_ins_52(rport_io_ins_52),
    .io_ins_53(rport_io_ins_53),
    .io_ins_54(rport_io_ins_54),
    .io_ins_55(rport_io_ins_55),
    .io_ins_56(rport_io_ins_56),
    .io_ins_57(rport_io_ins_57),
    .io_ins_58(rport_io_ins_58),
    .io_ins_59(rport_io_ins_59),
    .io_ins_60(rport_io_ins_60),
    .io_ins_61(rport_io_ins_61),
    .io_ins_62(rport_io_ins_62),
    .io_ins_63(rport_io_ins_63),
    .io_ins_64(rport_io_ins_64),
    .io_ins_65(rport_io_ins_65),
    .io_ins_66(rport_io_ins_66),
    .io_ins_67(rport_io_ins_67),
    .io_ins_68(rport_io_ins_68),
    .io_ins_69(rport_io_ins_69),
    .io_ins_70(rport_io_ins_70),
    .io_ins_71(rport_io_ins_71),
    .io_ins_72(rport_io_ins_72),
    .io_ins_73(rport_io_ins_73),
    .io_ins_74(rport_io_ins_74),
    .io_ins_75(rport_io_ins_75),
    .io_ins_76(rport_io_ins_76),
    .io_ins_77(rport_io_ins_77),
    .io_ins_78(rport_io_ins_78),
    .io_ins_79(rport_io_ins_79),
    .io_ins_80(rport_io_ins_80),
    .io_ins_81(rport_io_ins_81),
    .io_ins_82(rport_io_ins_82),
    .io_ins_83(rport_io_ins_83),
    .io_ins_84(rport_io_ins_84),
    .io_ins_85(rport_io_ins_85),
    .io_ins_86(rport_io_ins_86),
    .io_ins_87(rport_io_ins_87),
    .io_ins_88(rport_io_ins_88),
    .io_ins_89(rport_io_ins_89),
    .io_ins_90(rport_io_ins_90),
    .io_ins_91(rport_io_ins_91),
    .io_ins_92(rport_io_ins_92),
    .io_ins_93(rport_io_ins_93),
    .io_ins_94(rport_io_ins_94),
    .io_ins_95(rport_io_ins_95),
    .io_ins_96(rport_io_ins_96),
    .io_ins_97(rport_io_ins_97),
    .io_ins_98(rport_io_ins_98),
    .io_ins_99(rport_io_ins_99),
    .io_ins_100(rport_io_ins_100),
    .io_ins_101(rport_io_ins_101),
    .io_ins_102(rport_io_ins_102),
    .io_ins_103(rport_io_ins_103),
    .io_ins_104(rport_io_ins_104),
    .io_ins_105(rport_io_ins_105),
    .io_ins_106(rport_io_ins_106),
    .io_ins_107(rport_io_ins_107),
    .io_ins_108(rport_io_ins_108),
    .io_ins_109(rport_io_ins_109),
    .io_ins_110(rport_io_ins_110),
    .io_ins_111(rport_io_ins_111),
    .io_ins_112(rport_io_ins_112),
    .io_ins_113(rport_io_ins_113),
    .io_ins_114(rport_io_ins_114),
    .io_ins_115(rport_io_ins_115),
    .io_ins_116(rport_io_ins_116),
    .io_ins_117(rport_io_ins_117),
    .io_ins_118(rport_io_ins_118),
    .io_ins_119(rport_io_ins_119),
    .io_ins_120(rport_io_ins_120),
    .io_ins_121(rport_io_ins_121),
    .io_ins_122(rport_io_ins_122),
    .io_ins_123(rport_io_ins_123),
    .io_ins_124(rport_io_ins_124),
    .io_ins_125(rport_io_ins_125),
    .io_ins_126(rport_io_ins_126),
    .io_ins_127(rport_io_ins_127),
    .io_ins_128(rport_io_ins_128),
    .io_ins_129(rport_io_ins_129),
    .io_ins_130(rport_io_ins_130),
    .io_ins_131(rport_io_ins_131),
    .io_ins_132(rport_io_ins_132),
    .io_ins_133(rport_io_ins_133),
    .io_ins_134(rport_io_ins_134),
    .io_ins_135(rport_io_ins_135),
    .io_ins_136(rport_io_ins_136),
    .io_ins_137(rport_io_ins_137),
    .io_ins_138(rport_io_ins_138),
    .io_ins_139(rport_io_ins_139),
    .io_ins_140(rport_io_ins_140),
    .io_ins_141(rport_io_ins_141),
    .io_ins_142(rport_io_ins_142),
    .io_ins_143(rport_io_ins_143),
    .io_ins_144(rport_io_ins_144),
    .io_ins_145(rport_io_ins_145),
    .io_ins_146(rport_io_ins_146),
    .io_ins_147(rport_io_ins_147),
    .io_ins_148(rport_io_ins_148),
    .io_ins_149(rport_io_ins_149),
    .io_ins_150(rport_io_ins_150),
    .io_ins_151(rport_io_ins_151),
    .io_ins_152(rport_io_ins_152),
    .io_ins_153(rport_io_ins_153),
    .io_ins_154(rport_io_ins_154),
    .io_ins_155(rport_io_ins_155),
    .io_ins_156(rport_io_ins_156),
    .io_ins_157(rport_io_ins_157),
    .io_ins_158(rport_io_ins_158),
    .io_ins_159(rport_io_ins_159),
    .io_ins_160(rport_io_ins_160),
    .io_ins_161(rport_io_ins_161),
    .io_ins_162(rport_io_ins_162),
    .io_ins_163(rport_io_ins_163),
    .io_ins_164(rport_io_ins_164),
    .io_ins_165(rport_io_ins_165),
    .io_ins_166(rport_io_ins_166),
    .io_ins_167(rport_io_ins_167),
    .io_ins_168(rport_io_ins_168),
    .io_ins_169(rport_io_ins_169),
    .io_ins_170(rport_io_ins_170),
    .io_ins_171(rport_io_ins_171),
    .io_ins_172(rport_io_ins_172),
    .io_ins_173(rport_io_ins_173),
    .io_ins_174(rport_io_ins_174),
    .io_ins_175(rport_io_ins_175),
    .io_ins_176(rport_io_ins_176),
    .io_ins_177(rport_io_ins_177),
    .io_ins_178(rport_io_ins_178),
    .io_ins_179(rport_io_ins_179),
    .io_ins_180(rport_io_ins_180),
    .io_ins_181(rport_io_ins_181),
    .io_ins_182(rport_io_ins_182),
    .io_ins_183(rport_io_ins_183),
    .io_ins_184(rport_io_ins_184),
    .io_ins_185(rport_io_ins_185),
    .io_ins_186(rport_io_ins_186),
    .io_ins_187(rport_io_ins_187),
    .io_ins_188(rport_io_ins_188),
    .io_ins_189(rport_io_ins_189),
    .io_ins_190(rport_io_ins_190),
    .io_ins_191(rport_io_ins_191),
    .io_ins_192(rport_io_ins_192),
    .io_ins_193(rport_io_ins_193),
    .io_ins_194(rport_io_ins_194),
    .io_ins_195(rport_io_ins_195),
    .io_ins_196(rport_io_ins_196),
    .io_ins_197(rport_io_ins_197),
    .io_ins_198(rport_io_ins_198),
    .io_ins_199(rport_io_ins_199),
    .io_ins_200(rport_io_ins_200),
    .io_ins_201(rport_io_ins_201),
    .io_ins_202(rport_io_ins_202),
    .io_ins_203(rport_io_ins_203),
    .io_ins_204(rport_io_ins_204),
    .io_ins_205(rport_io_ins_205),
    .io_ins_206(rport_io_ins_206),
    .io_ins_207(rport_io_ins_207),
    .io_ins_208(rport_io_ins_208),
    .io_ins_209(rport_io_ins_209),
    .io_ins_210(rport_io_ins_210),
    .io_ins_211(rport_io_ins_211),
    .io_ins_212(rport_io_ins_212),
    .io_ins_213(rport_io_ins_213),
    .io_ins_214(rport_io_ins_214),
    .io_ins_215(rport_io_ins_215),
    .io_ins_216(rport_io_ins_216),
    .io_ins_217(rport_io_ins_217),
    .io_ins_218(rport_io_ins_218),
    .io_ins_219(rport_io_ins_219),
    .io_ins_220(rport_io_ins_220),
    .io_ins_221(rport_io_ins_221),
    .io_ins_222(rport_io_ins_222),
    .io_ins_223(rport_io_ins_223),
    .io_ins_224(rport_io_ins_224),
    .io_ins_225(rport_io_ins_225),
    .io_ins_226(rport_io_ins_226),
    .io_ins_227(rport_io_ins_227),
    .io_ins_228(rport_io_ins_228),
    .io_ins_229(rport_io_ins_229),
    .io_ins_230(rport_io_ins_230),
    .io_ins_231(rport_io_ins_231),
    .io_ins_232(rport_io_ins_232),
    .io_ins_233(rport_io_ins_233),
    .io_ins_234(rport_io_ins_234),
    .io_ins_235(rport_io_ins_235),
    .io_ins_236(rport_io_ins_236),
    .io_ins_237(rport_io_ins_237),
    .io_ins_238(rport_io_ins_238),
    .io_ins_239(rport_io_ins_239),
    .io_ins_240(rport_io_ins_240),
    .io_ins_241(rport_io_ins_241),
    .io_ins_242(rport_io_ins_242),
    .io_ins_243(rport_io_ins_243),
    .io_ins_244(rport_io_ins_244),
    .io_ins_245(rport_io_ins_245),
    .io_ins_246(rport_io_ins_246),
    .io_ins_247(rport_io_ins_247),
    .io_ins_248(rport_io_ins_248),
    .io_ins_249(rport_io_ins_249),
    .io_ins_250(rport_io_ins_250),
    .io_ins_251(rport_io_ins_251),
    .io_ins_252(rport_io_ins_252),
    .io_ins_253(rport_io_ins_253),
    .io_ins_254(rport_io_ins_254),
    .io_ins_255(rport_io_ins_255),
    .io_ins_256(rport_io_ins_256),
    .io_ins_257(rport_io_ins_257),
    .io_ins_258(rport_io_ins_258),
    .io_ins_259(rport_io_ins_259),
    .io_ins_260(rport_io_ins_260),
    .io_ins_261(rport_io_ins_261),
    .io_ins_262(rport_io_ins_262),
    .io_ins_263(rport_io_ins_263),
    .io_ins_264(rport_io_ins_264),
    .io_ins_265(rport_io_ins_265),
    .io_ins_266(rport_io_ins_266),
    .io_ins_267(rport_io_ins_267),
    .io_ins_268(rport_io_ins_268),
    .io_ins_269(rport_io_ins_269),
    .io_ins_270(rport_io_ins_270),
    .io_ins_271(rport_io_ins_271),
    .io_ins_272(rport_io_ins_272),
    .io_ins_273(rport_io_ins_273),
    .io_ins_274(rport_io_ins_274),
    .io_ins_275(rport_io_ins_275),
    .io_ins_276(rport_io_ins_276),
    .io_ins_277(rport_io_ins_277),
    .io_ins_278(rport_io_ins_278),
    .io_ins_279(rport_io_ins_279),
    .io_ins_280(rport_io_ins_280),
    .io_ins_281(rport_io_ins_281),
    .io_ins_282(rport_io_ins_282),
    .io_ins_283(rport_io_ins_283),
    .io_ins_284(rport_io_ins_284),
    .io_ins_285(rport_io_ins_285),
    .io_ins_286(rport_io_ins_286),
    .io_ins_287(rport_io_ins_287),
    .io_ins_288(rport_io_ins_288),
    .io_ins_289(rport_io_ins_289),
    .io_ins_290(rport_io_ins_290),
    .io_ins_291(rport_io_ins_291),
    .io_ins_292(rport_io_ins_292),
    .io_ins_293(rport_io_ins_293),
    .io_ins_294(rport_io_ins_294),
    .io_ins_295(rport_io_ins_295),
    .io_ins_296(rport_io_ins_296),
    .io_ins_297(rport_io_ins_297),
    .io_ins_298(rport_io_ins_298),
    .io_ins_299(rport_io_ins_299),
    .io_ins_300(rport_io_ins_300),
    .io_ins_301(rport_io_ins_301),
    .io_ins_302(rport_io_ins_302),
    .io_ins_303(rport_io_ins_303),
    .io_ins_304(rport_io_ins_304),
    .io_ins_305(rport_io_ins_305),
    .io_ins_306(rport_io_ins_306),
    .io_ins_307(rport_io_ins_307),
    .io_ins_308(rport_io_ins_308),
    .io_ins_309(rport_io_ins_309),
    .io_ins_310(rport_io_ins_310),
    .io_ins_311(rport_io_ins_311),
    .io_ins_312(rport_io_ins_312),
    .io_ins_313(rport_io_ins_313),
    .io_ins_314(rport_io_ins_314),
    .io_ins_315(rport_io_ins_315),
    .io_ins_316(rport_io_ins_316),
    .io_ins_317(rport_io_ins_317),
    .io_ins_318(rport_io_ins_318),
    .io_ins_319(rport_io_ins_319),
    .io_ins_320(rport_io_ins_320),
    .io_ins_321(rport_io_ins_321),
    .io_ins_322(rport_io_ins_322),
    .io_ins_323(rport_io_ins_323),
    .io_ins_324(rport_io_ins_324),
    .io_ins_325(rport_io_ins_325),
    .io_ins_326(rport_io_ins_326),
    .io_ins_327(rport_io_ins_327),
    .io_ins_328(rport_io_ins_328),
    .io_ins_329(rport_io_ins_329),
    .io_ins_330(rport_io_ins_330),
    .io_ins_331(rport_io_ins_331),
    .io_ins_332(rport_io_ins_332),
    .io_ins_333(rport_io_ins_333),
    .io_ins_334(rport_io_ins_334),
    .io_ins_335(rport_io_ins_335),
    .io_ins_336(rport_io_ins_336),
    .io_ins_337(rport_io_ins_337),
    .io_ins_338(rport_io_ins_338),
    .io_ins_339(rport_io_ins_339),
    .io_ins_340(rport_io_ins_340),
    .io_ins_341(rport_io_ins_341),
    .io_ins_342(rport_io_ins_342),
    .io_ins_343(rport_io_ins_343),
    .io_ins_344(rport_io_ins_344),
    .io_ins_345(rport_io_ins_345),
    .io_ins_346(rport_io_ins_346),
    .io_ins_347(rport_io_ins_347),
    .io_ins_348(rport_io_ins_348),
    .io_ins_349(rport_io_ins_349),
    .io_ins_350(rport_io_ins_350),
    .io_ins_351(rport_io_ins_351),
    .io_ins_352(rport_io_ins_352),
    .io_ins_353(rport_io_ins_353),
    .io_ins_354(rport_io_ins_354),
    .io_ins_355(rport_io_ins_355),
    .io_ins_356(rport_io_ins_356),
    .io_ins_357(rport_io_ins_357),
    .io_ins_358(rport_io_ins_358),
    .io_ins_359(rport_io_ins_359),
    .io_ins_360(rport_io_ins_360),
    .io_ins_361(rport_io_ins_361),
    .io_ins_362(rport_io_ins_362),
    .io_ins_363(rport_io_ins_363),
    .io_ins_364(rport_io_ins_364),
    .io_ins_365(rport_io_ins_365),
    .io_ins_366(rport_io_ins_366),
    .io_ins_367(rport_io_ins_367),
    .io_ins_368(rport_io_ins_368),
    .io_ins_369(rport_io_ins_369),
    .io_ins_370(rport_io_ins_370),
    .io_ins_371(rport_io_ins_371),
    .io_ins_372(rport_io_ins_372),
    .io_ins_373(rport_io_ins_373),
    .io_ins_374(rport_io_ins_374),
    .io_ins_375(rport_io_ins_375),
    .io_ins_376(rport_io_ins_376),
    .io_ins_377(rport_io_ins_377),
    .io_ins_378(rport_io_ins_378),
    .io_ins_379(rport_io_ins_379),
    .io_ins_380(rport_io_ins_380),
    .io_ins_381(rport_io_ins_381),
    .io_ins_382(rport_io_ins_382),
    .io_ins_383(rport_io_ins_383),
    .io_ins_384(rport_io_ins_384),
    .io_ins_385(rport_io_ins_385),
    .io_ins_386(rport_io_ins_386),
    .io_ins_387(rport_io_ins_387),
    .io_ins_388(rport_io_ins_388),
    .io_ins_389(rport_io_ins_389),
    .io_ins_390(rport_io_ins_390),
    .io_ins_391(rport_io_ins_391),
    .io_ins_392(rport_io_ins_392),
    .io_ins_393(rport_io_ins_393),
    .io_ins_394(rport_io_ins_394),
    .io_ins_395(rport_io_ins_395),
    .io_ins_396(rport_io_ins_396),
    .io_ins_397(rport_io_ins_397),
    .io_ins_398(rport_io_ins_398),
    .io_ins_399(rport_io_ins_399),
    .io_ins_400(rport_io_ins_400),
    .io_ins_401(rport_io_ins_401),
    .io_ins_402(rport_io_ins_402),
    .io_ins_403(rport_io_ins_403),
    .io_ins_404(rport_io_ins_404),
    .io_ins_405(rport_io_ins_405),
    .io_ins_406(rport_io_ins_406),
    .io_ins_407(rport_io_ins_407),
    .io_ins_408(rport_io_ins_408),
    .io_ins_409(rport_io_ins_409),
    .io_ins_410(rport_io_ins_410),
    .io_ins_411(rport_io_ins_411),
    .io_ins_412(rport_io_ins_412),
    .io_ins_413(rport_io_ins_413),
    .io_ins_414(rport_io_ins_414),
    .io_ins_415(rport_io_ins_415),
    .io_ins_416(rport_io_ins_416),
    .io_ins_417(rport_io_ins_417),
    .io_ins_418(rport_io_ins_418),
    .io_ins_419(rport_io_ins_419),
    .io_ins_420(rport_io_ins_420),
    .io_ins_421(rport_io_ins_421),
    .io_ins_422(rport_io_ins_422),
    .io_ins_423(rport_io_ins_423),
    .io_ins_424(rport_io_ins_424),
    .io_ins_425(rport_io_ins_425),
    .io_ins_426(rport_io_ins_426),
    .io_ins_427(rport_io_ins_427),
    .io_ins_428(rport_io_ins_428),
    .io_ins_429(rport_io_ins_429),
    .io_ins_430(rport_io_ins_430),
    .io_ins_431(rport_io_ins_431),
    .io_ins_432(rport_io_ins_432),
    .io_ins_433(rport_io_ins_433),
    .io_ins_434(rport_io_ins_434),
    .io_ins_435(rport_io_ins_435),
    .io_ins_436(rport_io_ins_436),
    .io_ins_437(rport_io_ins_437),
    .io_ins_438(rport_io_ins_438),
    .io_ins_439(rport_io_ins_439),
    .io_ins_440(rport_io_ins_440),
    .io_ins_441(rport_io_ins_441),
    .io_ins_442(rport_io_ins_442),
    .io_ins_443(rport_io_ins_443),
    .io_ins_444(rport_io_ins_444),
    .io_ins_445(rport_io_ins_445),
    .io_ins_446(rport_io_ins_446),
    .io_ins_447(rport_io_ins_447),
    .io_ins_448(rport_io_ins_448),
    .io_ins_449(rport_io_ins_449),
    .io_ins_450(rport_io_ins_450),
    .io_ins_451(rport_io_ins_451),
    .io_ins_452(rport_io_ins_452),
    .io_ins_453(rport_io_ins_453),
    .io_ins_454(rport_io_ins_454),
    .io_ins_455(rport_io_ins_455),
    .io_ins_456(rport_io_ins_456),
    .io_ins_457(rport_io_ins_457),
    .io_ins_458(rport_io_ins_458),
    .io_ins_459(rport_io_ins_459),
    .io_ins_460(rport_io_ins_460),
    .io_ins_461(rport_io_ins_461),
    .io_ins_462(rport_io_ins_462),
    .io_ins_463(rport_io_ins_463),
    .io_ins_464(rport_io_ins_464),
    .io_ins_465(rport_io_ins_465),
    .io_ins_466(rport_io_ins_466),
    .io_ins_467(rport_io_ins_467),
    .io_ins_468(rport_io_ins_468),
    .io_ins_469(rport_io_ins_469),
    .io_ins_470(rport_io_ins_470),
    .io_ins_471(rport_io_ins_471),
    .io_ins_472(rport_io_ins_472),
    .io_ins_473(rport_io_ins_473),
    .io_ins_474(rport_io_ins_474),
    .io_ins_475(rport_io_ins_475),
    .io_ins_476(rport_io_ins_476),
    .io_ins_477(rport_io_ins_477),
    .io_ins_478(rport_io_ins_478),
    .io_ins_479(rport_io_ins_479),
    .io_ins_480(rport_io_ins_480),
    .io_ins_481(rport_io_ins_481),
    .io_ins_482(rport_io_ins_482),
    .io_ins_483(rport_io_ins_483),
    .io_ins_484(rport_io_ins_484),
    .io_ins_485(rport_io_ins_485),
    .io_ins_486(rport_io_ins_486),
    .io_ins_487(rport_io_ins_487),
    .io_ins_488(rport_io_ins_488),
    .io_ins_489(rport_io_ins_489),
    .io_ins_490(rport_io_ins_490),
    .io_ins_491(rport_io_ins_491),
    .io_ins_492(rport_io_ins_492),
    .io_ins_493(rport_io_ins_493),
    .io_ins_494(rport_io_ins_494),
    .io_ins_495(rport_io_ins_495),
    .io_ins_496(rport_io_ins_496),
    .io_ins_497(rport_io_ins_497),
    .io_ins_498(rport_io_ins_498),
    .io_ins_499(rport_io_ins_499),
    .io_ins_500(rport_io_ins_500),
    .io_ins_501(rport_io_ins_501),
    .io_ins_502(rport_io_ins_502),
    .io_ins_503(rport_io_ins_503),
    .io_ins_504(rport_io_ins_504),
    .io_ins_505(rport_io_ins_505),
    .io_ins_506(rport_io_ins_506),
    .io_ins_507(rport_io_ins_507),
    .io_ins_508(rport_io_ins_508),
    .io_ins_509(rport_io_ins_509),
    .io_ins_510(rport_io_ins_510),
    .io_ins_511(rport_io_ins_511),
    .io_ins_512(rport_io_ins_512),
    .io_ins_513(rport_io_ins_513),
    .io_ins_514(rport_io_ins_514),
    .io_ins_515(rport_io_ins_515),
    .io_ins_516(rport_io_ins_516),
    .io_ins_517(rport_io_ins_517),
    .io_ins_518(rport_io_ins_518),
    .io_ins_519(rport_io_ins_519),
    .io_ins_520(rport_io_ins_520),
    .io_ins_521(rport_io_ins_521),
    .io_ins_522(rport_io_ins_522),
    .io_ins_523(rport_io_ins_523),
    .io_ins_524(rport_io_ins_524),
    .io_ins_525(rport_io_ins_525),
    .io_ins_526(rport_io_ins_526),
    .io_ins_527(rport_io_ins_527),
    .io_ins_528(rport_io_ins_528),
    .io_ins_529(rport_io_ins_529),
    .io_ins_530(rport_io_ins_530),
    .io_ins_531(rport_io_ins_531),
    .io_ins_532(rport_io_ins_532),
    .io_ins_533(rport_io_ins_533),
    .io_sel(rport_io_sel),
    .io_out(rport_io_out)
  );
  assign _T_3262 = io_waddr == 32'h0; // @[RegFile.scala 80:42:@41723.4]
  assign _T_3268 = io_waddr == 32'h1; // @[RegFile.scala 68:46:@41735.4]
  assign _T_3269 = io_wen & _T_3268; // @[RegFile.scala 68:34:@41736.4]
  assign _T_3282 = io_waddr == 32'h2; // @[RegFile.scala 80:42:@41754.4]
  assign _T_3288 = io_waddr == 32'h3; // @[RegFile.scala 74:80:@41766.4]
  assign _T_3289 = io_wen & _T_3288; // @[RegFile.scala 74:68:@41767.4]
  assign _T_3295 = io_waddr == 32'h4; // @[RegFile.scala 74:80:@41780.4]
  assign _T_3296 = io_wen & _T_3295; // @[RegFile.scala 74:68:@41781.4]
  assign _T_3302 = io_waddr == 32'h5; // @[RegFile.scala 74:80:@41794.4]
  assign _T_3303 = io_wen & _T_3302; // @[RegFile.scala 74:68:@41795.4]
  assign _T_3309 = io_waddr == 32'h6; // @[RegFile.scala 74:80:@41808.4]
  assign _T_3310 = io_wen & _T_3309; // @[RegFile.scala 74:68:@41809.4]
  assign _T_3316 = io_waddr == 32'h7; // @[RegFile.scala 74:80:@41822.4]
  assign _T_3317 = io_wen & _T_3316; // @[RegFile.scala 74:68:@41823.4]
  assign _T_3323 = io_waddr == 32'h8; // @[RegFile.scala 74:80:@41836.4]
  assign _T_3324 = io_wen & _T_3323; // @[RegFile.scala 74:68:@41837.4]
  assign _T_3330 = io_waddr == 32'h9; // @[RegFile.scala 74:80:@41850.4]
  assign _T_3331 = io_wen & _T_3330; // @[RegFile.scala 74:68:@41851.4]
  assign _T_3337 = io_waddr == 32'ha; // @[RegFile.scala 74:80:@41864.4]
  assign _T_3338 = io_wen & _T_3337; // @[RegFile.scala 74:68:@41865.4]
  assign _T_3344 = io_waddr == 32'hb; // @[RegFile.scala 74:80:@41878.4]
  assign _T_3345 = io_wen & _T_3344; // @[RegFile.scala 74:68:@41879.4]
  assign _T_3351 = io_waddr == 32'hc; // @[RegFile.scala 74:80:@41892.4]
  assign _T_3352 = io_wen & _T_3351; // @[RegFile.scala 74:68:@41893.4]
  assign _T_3358 = io_waddr == 32'hd; // @[RegFile.scala 74:80:@41906.4]
  assign _T_3359 = io_wen & _T_3358; // @[RegFile.scala 74:68:@41907.4]
  assign _T_3365 = io_waddr == 32'he; // @[RegFile.scala 74:80:@41920.4]
  assign _T_3366 = io_wen & _T_3365; // @[RegFile.scala 74:68:@41921.4]
  assign _T_3372 = io_waddr == 32'hf; // @[RegFile.scala 74:80:@41934.4]
  assign _T_3373 = io_wen & _T_3372; // @[RegFile.scala 74:68:@41935.4]
  assign _T_3379 = io_waddr == 32'h10; // @[RegFile.scala 74:80:@41948.4]
  assign _T_3380 = io_wen & _T_3379; // @[RegFile.scala 74:68:@41949.4]
  assign _T_3386 = io_waddr == 32'h11; // @[RegFile.scala 74:80:@41962.4]
  assign _T_3387 = io_wen & _T_3386; // @[RegFile.scala 74:68:@41963.4]
  assign _T_3393 = io_waddr == 32'h12; // @[RegFile.scala 74:80:@41976.4]
  assign _T_3394 = io_wen & _T_3393; // @[RegFile.scala 74:68:@41977.4]
  assign _T_3400 = io_waddr == 32'h13; // @[RegFile.scala 74:80:@41990.4]
  assign _T_3401 = io_wen & _T_3400; // @[RegFile.scala 74:68:@41991.4]
  assign _T_3407 = io_waddr == 32'h14; // @[RegFile.scala 74:80:@42004.4]
  assign _T_3408 = io_wen & _T_3407; // @[RegFile.scala 74:68:@42005.4]
  assign _T_3414 = io_waddr == 32'h15; // @[RegFile.scala 74:80:@42018.4]
  assign _T_3415 = io_wen & _T_3414; // @[RegFile.scala 74:68:@42019.4]
  assign _T_3421 = io_waddr == 32'h16; // @[RegFile.scala 74:80:@42032.4]
  assign _T_3422 = io_wen & _T_3421; // @[RegFile.scala 74:68:@42033.4]
  assign _T_3428 = io_waddr == 32'h17; // @[RegFile.scala 74:80:@42046.4]
  assign _T_3429 = io_wen & _T_3428; // @[RegFile.scala 74:68:@42047.4]
  assign _T_3435 = io_waddr == 32'h18; // @[RegFile.scala 74:80:@42060.4]
  assign _T_3436 = io_wen & _T_3435; // @[RegFile.scala 74:68:@42061.4]
  assign _T_3442 = io_waddr == 32'h19; // @[RegFile.scala 74:80:@42074.4]
  assign _T_3443 = io_wen & _T_3442; // @[RegFile.scala 74:68:@42075.4]
  assign _T_3449 = io_waddr == 32'h1a; // @[RegFile.scala 74:80:@42088.4]
  assign _T_3450 = io_wen & _T_3449; // @[RegFile.scala 74:68:@42089.4]
  assign _T_3456 = io_waddr == 32'h1b; // @[RegFile.scala 74:80:@42102.4]
  assign _T_3457 = io_wen & _T_3456; // @[RegFile.scala 74:68:@42103.4]
  assign _T_3463 = io_waddr == 32'h1c; // @[RegFile.scala 74:80:@42116.4]
  assign _T_3464 = io_wen & _T_3463; // @[RegFile.scala 74:68:@42117.4]
  assign _T_3470 = io_waddr == 32'h1d; // @[RegFile.scala 74:80:@42130.4]
  assign _T_3471 = io_wen & _T_3470; // @[RegFile.scala 74:68:@42131.4]
  assign _T_3477 = io_waddr == 32'h1e; // @[RegFile.scala 74:80:@42144.4]
  assign _T_3478 = io_wen & _T_3477; // @[RegFile.scala 74:68:@42145.4]
  assign _T_3484 = io_waddr == 32'h1f; // @[RegFile.scala 74:80:@42158.4]
  assign _T_3485 = io_wen & _T_3484; // @[RegFile.scala 74:68:@42159.4]
  assign _T_3491 = io_waddr == 32'h20; // @[RegFile.scala 74:80:@42172.4]
  assign _T_3492 = io_wen & _T_3491; // @[RegFile.scala 74:68:@42173.4]
  assign _T_3498 = io_waddr == 32'h21; // @[RegFile.scala 74:80:@42186.4]
  assign _T_3499 = io_wen & _T_3498; // @[RegFile.scala 74:68:@42187.4]
  assign _T_3505 = io_waddr == 32'h22; // @[RegFile.scala 74:80:@42200.4]
  assign _T_3506 = io_wen & _T_3505; // @[RegFile.scala 74:68:@42201.4]
  assign io_rdata = rport_io_out; // @[RegFile.scala 107:14:@50270.4]
  assign io_argIns_0 = regs_0_io_out; // @[RegFile.scala 111:13:@50275.4]
  assign io_argIns_1 = regs_1_io_out; // @[RegFile.scala 111:13:@50276.4]
  assign io_argIns_2 = regs_2_io_out; // @[RegFile.scala 111:13:@50277.4]
  assign regs_0_clock = clock; // @[:@41721.4]
  assign regs_0_reset = reset; // @[:@41722.4 RegFile.scala 82:16:@41728.4]
  assign regs_0_io_in = io_wdata; // @[RegFile.scala 81:16:@41726.4]
  assign regs_0_io_reset = reset; // @[RegFile.scala 83:19:@41730.4]
  assign regs_0_io_enable = io_wen & _T_3262; // @[RegFile.scala 80:20:@41725.4]
  assign regs_1_clock = clock; // @[:@41733.4]
  assign regs_1_reset = reset; // @[:@41734.4 RegFile.scala 70:16:@41746.4]
  assign regs_1_io_in = _T_3269 ? io_wdata : io_argOuts_0_bits; // @[RegFile.scala 69:16:@41744.4]
  assign regs_1_io_reset = reset; // @[RegFile.scala 72:19:@41749.4]
  assign regs_1_io_enable = _T_3269 ? _T_3269 : io_argOuts_0_valid; // @[RegFile.scala 68:20:@41740.4]
  assign regs_2_clock = clock; // @[:@41752.4]
  assign regs_2_reset = reset; // @[:@41753.4 RegFile.scala 82:16:@41759.4]
  assign regs_2_io_in = io_wdata; // @[RegFile.scala 81:16:@41757.4]
  assign regs_2_io_reset = reset; // @[RegFile.scala 83:19:@41761.4]
  assign regs_2_io_enable = io_wen & _T_3282; // @[RegFile.scala 80:20:@41756.4]
  assign regs_3_clock = clock; // @[:@41764.4]
  assign regs_3_reset = io_reset; // @[:@41765.4 RegFile.scala 76:16:@41772.4]
  assign regs_3_io_in = io_argOuts_1_valid ? io_argOuts_1_bits : io_wdata; // @[RegFile.scala 75:16:@41771.4]
  assign regs_3_io_reset = reset; // @[RegFile.scala 78:19:@41775.4]
  assign regs_3_io_enable = io_argOuts_1_valid | _T_3289; // @[RegFile.scala 74:20:@41769.4]
  assign regs_4_clock = clock; // @[:@41778.4]
  assign regs_4_reset = io_reset; // @[:@41779.4 RegFile.scala 76:16:@41786.4]
  assign regs_4_io_in = io_argOuts_2_valid ? io_argOuts_2_bits : io_wdata; // @[RegFile.scala 75:16:@41785.4]
  assign regs_4_io_reset = reset; // @[RegFile.scala 78:19:@41789.4]
  assign regs_4_io_enable = io_argOuts_2_valid | _T_3296; // @[RegFile.scala 74:20:@41783.4]
  assign regs_5_clock = clock; // @[:@41792.4]
  assign regs_5_reset = io_reset; // @[:@41793.4 RegFile.scala 76:16:@41800.4]
  assign regs_5_io_in = io_argOuts_3_valid ? io_argOuts_3_bits : io_wdata; // @[RegFile.scala 75:16:@41799.4]
  assign regs_5_io_reset = reset; // @[RegFile.scala 78:19:@41803.4]
  assign regs_5_io_enable = io_argOuts_3_valid | _T_3303; // @[RegFile.scala 74:20:@41797.4]
  assign regs_6_clock = clock; // @[:@41806.4]
  assign regs_6_reset = io_reset; // @[:@41807.4 RegFile.scala 76:16:@41814.4]
  assign regs_6_io_in = io_argOuts_4_valid ? io_argOuts_4_bits : io_wdata; // @[RegFile.scala 75:16:@41813.4]
  assign regs_6_io_reset = reset; // @[RegFile.scala 78:19:@41817.4]
  assign regs_6_io_enable = io_argOuts_4_valid | _T_3310; // @[RegFile.scala 74:20:@41811.4]
  assign regs_7_clock = clock; // @[:@41820.4]
  assign regs_7_reset = io_reset; // @[:@41821.4 RegFile.scala 76:16:@41828.4]
  assign regs_7_io_in = io_argOuts_5_valid ? io_argOuts_5_bits : io_wdata; // @[RegFile.scala 75:16:@41827.4]
  assign regs_7_io_reset = reset; // @[RegFile.scala 78:19:@41831.4]
  assign regs_7_io_enable = io_argOuts_5_valid | _T_3317; // @[RegFile.scala 74:20:@41825.4]
  assign regs_8_clock = clock; // @[:@41834.4]
  assign regs_8_reset = io_reset; // @[:@41835.4 RegFile.scala 76:16:@41842.4]
  assign regs_8_io_in = io_argOuts_6_valid ? io_argOuts_6_bits : io_wdata; // @[RegFile.scala 75:16:@41841.4]
  assign regs_8_io_reset = reset; // @[RegFile.scala 78:19:@41845.4]
  assign regs_8_io_enable = io_argOuts_6_valid | _T_3324; // @[RegFile.scala 74:20:@41839.4]
  assign regs_9_clock = clock; // @[:@41848.4]
  assign regs_9_reset = io_reset; // @[:@41849.4 RegFile.scala 76:16:@41856.4]
  assign regs_9_io_in = io_argOuts_7_valid ? io_argOuts_7_bits : io_wdata; // @[RegFile.scala 75:16:@41855.4]
  assign regs_9_io_reset = reset; // @[RegFile.scala 78:19:@41859.4]
  assign regs_9_io_enable = io_argOuts_7_valid | _T_3331; // @[RegFile.scala 74:20:@41853.4]
  assign regs_10_clock = clock; // @[:@41862.4]
  assign regs_10_reset = io_reset; // @[:@41863.4 RegFile.scala 76:16:@41870.4]
  assign regs_10_io_in = io_argOuts_8_valid ? io_argOuts_8_bits : io_wdata; // @[RegFile.scala 75:16:@41869.4]
  assign regs_10_io_reset = reset; // @[RegFile.scala 78:19:@41873.4]
  assign regs_10_io_enable = io_argOuts_8_valid | _T_3338; // @[RegFile.scala 74:20:@41867.4]
  assign regs_11_clock = clock; // @[:@41876.4]
  assign regs_11_reset = io_reset; // @[:@41877.4 RegFile.scala 76:16:@41884.4]
  assign regs_11_io_in = io_argOuts_9_valid ? io_argOuts_9_bits : io_wdata; // @[RegFile.scala 75:16:@41883.4]
  assign regs_11_io_reset = reset; // @[RegFile.scala 78:19:@41887.4]
  assign regs_11_io_enable = io_argOuts_9_valid | _T_3345; // @[RegFile.scala 74:20:@41881.4]
  assign regs_12_clock = clock; // @[:@41890.4]
  assign regs_12_reset = io_reset; // @[:@41891.4 RegFile.scala 76:16:@41898.4]
  assign regs_12_io_in = io_argOuts_10_valid ? io_argOuts_10_bits : io_wdata; // @[RegFile.scala 75:16:@41897.4]
  assign regs_12_io_reset = reset; // @[RegFile.scala 78:19:@41901.4]
  assign regs_12_io_enable = io_argOuts_10_valid | _T_3352; // @[RegFile.scala 74:20:@41895.4]
  assign regs_13_clock = clock; // @[:@41904.4]
  assign regs_13_reset = io_reset; // @[:@41905.4 RegFile.scala 76:16:@41912.4]
  assign regs_13_io_in = io_argOuts_11_valid ? io_argOuts_11_bits : io_wdata; // @[RegFile.scala 75:16:@41911.4]
  assign regs_13_io_reset = reset; // @[RegFile.scala 78:19:@41915.4]
  assign regs_13_io_enable = io_argOuts_11_valid | _T_3359; // @[RegFile.scala 74:20:@41909.4]
  assign regs_14_clock = clock; // @[:@41918.4]
  assign regs_14_reset = io_reset; // @[:@41919.4 RegFile.scala 76:16:@41926.4]
  assign regs_14_io_in = io_argOuts_12_valid ? io_argOuts_12_bits : io_wdata; // @[RegFile.scala 75:16:@41925.4]
  assign regs_14_io_reset = reset; // @[RegFile.scala 78:19:@41929.4]
  assign regs_14_io_enable = io_argOuts_12_valid | _T_3366; // @[RegFile.scala 74:20:@41923.4]
  assign regs_15_clock = clock; // @[:@41932.4]
  assign regs_15_reset = io_reset; // @[:@41933.4 RegFile.scala 76:16:@41940.4]
  assign regs_15_io_in = io_argOuts_13_valid ? io_argOuts_13_bits : io_wdata; // @[RegFile.scala 75:16:@41939.4]
  assign regs_15_io_reset = reset; // @[RegFile.scala 78:19:@41943.4]
  assign regs_15_io_enable = io_argOuts_13_valid | _T_3373; // @[RegFile.scala 74:20:@41937.4]
  assign regs_16_clock = clock; // @[:@41946.4]
  assign regs_16_reset = io_reset; // @[:@41947.4 RegFile.scala 76:16:@41954.4]
  assign regs_16_io_in = io_argOuts_14_valid ? io_argOuts_14_bits : io_wdata; // @[RegFile.scala 75:16:@41953.4]
  assign regs_16_io_reset = reset; // @[RegFile.scala 78:19:@41957.4]
  assign regs_16_io_enable = io_argOuts_14_valid | _T_3380; // @[RegFile.scala 74:20:@41951.4]
  assign regs_17_clock = clock; // @[:@41960.4]
  assign regs_17_reset = io_reset; // @[:@41961.4 RegFile.scala 76:16:@41968.4]
  assign regs_17_io_in = io_argOuts_15_valid ? io_argOuts_15_bits : io_wdata; // @[RegFile.scala 75:16:@41967.4]
  assign regs_17_io_reset = reset; // @[RegFile.scala 78:19:@41971.4]
  assign regs_17_io_enable = io_argOuts_15_valid | _T_3387; // @[RegFile.scala 74:20:@41965.4]
  assign regs_18_clock = clock; // @[:@41974.4]
  assign regs_18_reset = io_reset; // @[:@41975.4 RegFile.scala 76:16:@41982.4]
  assign regs_18_io_in = io_argOuts_16_valid ? io_argOuts_16_bits : io_wdata; // @[RegFile.scala 75:16:@41981.4]
  assign regs_18_io_reset = reset; // @[RegFile.scala 78:19:@41985.4]
  assign regs_18_io_enable = io_argOuts_16_valid | _T_3394; // @[RegFile.scala 74:20:@41979.4]
  assign regs_19_clock = clock; // @[:@41988.4]
  assign regs_19_reset = io_reset; // @[:@41989.4 RegFile.scala 76:16:@41996.4]
  assign regs_19_io_in = io_argOuts_17_valid ? io_argOuts_17_bits : io_wdata; // @[RegFile.scala 75:16:@41995.4]
  assign regs_19_io_reset = reset; // @[RegFile.scala 78:19:@41999.4]
  assign regs_19_io_enable = io_argOuts_17_valid | _T_3401; // @[RegFile.scala 74:20:@41993.4]
  assign regs_20_clock = clock; // @[:@42002.4]
  assign regs_20_reset = io_reset; // @[:@42003.4 RegFile.scala 76:16:@42010.4]
  assign regs_20_io_in = io_argOuts_18_valid ? io_argOuts_18_bits : io_wdata; // @[RegFile.scala 75:16:@42009.4]
  assign regs_20_io_reset = reset; // @[RegFile.scala 78:19:@42013.4]
  assign regs_20_io_enable = io_argOuts_18_valid | _T_3408; // @[RegFile.scala 74:20:@42007.4]
  assign regs_21_clock = clock; // @[:@42016.4]
  assign regs_21_reset = io_reset; // @[:@42017.4 RegFile.scala 76:16:@42024.4]
  assign regs_21_io_in = io_argOuts_19_valid ? io_argOuts_19_bits : io_wdata; // @[RegFile.scala 75:16:@42023.4]
  assign regs_21_io_reset = reset; // @[RegFile.scala 78:19:@42027.4]
  assign regs_21_io_enable = io_argOuts_19_valid | _T_3415; // @[RegFile.scala 74:20:@42021.4]
  assign regs_22_clock = clock; // @[:@42030.4]
  assign regs_22_reset = io_reset; // @[:@42031.4 RegFile.scala 76:16:@42038.4]
  assign regs_22_io_in = io_argOuts_20_valid ? io_argOuts_20_bits : io_wdata; // @[RegFile.scala 75:16:@42037.4]
  assign regs_22_io_reset = reset; // @[RegFile.scala 78:19:@42041.4]
  assign regs_22_io_enable = io_argOuts_20_valid | _T_3422; // @[RegFile.scala 74:20:@42035.4]
  assign regs_23_clock = clock; // @[:@42044.4]
  assign regs_23_reset = io_reset; // @[:@42045.4 RegFile.scala 76:16:@42052.4]
  assign regs_23_io_in = io_argOuts_21_valid ? io_argOuts_21_bits : io_wdata; // @[RegFile.scala 75:16:@42051.4]
  assign regs_23_io_reset = reset; // @[RegFile.scala 78:19:@42055.4]
  assign regs_23_io_enable = io_argOuts_21_valid | _T_3429; // @[RegFile.scala 74:20:@42049.4]
  assign regs_24_clock = clock; // @[:@42058.4]
  assign regs_24_reset = io_reset; // @[:@42059.4 RegFile.scala 76:16:@42066.4]
  assign regs_24_io_in = io_argOuts_22_valid ? io_argOuts_22_bits : io_wdata; // @[RegFile.scala 75:16:@42065.4]
  assign regs_24_io_reset = reset; // @[RegFile.scala 78:19:@42069.4]
  assign regs_24_io_enable = io_argOuts_22_valid | _T_3436; // @[RegFile.scala 74:20:@42063.4]
  assign regs_25_clock = clock; // @[:@42072.4]
  assign regs_25_reset = io_reset; // @[:@42073.4 RegFile.scala 76:16:@42080.4]
  assign regs_25_io_in = io_argOuts_23_valid ? io_argOuts_23_bits : io_wdata; // @[RegFile.scala 75:16:@42079.4]
  assign regs_25_io_reset = reset; // @[RegFile.scala 78:19:@42083.4]
  assign regs_25_io_enable = io_argOuts_23_valid | _T_3443; // @[RegFile.scala 74:20:@42077.4]
  assign regs_26_clock = clock; // @[:@42086.4]
  assign regs_26_reset = io_reset; // @[:@42087.4 RegFile.scala 76:16:@42094.4]
  assign regs_26_io_in = io_argOuts_24_valid ? io_argOuts_24_bits : io_wdata; // @[RegFile.scala 75:16:@42093.4]
  assign regs_26_io_reset = reset; // @[RegFile.scala 78:19:@42097.4]
  assign regs_26_io_enable = io_argOuts_24_valid | _T_3450; // @[RegFile.scala 74:20:@42091.4]
  assign regs_27_clock = clock; // @[:@42100.4]
  assign regs_27_reset = io_reset; // @[:@42101.4 RegFile.scala 76:16:@42108.4]
  assign regs_27_io_in = io_argOuts_25_valid ? io_argOuts_25_bits : io_wdata; // @[RegFile.scala 75:16:@42107.4]
  assign regs_27_io_reset = reset; // @[RegFile.scala 78:19:@42111.4]
  assign regs_27_io_enable = io_argOuts_25_valid | _T_3457; // @[RegFile.scala 74:20:@42105.4]
  assign regs_28_clock = clock; // @[:@42114.4]
  assign regs_28_reset = io_reset; // @[:@42115.4 RegFile.scala 76:16:@42122.4]
  assign regs_28_io_in = io_argOuts_26_valid ? io_argOuts_26_bits : io_wdata; // @[RegFile.scala 75:16:@42121.4]
  assign regs_28_io_reset = reset; // @[RegFile.scala 78:19:@42125.4]
  assign regs_28_io_enable = io_argOuts_26_valid | _T_3464; // @[RegFile.scala 74:20:@42119.4]
  assign regs_29_clock = clock; // @[:@42128.4]
  assign regs_29_reset = io_reset; // @[:@42129.4 RegFile.scala 76:16:@42136.4]
  assign regs_29_io_in = io_argOuts_27_valid ? io_argOuts_27_bits : io_wdata; // @[RegFile.scala 75:16:@42135.4]
  assign regs_29_io_reset = reset; // @[RegFile.scala 78:19:@42139.4]
  assign regs_29_io_enable = io_argOuts_27_valid | _T_3471; // @[RegFile.scala 74:20:@42133.4]
  assign regs_30_clock = clock; // @[:@42142.4]
  assign regs_30_reset = io_reset; // @[:@42143.4 RegFile.scala 76:16:@42150.4]
  assign regs_30_io_in = io_argOuts_28_valid ? io_argOuts_28_bits : io_wdata; // @[RegFile.scala 75:16:@42149.4]
  assign regs_30_io_reset = reset; // @[RegFile.scala 78:19:@42153.4]
  assign regs_30_io_enable = io_argOuts_28_valid | _T_3478; // @[RegFile.scala 74:20:@42147.4]
  assign regs_31_clock = clock; // @[:@42156.4]
  assign regs_31_reset = io_reset; // @[:@42157.4 RegFile.scala 76:16:@42164.4]
  assign regs_31_io_in = io_argOuts_29_valid ? io_argOuts_29_bits : io_wdata; // @[RegFile.scala 75:16:@42163.4]
  assign regs_31_io_reset = reset; // @[RegFile.scala 78:19:@42167.4]
  assign regs_31_io_enable = io_argOuts_29_valid | _T_3485; // @[RegFile.scala 74:20:@42161.4]
  assign regs_32_clock = clock; // @[:@42170.4]
  assign regs_32_reset = io_reset; // @[:@42171.4 RegFile.scala 76:16:@42178.4]
  assign regs_32_io_in = io_argOuts_30_valid ? io_argOuts_30_bits : io_wdata; // @[RegFile.scala 75:16:@42177.4]
  assign regs_32_io_reset = reset; // @[RegFile.scala 78:19:@42181.4]
  assign regs_32_io_enable = io_argOuts_30_valid | _T_3492; // @[RegFile.scala 74:20:@42175.4]
  assign regs_33_clock = clock; // @[:@42184.4]
  assign regs_33_reset = io_reset; // @[:@42185.4 RegFile.scala 76:16:@42192.4]
  assign regs_33_io_in = io_argOuts_31_valid ? io_argOuts_31_bits : io_wdata; // @[RegFile.scala 75:16:@42191.4]
  assign regs_33_io_reset = reset; // @[RegFile.scala 78:19:@42195.4]
  assign regs_33_io_enable = io_argOuts_31_valid | _T_3499; // @[RegFile.scala 74:20:@42189.4]
  assign regs_34_clock = clock; // @[:@42198.4]
  assign regs_34_reset = io_reset; // @[:@42199.4 RegFile.scala 76:16:@42206.4]
  assign regs_34_io_in = io_argOuts_32_valid ? io_argOuts_32_bits : io_wdata; // @[RegFile.scala 75:16:@42205.4]
  assign regs_34_io_reset = reset; // @[RegFile.scala 78:19:@42209.4]
  assign regs_34_io_enable = io_argOuts_32_valid | _T_3506; // @[RegFile.scala 74:20:@42203.4]
  assign regs_35_clock = clock; // @[:@42212.4]
  assign regs_35_reset = io_reset; // @[:@42213.4 RegFile.scala 76:16:@42220.4]
  assign regs_35_io_in = 64'h0; // @[RegFile.scala 75:16:@42219.4]
  assign regs_35_io_reset = reset; // @[RegFile.scala 78:19:@42223.4]
  assign regs_35_io_enable = 1'h1; // @[RegFile.scala 74:20:@42217.4]
  assign regs_36_clock = clock; // @[:@42226.4]
  assign regs_36_reset = io_reset; // @[:@42227.4 RegFile.scala 76:16:@42234.4]
  assign regs_36_io_in = 64'h0; // @[RegFile.scala 75:16:@42233.4]
  assign regs_36_io_reset = reset; // @[RegFile.scala 78:19:@42237.4]
  assign regs_36_io_enable = 1'h1; // @[RegFile.scala 74:20:@42231.4]
  assign regs_37_clock = clock; // @[:@42240.4]
  assign regs_37_reset = io_reset; // @[:@42241.4 RegFile.scala 76:16:@42248.4]
  assign regs_37_io_in = 64'h0; // @[RegFile.scala 75:16:@42247.4]
  assign regs_37_io_reset = reset; // @[RegFile.scala 78:19:@42251.4]
  assign regs_37_io_enable = 1'h1; // @[RegFile.scala 74:20:@42245.4]
  assign regs_38_clock = clock; // @[:@42254.4]
  assign regs_38_reset = io_reset; // @[:@42255.4 RegFile.scala 76:16:@42262.4]
  assign regs_38_io_in = 64'h0; // @[RegFile.scala 75:16:@42261.4]
  assign regs_38_io_reset = reset; // @[RegFile.scala 78:19:@42265.4]
  assign regs_38_io_enable = 1'h1; // @[RegFile.scala 74:20:@42259.4]
  assign regs_39_clock = clock; // @[:@42268.4]
  assign regs_39_reset = io_reset; // @[:@42269.4 RegFile.scala 76:16:@42276.4]
  assign regs_39_io_in = 64'h0; // @[RegFile.scala 75:16:@42275.4]
  assign regs_39_io_reset = reset; // @[RegFile.scala 78:19:@42279.4]
  assign regs_39_io_enable = 1'h1; // @[RegFile.scala 74:20:@42273.4]
  assign regs_40_clock = clock; // @[:@42282.4]
  assign regs_40_reset = io_reset; // @[:@42283.4 RegFile.scala 76:16:@42290.4]
  assign regs_40_io_in = 64'h0; // @[RegFile.scala 75:16:@42289.4]
  assign regs_40_io_reset = reset; // @[RegFile.scala 78:19:@42293.4]
  assign regs_40_io_enable = 1'h1; // @[RegFile.scala 74:20:@42287.4]
  assign regs_41_clock = clock; // @[:@42296.4]
  assign regs_41_reset = io_reset; // @[:@42297.4 RegFile.scala 76:16:@42304.4]
  assign regs_41_io_in = 64'h0; // @[RegFile.scala 75:16:@42303.4]
  assign regs_41_io_reset = reset; // @[RegFile.scala 78:19:@42307.4]
  assign regs_41_io_enable = 1'h1; // @[RegFile.scala 74:20:@42301.4]
  assign regs_42_clock = clock; // @[:@42310.4]
  assign regs_42_reset = io_reset; // @[:@42311.4 RegFile.scala 76:16:@42318.4]
  assign regs_42_io_in = 64'h0; // @[RegFile.scala 75:16:@42317.4]
  assign regs_42_io_reset = reset; // @[RegFile.scala 78:19:@42321.4]
  assign regs_42_io_enable = 1'h1; // @[RegFile.scala 74:20:@42315.4]
  assign regs_43_clock = clock; // @[:@42324.4]
  assign regs_43_reset = io_reset; // @[:@42325.4 RegFile.scala 76:16:@42332.4]
  assign regs_43_io_in = 64'h0; // @[RegFile.scala 75:16:@42331.4]
  assign regs_43_io_reset = reset; // @[RegFile.scala 78:19:@42335.4]
  assign regs_43_io_enable = 1'h1; // @[RegFile.scala 74:20:@42329.4]
  assign regs_44_clock = clock; // @[:@42338.4]
  assign regs_44_reset = io_reset; // @[:@42339.4 RegFile.scala 76:16:@42346.4]
  assign regs_44_io_in = 64'h0; // @[RegFile.scala 75:16:@42345.4]
  assign regs_44_io_reset = reset; // @[RegFile.scala 78:19:@42349.4]
  assign regs_44_io_enable = 1'h1; // @[RegFile.scala 74:20:@42343.4]
  assign regs_45_clock = clock; // @[:@42352.4]
  assign regs_45_reset = io_reset; // @[:@42353.4 RegFile.scala 76:16:@42360.4]
  assign regs_45_io_in = 64'h0; // @[RegFile.scala 75:16:@42359.4]
  assign regs_45_io_reset = reset; // @[RegFile.scala 78:19:@42363.4]
  assign regs_45_io_enable = 1'h1; // @[RegFile.scala 74:20:@42357.4]
  assign regs_46_clock = clock; // @[:@42366.4]
  assign regs_46_reset = io_reset; // @[:@42367.4 RegFile.scala 76:16:@42374.4]
  assign regs_46_io_in = 64'h0; // @[RegFile.scala 75:16:@42373.4]
  assign regs_46_io_reset = reset; // @[RegFile.scala 78:19:@42377.4]
  assign regs_46_io_enable = 1'h1; // @[RegFile.scala 74:20:@42371.4]
  assign regs_47_clock = clock; // @[:@42380.4]
  assign regs_47_reset = io_reset; // @[:@42381.4 RegFile.scala 76:16:@42388.4]
  assign regs_47_io_in = 64'h0; // @[RegFile.scala 75:16:@42387.4]
  assign regs_47_io_reset = reset; // @[RegFile.scala 78:19:@42391.4]
  assign regs_47_io_enable = 1'h1; // @[RegFile.scala 74:20:@42385.4]
  assign regs_48_clock = clock; // @[:@42394.4]
  assign regs_48_reset = io_reset; // @[:@42395.4 RegFile.scala 76:16:@42402.4]
  assign regs_48_io_in = 64'h0; // @[RegFile.scala 75:16:@42401.4]
  assign regs_48_io_reset = reset; // @[RegFile.scala 78:19:@42405.4]
  assign regs_48_io_enable = 1'h1; // @[RegFile.scala 74:20:@42399.4]
  assign regs_49_clock = clock; // @[:@42408.4]
  assign regs_49_reset = io_reset; // @[:@42409.4 RegFile.scala 76:16:@42416.4]
  assign regs_49_io_in = 64'h0; // @[RegFile.scala 75:16:@42415.4]
  assign regs_49_io_reset = reset; // @[RegFile.scala 78:19:@42419.4]
  assign regs_49_io_enable = 1'h1; // @[RegFile.scala 74:20:@42413.4]
  assign regs_50_clock = clock; // @[:@42422.4]
  assign regs_50_reset = io_reset; // @[:@42423.4 RegFile.scala 76:16:@42430.4]
  assign regs_50_io_in = 64'h0; // @[RegFile.scala 75:16:@42429.4]
  assign regs_50_io_reset = reset; // @[RegFile.scala 78:19:@42433.4]
  assign regs_50_io_enable = 1'h1; // @[RegFile.scala 74:20:@42427.4]
  assign regs_51_clock = clock; // @[:@42436.4]
  assign regs_51_reset = io_reset; // @[:@42437.4 RegFile.scala 76:16:@42444.4]
  assign regs_51_io_in = 64'h0; // @[RegFile.scala 75:16:@42443.4]
  assign regs_51_io_reset = reset; // @[RegFile.scala 78:19:@42447.4]
  assign regs_51_io_enable = 1'h1; // @[RegFile.scala 74:20:@42441.4]
  assign regs_52_clock = clock; // @[:@42450.4]
  assign regs_52_reset = io_reset; // @[:@42451.4 RegFile.scala 76:16:@42458.4]
  assign regs_52_io_in = 64'h0; // @[RegFile.scala 75:16:@42457.4]
  assign regs_52_io_reset = reset; // @[RegFile.scala 78:19:@42461.4]
  assign regs_52_io_enable = 1'h1; // @[RegFile.scala 74:20:@42455.4]
  assign regs_53_clock = clock; // @[:@42464.4]
  assign regs_53_reset = io_reset; // @[:@42465.4 RegFile.scala 76:16:@42472.4]
  assign regs_53_io_in = 64'h0; // @[RegFile.scala 75:16:@42471.4]
  assign regs_53_io_reset = reset; // @[RegFile.scala 78:19:@42475.4]
  assign regs_53_io_enable = 1'h1; // @[RegFile.scala 74:20:@42469.4]
  assign regs_54_clock = clock; // @[:@42478.4]
  assign regs_54_reset = io_reset; // @[:@42479.4 RegFile.scala 76:16:@42486.4]
  assign regs_54_io_in = 64'h0; // @[RegFile.scala 75:16:@42485.4]
  assign regs_54_io_reset = reset; // @[RegFile.scala 78:19:@42489.4]
  assign regs_54_io_enable = 1'h1; // @[RegFile.scala 74:20:@42483.4]
  assign regs_55_clock = clock; // @[:@42492.4]
  assign regs_55_reset = io_reset; // @[:@42493.4 RegFile.scala 76:16:@42500.4]
  assign regs_55_io_in = 64'h0; // @[RegFile.scala 75:16:@42499.4]
  assign regs_55_io_reset = reset; // @[RegFile.scala 78:19:@42503.4]
  assign regs_55_io_enable = 1'h1; // @[RegFile.scala 74:20:@42497.4]
  assign regs_56_clock = clock; // @[:@42506.4]
  assign regs_56_reset = io_reset; // @[:@42507.4 RegFile.scala 76:16:@42514.4]
  assign regs_56_io_in = 64'h0; // @[RegFile.scala 75:16:@42513.4]
  assign regs_56_io_reset = reset; // @[RegFile.scala 78:19:@42517.4]
  assign regs_56_io_enable = 1'h1; // @[RegFile.scala 74:20:@42511.4]
  assign regs_57_clock = clock; // @[:@42520.4]
  assign regs_57_reset = io_reset; // @[:@42521.4 RegFile.scala 76:16:@42528.4]
  assign regs_57_io_in = 64'h0; // @[RegFile.scala 75:16:@42527.4]
  assign regs_57_io_reset = reset; // @[RegFile.scala 78:19:@42531.4]
  assign regs_57_io_enable = 1'h1; // @[RegFile.scala 74:20:@42525.4]
  assign regs_58_clock = clock; // @[:@42534.4]
  assign regs_58_reset = io_reset; // @[:@42535.4 RegFile.scala 76:16:@42542.4]
  assign regs_58_io_in = 64'h0; // @[RegFile.scala 75:16:@42541.4]
  assign regs_58_io_reset = reset; // @[RegFile.scala 78:19:@42545.4]
  assign regs_58_io_enable = 1'h1; // @[RegFile.scala 74:20:@42539.4]
  assign regs_59_clock = clock; // @[:@42548.4]
  assign regs_59_reset = io_reset; // @[:@42549.4 RegFile.scala 76:16:@42556.4]
  assign regs_59_io_in = 64'h0; // @[RegFile.scala 75:16:@42555.4]
  assign regs_59_io_reset = reset; // @[RegFile.scala 78:19:@42559.4]
  assign regs_59_io_enable = 1'h1; // @[RegFile.scala 74:20:@42553.4]
  assign regs_60_clock = clock; // @[:@42562.4]
  assign regs_60_reset = io_reset; // @[:@42563.4 RegFile.scala 76:16:@42570.4]
  assign regs_60_io_in = 64'h0; // @[RegFile.scala 75:16:@42569.4]
  assign regs_60_io_reset = reset; // @[RegFile.scala 78:19:@42573.4]
  assign regs_60_io_enable = 1'h1; // @[RegFile.scala 74:20:@42567.4]
  assign regs_61_clock = clock; // @[:@42576.4]
  assign regs_61_reset = io_reset; // @[:@42577.4 RegFile.scala 76:16:@42584.4]
  assign regs_61_io_in = 64'h0; // @[RegFile.scala 75:16:@42583.4]
  assign regs_61_io_reset = reset; // @[RegFile.scala 78:19:@42587.4]
  assign regs_61_io_enable = 1'h1; // @[RegFile.scala 74:20:@42581.4]
  assign regs_62_clock = clock; // @[:@42590.4]
  assign regs_62_reset = io_reset; // @[:@42591.4 RegFile.scala 76:16:@42598.4]
  assign regs_62_io_in = 64'h0; // @[RegFile.scala 75:16:@42597.4]
  assign regs_62_io_reset = reset; // @[RegFile.scala 78:19:@42601.4]
  assign regs_62_io_enable = 1'h1; // @[RegFile.scala 74:20:@42595.4]
  assign regs_63_clock = clock; // @[:@42604.4]
  assign regs_63_reset = io_reset; // @[:@42605.4 RegFile.scala 76:16:@42612.4]
  assign regs_63_io_in = 64'h0; // @[RegFile.scala 75:16:@42611.4]
  assign regs_63_io_reset = reset; // @[RegFile.scala 78:19:@42615.4]
  assign regs_63_io_enable = 1'h1; // @[RegFile.scala 74:20:@42609.4]
  assign regs_64_clock = clock; // @[:@42618.4]
  assign regs_64_reset = io_reset; // @[:@42619.4 RegFile.scala 76:16:@42626.4]
  assign regs_64_io_in = 64'h0; // @[RegFile.scala 75:16:@42625.4]
  assign regs_64_io_reset = reset; // @[RegFile.scala 78:19:@42629.4]
  assign regs_64_io_enable = 1'h1; // @[RegFile.scala 74:20:@42623.4]
  assign regs_65_clock = clock; // @[:@42632.4]
  assign regs_65_reset = io_reset; // @[:@42633.4 RegFile.scala 76:16:@42640.4]
  assign regs_65_io_in = 64'h0; // @[RegFile.scala 75:16:@42639.4]
  assign regs_65_io_reset = reset; // @[RegFile.scala 78:19:@42643.4]
  assign regs_65_io_enable = 1'h1; // @[RegFile.scala 74:20:@42637.4]
  assign regs_66_clock = clock; // @[:@42646.4]
  assign regs_66_reset = io_reset; // @[:@42647.4 RegFile.scala 76:16:@42654.4]
  assign regs_66_io_in = 64'h0; // @[RegFile.scala 75:16:@42653.4]
  assign regs_66_io_reset = reset; // @[RegFile.scala 78:19:@42657.4]
  assign regs_66_io_enable = 1'h1; // @[RegFile.scala 74:20:@42651.4]
  assign regs_67_clock = clock; // @[:@42660.4]
  assign regs_67_reset = io_reset; // @[:@42661.4 RegFile.scala 76:16:@42668.4]
  assign regs_67_io_in = 64'h0; // @[RegFile.scala 75:16:@42667.4]
  assign regs_67_io_reset = reset; // @[RegFile.scala 78:19:@42671.4]
  assign regs_67_io_enable = 1'h1; // @[RegFile.scala 74:20:@42665.4]
  assign regs_68_clock = clock; // @[:@42674.4]
  assign regs_68_reset = io_reset; // @[:@42675.4 RegFile.scala 76:16:@42682.4]
  assign regs_68_io_in = 64'h0; // @[RegFile.scala 75:16:@42681.4]
  assign regs_68_io_reset = reset; // @[RegFile.scala 78:19:@42685.4]
  assign regs_68_io_enable = 1'h1; // @[RegFile.scala 74:20:@42679.4]
  assign regs_69_clock = clock; // @[:@42688.4]
  assign regs_69_reset = io_reset; // @[:@42689.4 RegFile.scala 76:16:@42696.4]
  assign regs_69_io_in = 64'h0; // @[RegFile.scala 75:16:@42695.4]
  assign regs_69_io_reset = reset; // @[RegFile.scala 78:19:@42699.4]
  assign regs_69_io_enable = 1'h1; // @[RegFile.scala 74:20:@42693.4]
  assign regs_70_clock = clock; // @[:@42702.4]
  assign regs_70_reset = io_reset; // @[:@42703.4 RegFile.scala 76:16:@42710.4]
  assign regs_70_io_in = 64'h0; // @[RegFile.scala 75:16:@42709.4]
  assign regs_70_io_reset = reset; // @[RegFile.scala 78:19:@42713.4]
  assign regs_70_io_enable = 1'h1; // @[RegFile.scala 74:20:@42707.4]
  assign regs_71_clock = clock; // @[:@42716.4]
  assign regs_71_reset = io_reset; // @[:@42717.4 RegFile.scala 76:16:@42724.4]
  assign regs_71_io_in = 64'h0; // @[RegFile.scala 75:16:@42723.4]
  assign regs_71_io_reset = reset; // @[RegFile.scala 78:19:@42727.4]
  assign regs_71_io_enable = 1'h1; // @[RegFile.scala 74:20:@42721.4]
  assign regs_72_clock = clock; // @[:@42730.4]
  assign regs_72_reset = io_reset; // @[:@42731.4 RegFile.scala 76:16:@42738.4]
  assign regs_72_io_in = 64'h0; // @[RegFile.scala 75:16:@42737.4]
  assign regs_72_io_reset = reset; // @[RegFile.scala 78:19:@42741.4]
  assign regs_72_io_enable = 1'h1; // @[RegFile.scala 74:20:@42735.4]
  assign regs_73_clock = clock; // @[:@42744.4]
  assign regs_73_reset = io_reset; // @[:@42745.4 RegFile.scala 76:16:@42752.4]
  assign regs_73_io_in = 64'h0; // @[RegFile.scala 75:16:@42751.4]
  assign regs_73_io_reset = reset; // @[RegFile.scala 78:19:@42755.4]
  assign regs_73_io_enable = 1'h1; // @[RegFile.scala 74:20:@42749.4]
  assign regs_74_clock = clock; // @[:@42758.4]
  assign regs_74_reset = io_reset; // @[:@42759.4 RegFile.scala 76:16:@42766.4]
  assign regs_74_io_in = 64'h0; // @[RegFile.scala 75:16:@42765.4]
  assign regs_74_io_reset = reset; // @[RegFile.scala 78:19:@42769.4]
  assign regs_74_io_enable = 1'h1; // @[RegFile.scala 74:20:@42763.4]
  assign regs_75_clock = clock; // @[:@42772.4]
  assign regs_75_reset = io_reset; // @[:@42773.4 RegFile.scala 76:16:@42780.4]
  assign regs_75_io_in = 64'h0; // @[RegFile.scala 75:16:@42779.4]
  assign regs_75_io_reset = reset; // @[RegFile.scala 78:19:@42783.4]
  assign regs_75_io_enable = 1'h1; // @[RegFile.scala 74:20:@42777.4]
  assign regs_76_clock = clock; // @[:@42786.4]
  assign regs_76_reset = io_reset; // @[:@42787.4 RegFile.scala 76:16:@42794.4]
  assign regs_76_io_in = 64'h0; // @[RegFile.scala 75:16:@42793.4]
  assign regs_76_io_reset = reset; // @[RegFile.scala 78:19:@42797.4]
  assign regs_76_io_enable = 1'h1; // @[RegFile.scala 74:20:@42791.4]
  assign regs_77_clock = clock; // @[:@42800.4]
  assign regs_77_reset = io_reset; // @[:@42801.4 RegFile.scala 76:16:@42808.4]
  assign regs_77_io_in = 64'h0; // @[RegFile.scala 75:16:@42807.4]
  assign regs_77_io_reset = reset; // @[RegFile.scala 78:19:@42811.4]
  assign regs_77_io_enable = 1'h1; // @[RegFile.scala 74:20:@42805.4]
  assign regs_78_clock = clock; // @[:@42814.4]
  assign regs_78_reset = io_reset; // @[:@42815.4 RegFile.scala 76:16:@42822.4]
  assign regs_78_io_in = 64'h0; // @[RegFile.scala 75:16:@42821.4]
  assign regs_78_io_reset = reset; // @[RegFile.scala 78:19:@42825.4]
  assign regs_78_io_enable = 1'h1; // @[RegFile.scala 74:20:@42819.4]
  assign regs_79_clock = clock; // @[:@42828.4]
  assign regs_79_reset = io_reset; // @[:@42829.4 RegFile.scala 76:16:@42836.4]
  assign regs_79_io_in = 64'h0; // @[RegFile.scala 75:16:@42835.4]
  assign regs_79_io_reset = reset; // @[RegFile.scala 78:19:@42839.4]
  assign regs_79_io_enable = 1'h1; // @[RegFile.scala 74:20:@42833.4]
  assign regs_80_clock = clock; // @[:@42842.4]
  assign regs_80_reset = io_reset; // @[:@42843.4 RegFile.scala 76:16:@42850.4]
  assign regs_80_io_in = 64'h0; // @[RegFile.scala 75:16:@42849.4]
  assign regs_80_io_reset = reset; // @[RegFile.scala 78:19:@42853.4]
  assign regs_80_io_enable = 1'h1; // @[RegFile.scala 74:20:@42847.4]
  assign regs_81_clock = clock; // @[:@42856.4]
  assign regs_81_reset = io_reset; // @[:@42857.4 RegFile.scala 76:16:@42864.4]
  assign regs_81_io_in = 64'h0; // @[RegFile.scala 75:16:@42863.4]
  assign regs_81_io_reset = reset; // @[RegFile.scala 78:19:@42867.4]
  assign regs_81_io_enable = 1'h1; // @[RegFile.scala 74:20:@42861.4]
  assign regs_82_clock = clock; // @[:@42870.4]
  assign regs_82_reset = io_reset; // @[:@42871.4 RegFile.scala 76:16:@42878.4]
  assign regs_82_io_in = 64'h0; // @[RegFile.scala 75:16:@42877.4]
  assign regs_82_io_reset = reset; // @[RegFile.scala 78:19:@42881.4]
  assign regs_82_io_enable = 1'h1; // @[RegFile.scala 74:20:@42875.4]
  assign regs_83_clock = clock; // @[:@42884.4]
  assign regs_83_reset = io_reset; // @[:@42885.4 RegFile.scala 76:16:@42892.4]
  assign regs_83_io_in = 64'h0; // @[RegFile.scala 75:16:@42891.4]
  assign regs_83_io_reset = reset; // @[RegFile.scala 78:19:@42895.4]
  assign regs_83_io_enable = 1'h1; // @[RegFile.scala 74:20:@42889.4]
  assign regs_84_clock = clock; // @[:@42898.4]
  assign regs_84_reset = io_reset; // @[:@42899.4 RegFile.scala 76:16:@42906.4]
  assign regs_84_io_in = 64'h0; // @[RegFile.scala 75:16:@42905.4]
  assign regs_84_io_reset = reset; // @[RegFile.scala 78:19:@42909.4]
  assign regs_84_io_enable = 1'h1; // @[RegFile.scala 74:20:@42903.4]
  assign regs_85_clock = clock; // @[:@42912.4]
  assign regs_85_reset = io_reset; // @[:@42913.4 RegFile.scala 76:16:@42920.4]
  assign regs_85_io_in = 64'h0; // @[RegFile.scala 75:16:@42919.4]
  assign regs_85_io_reset = reset; // @[RegFile.scala 78:19:@42923.4]
  assign regs_85_io_enable = 1'h1; // @[RegFile.scala 74:20:@42917.4]
  assign regs_86_clock = clock; // @[:@42926.4]
  assign regs_86_reset = io_reset; // @[:@42927.4 RegFile.scala 76:16:@42934.4]
  assign regs_86_io_in = 64'h0; // @[RegFile.scala 75:16:@42933.4]
  assign regs_86_io_reset = reset; // @[RegFile.scala 78:19:@42937.4]
  assign regs_86_io_enable = 1'h1; // @[RegFile.scala 74:20:@42931.4]
  assign regs_87_clock = clock; // @[:@42940.4]
  assign regs_87_reset = io_reset; // @[:@42941.4 RegFile.scala 76:16:@42948.4]
  assign regs_87_io_in = 64'h0; // @[RegFile.scala 75:16:@42947.4]
  assign regs_87_io_reset = reset; // @[RegFile.scala 78:19:@42951.4]
  assign regs_87_io_enable = 1'h1; // @[RegFile.scala 74:20:@42945.4]
  assign regs_88_clock = clock; // @[:@42954.4]
  assign regs_88_reset = io_reset; // @[:@42955.4 RegFile.scala 76:16:@42962.4]
  assign regs_88_io_in = 64'h0; // @[RegFile.scala 75:16:@42961.4]
  assign regs_88_io_reset = reset; // @[RegFile.scala 78:19:@42965.4]
  assign regs_88_io_enable = 1'h1; // @[RegFile.scala 74:20:@42959.4]
  assign regs_89_clock = clock; // @[:@42968.4]
  assign regs_89_reset = io_reset; // @[:@42969.4 RegFile.scala 76:16:@42976.4]
  assign regs_89_io_in = 64'h0; // @[RegFile.scala 75:16:@42975.4]
  assign regs_89_io_reset = reset; // @[RegFile.scala 78:19:@42979.4]
  assign regs_89_io_enable = 1'h1; // @[RegFile.scala 74:20:@42973.4]
  assign regs_90_clock = clock; // @[:@42982.4]
  assign regs_90_reset = io_reset; // @[:@42983.4 RegFile.scala 76:16:@42990.4]
  assign regs_90_io_in = 64'h0; // @[RegFile.scala 75:16:@42989.4]
  assign regs_90_io_reset = reset; // @[RegFile.scala 78:19:@42993.4]
  assign regs_90_io_enable = 1'h1; // @[RegFile.scala 74:20:@42987.4]
  assign regs_91_clock = clock; // @[:@42996.4]
  assign regs_91_reset = io_reset; // @[:@42997.4 RegFile.scala 76:16:@43004.4]
  assign regs_91_io_in = 64'h0; // @[RegFile.scala 75:16:@43003.4]
  assign regs_91_io_reset = reset; // @[RegFile.scala 78:19:@43007.4]
  assign regs_91_io_enable = 1'h1; // @[RegFile.scala 74:20:@43001.4]
  assign regs_92_clock = clock; // @[:@43010.4]
  assign regs_92_reset = io_reset; // @[:@43011.4 RegFile.scala 76:16:@43018.4]
  assign regs_92_io_in = 64'h0; // @[RegFile.scala 75:16:@43017.4]
  assign regs_92_io_reset = reset; // @[RegFile.scala 78:19:@43021.4]
  assign regs_92_io_enable = 1'h1; // @[RegFile.scala 74:20:@43015.4]
  assign regs_93_clock = clock; // @[:@43024.4]
  assign regs_93_reset = io_reset; // @[:@43025.4 RegFile.scala 76:16:@43032.4]
  assign regs_93_io_in = 64'h0; // @[RegFile.scala 75:16:@43031.4]
  assign regs_93_io_reset = reset; // @[RegFile.scala 78:19:@43035.4]
  assign regs_93_io_enable = 1'h1; // @[RegFile.scala 74:20:@43029.4]
  assign regs_94_clock = clock; // @[:@43038.4]
  assign regs_94_reset = io_reset; // @[:@43039.4 RegFile.scala 76:16:@43046.4]
  assign regs_94_io_in = 64'h0; // @[RegFile.scala 75:16:@43045.4]
  assign regs_94_io_reset = reset; // @[RegFile.scala 78:19:@43049.4]
  assign regs_94_io_enable = 1'h1; // @[RegFile.scala 74:20:@43043.4]
  assign regs_95_clock = clock; // @[:@43052.4]
  assign regs_95_reset = io_reset; // @[:@43053.4 RegFile.scala 76:16:@43060.4]
  assign regs_95_io_in = 64'h0; // @[RegFile.scala 75:16:@43059.4]
  assign regs_95_io_reset = reset; // @[RegFile.scala 78:19:@43063.4]
  assign regs_95_io_enable = 1'h1; // @[RegFile.scala 74:20:@43057.4]
  assign regs_96_clock = clock; // @[:@43066.4]
  assign regs_96_reset = io_reset; // @[:@43067.4 RegFile.scala 76:16:@43074.4]
  assign regs_96_io_in = 64'h0; // @[RegFile.scala 75:16:@43073.4]
  assign regs_96_io_reset = reset; // @[RegFile.scala 78:19:@43077.4]
  assign regs_96_io_enable = 1'h1; // @[RegFile.scala 74:20:@43071.4]
  assign regs_97_clock = clock; // @[:@43080.4]
  assign regs_97_reset = io_reset; // @[:@43081.4 RegFile.scala 76:16:@43088.4]
  assign regs_97_io_in = 64'h0; // @[RegFile.scala 75:16:@43087.4]
  assign regs_97_io_reset = reset; // @[RegFile.scala 78:19:@43091.4]
  assign regs_97_io_enable = 1'h1; // @[RegFile.scala 74:20:@43085.4]
  assign regs_98_clock = clock; // @[:@43094.4]
  assign regs_98_reset = io_reset; // @[:@43095.4 RegFile.scala 76:16:@43102.4]
  assign regs_98_io_in = 64'h0; // @[RegFile.scala 75:16:@43101.4]
  assign regs_98_io_reset = reset; // @[RegFile.scala 78:19:@43105.4]
  assign regs_98_io_enable = 1'h1; // @[RegFile.scala 74:20:@43099.4]
  assign regs_99_clock = clock; // @[:@43108.4]
  assign regs_99_reset = io_reset; // @[:@43109.4 RegFile.scala 76:16:@43116.4]
  assign regs_99_io_in = 64'h0; // @[RegFile.scala 75:16:@43115.4]
  assign regs_99_io_reset = reset; // @[RegFile.scala 78:19:@43119.4]
  assign regs_99_io_enable = 1'h1; // @[RegFile.scala 74:20:@43113.4]
  assign regs_100_clock = clock; // @[:@43122.4]
  assign regs_100_reset = io_reset; // @[:@43123.4 RegFile.scala 76:16:@43130.4]
  assign regs_100_io_in = 64'h0; // @[RegFile.scala 75:16:@43129.4]
  assign regs_100_io_reset = reset; // @[RegFile.scala 78:19:@43133.4]
  assign regs_100_io_enable = 1'h1; // @[RegFile.scala 74:20:@43127.4]
  assign regs_101_clock = clock; // @[:@43136.4]
  assign regs_101_reset = io_reset; // @[:@43137.4 RegFile.scala 76:16:@43144.4]
  assign regs_101_io_in = 64'h0; // @[RegFile.scala 75:16:@43143.4]
  assign regs_101_io_reset = reset; // @[RegFile.scala 78:19:@43147.4]
  assign regs_101_io_enable = 1'h1; // @[RegFile.scala 74:20:@43141.4]
  assign regs_102_clock = clock; // @[:@43150.4]
  assign regs_102_reset = io_reset; // @[:@43151.4 RegFile.scala 76:16:@43158.4]
  assign regs_102_io_in = 64'h0; // @[RegFile.scala 75:16:@43157.4]
  assign regs_102_io_reset = reset; // @[RegFile.scala 78:19:@43161.4]
  assign regs_102_io_enable = 1'h1; // @[RegFile.scala 74:20:@43155.4]
  assign regs_103_clock = clock; // @[:@43164.4]
  assign regs_103_reset = io_reset; // @[:@43165.4 RegFile.scala 76:16:@43172.4]
  assign regs_103_io_in = 64'h0; // @[RegFile.scala 75:16:@43171.4]
  assign regs_103_io_reset = reset; // @[RegFile.scala 78:19:@43175.4]
  assign regs_103_io_enable = 1'h1; // @[RegFile.scala 74:20:@43169.4]
  assign regs_104_clock = clock; // @[:@43178.4]
  assign regs_104_reset = io_reset; // @[:@43179.4 RegFile.scala 76:16:@43186.4]
  assign regs_104_io_in = 64'h0; // @[RegFile.scala 75:16:@43185.4]
  assign regs_104_io_reset = reset; // @[RegFile.scala 78:19:@43189.4]
  assign regs_104_io_enable = 1'h1; // @[RegFile.scala 74:20:@43183.4]
  assign regs_105_clock = clock; // @[:@43192.4]
  assign regs_105_reset = io_reset; // @[:@43193.4 RegFile.scala 76:16:@43200.4]
  assign regs_105_io_in = 64'h0; // @[RegFile.scala 75:16:@43199.4]
  assign regs_105_io_reset = reset; // @[RegFile.scala 78:19:@43203.4]
  assign regs_105_io_enable = 1'h1; // @[RegFile.scala 74:20:@43197.4]
  assign regs_106_clock = clock; // @[:@43206.4]
  assign regs_106_reset = io_reset; // @[:@43207.4 RegFile.scala 76:16:@43214.4]
  assign regs_106_io_in = 64'h0; // @[RegFile.scala 75:16:@43213.4]
  assign regs_106_io_reset = reset; // @[RegFile.scala 78:19:@43217.4]
  assign regs_106_io_enable = 1'h1; // @[RegFile.scala 74:20:@43211.4]
  assign regs_107_clock = clock; // @[:@43220.4]
  assign regs_107_reset = io_reset; // @[:@43221.4 RegFile.scala 76:16:@43228.4]
  assign regs_107_io_in = 64'h0; // @[RegFile.scala 75:16:@43227.4]
  assign regs_107_io_reset = reset; // @[RegFile.scala 78:19:@43231.4]
  assign regs_107_io_enable = 1'h1; // @[RegFile.scala 74:20:@43225.4]
  assign regs_108_clock = clock; // @[:@43234.4]
  assign regs_108_reset = io_reset; // @[:@43235.4 RegFile.scala 76:16:@43242.4]
  assign regs_108_io_in = 64'h0; // @[RegFile.scala 75:16:@43241.4]
  assign regs_108_io_reset = reset; // @[RegFile.scala 78:19:@43245.4]
  assign regs_108_io_enable = 1'h1; // @[RegFile.scala 74:20:@43239.4]
  assign regs_109_clock = clock; // @[:@43248.4]
  assign regs_109_reset = io_reset; // @[:@43249.4 RegFile.scala 76:16:@43256.4]
  assign regs_109_io_in = 64'h0; // @[RegFile.scala 75:16:@43255.4]
  assign regs_109_io_reset = reset; // @[RegFile.scala 78:19:@43259.4]
  assign regs_109_io_enable = 1'h1; // @[RegFile.scala 74:20:@43253.4]
  assign regs_110_clock = clock; // @[:@43262.4]
  assign regs_110_reset = io_reset; // @[:@43263.4 RegFile.scala 76:16:@43270.4]
  assign regs_110_io_in = 64'h0; // @[RegFile.scala 75:16:@43269.4]
  assign regs_110_io_reset = reset; // @[RegFile.scala 78:19:@43273.4]
  assign regs_110_io_enable = 1'h1; // @[RegFile.scala 74:20:@43267.4]
  assign regs_111_clock = clock; // @[:@43276.4]
  assign regs_111_reset = io_reset; // @[:@43277.4 RegFile.scala 76:16:@43284.4]
  assign regs_111_io_in = 64'h0; // @[RegFile.scala 75:16:@43283.4]
  assign regs_111_io_reset = reset; // @[RegFile.scala 78:19:@43287.4]
  assign regs_111_io_enable = 1'h1; // @[RegFile.scala 74:20:@43281.4]
  assign regs_112_clock = clock; // @[:@43290.4]
  assign regs_112_reset = io_reset; // @[:@43291.4 RegFile.scala 76:16:@43298.4]
  assign regs_112_io_in = 64'h0; // @[RegFile.scala 75:16:@43297.4]
  assign regs_112_io_reset = reset; // @[RegFile.scala 78:19:@43301.4]
  assign regs_112_io_enable = 1'h1; // @[RegFile.scala 74:20:@43295.4]
  assign regs_113_clock = clock; // @[:@43304.4]
  assign regs_113_reset = io_reset; // @[:@43305.4 RegFile.scala 76:16:@43312.4]
  assign regs_113_io_in = 64'h0; // @[RegFile.scala 75:16:@43311.4]
  assign regs_113_io_reset = reset; // @[RegFile.scala 78:19:@43315.4]
  assign regs_113_io_enable = 1'h1; // @[RegFile.scala 74:20:@43309.4]
  assign regs_114_clock = clock; // @[:@43318.4]
  assign regs_114_reset = io_reset; // @[:@43319.4 RegFile.scala 76:16:@43326.4]
  assign regs_114_io_in = 64'h0; // @[RegFile.scala 75:16:@43325.4]
  assign regs_114_io_reset = reset; // @[RegFile.scala 78:19:@43329.4]
  assign regs_114_io_enable = 1'h1; // @[RegFile.scala 74:20:@43323.4]
  assign regs_115_clock = clock; // @[:@43332.4]
  assign regs_115_reset = io_reset; // @[:@43333.4 RegFile.scala 76:16:@43340.4]
  assign regs_115_io_in = 64'h0; // @[RegFile.scala 75:16:@43339.4]
  assign regs_115_io_reset = reset; // @[RegFile.scala 78:19:@43343.4]
  assign regs_115_io_enable = 1'h1; // @[RegFile.scala 74:20:@43337.4]
  assign regs_116_clock = clock; // @[:@43346.4]
  assign regs_116_reset = io_reset; // @[:@43347.4 RegFile.scala 76:16:@43354.4]
  assign regs_116_io_in = 64'h0; // @[RegFile.scala 75:16:@43353.4]
  assign regs_116_io_reset = reset; // @[RegFile.scala 78:19:@43357.4]
  assign regs_116_io_enable = 1'h1; // @[RegFile.scala 74:20:@43351.4]
  assign regs_117_clock = clock; // @[:@43360.4]
  assign regs_117_reset = io_reset; // @[:@43361.4 RegFile.scala 76:16:@43368.4]
  assign regs_117_io_in = 64'h0; // @[RegFile.scala 75:16:@43367.4]
  assign regs_117_io_reset = reset; // @[RegFile.scala 78:19:@43371.4]
  assign regs_117_io_enable = 1'h1; // @[RegFile.scala 74:20:@43365.4]
  assign regs_118_clock = clock; // @[:@43374.4]
  assign regs_118_reset = io_reset; // @[:@43375.4 RegFile.scala 76:16:@43382.4]
  assign regs_118_io_in = 64'h0; // @[RegFile.scala 75:16:@43381.4]
  assign regs_118_io_reset = reset; // @[RegFile.scala 78:19:@43385.4]
  assign regs_118_io_enable = 1'h1; // @[RegFile.scala 74:20:@43379.4]
  assign regs_119_clock = clock; // @[:@43388.4]
  assign regs_119_reset = io_reset; // @[:@43389.4 RegFile.scala 76:16:@43396.4]
  assign regs_119_io_in = 64'h0; // @[RegFile.scala 75:16:@43395.4]
  assign regs_119_io_reset = reset; // @[RegFile.scala 78:19:@43399.4]
  assign regs_119_io_enable = 1'h1; // @[RegFile.scala 74:20:@43393.4]
  assign regs_120_clock = clock; // @[:@43402.4]
  assign regs_120_reset = io_reset; // @[:@43403.4 RegFile.scala 76:16:@43410.4]
  assign regs_120_io_in = 64'h0; // @[RegFile.scala 75:16:@43409.4]
  assign regs_120_io_reset = reset; // @[RegFile.scala 78:19:@43413.4]
  assign regs_120_io_enable = 1'h1; // @[RegFile.scala 74:20:@43407.4]
  assign regs_121_clock = clock; // @[:@43416.4]
  assign regs_121_reset = io_reset; // @[:@43417.4 RegFile.scala 76:16:@43424.4]
  assign regs_121_io_in = 64'h0; // @[RegFile.scala 75:16:@43423.4]
  assign regs_121_io_reset = reset; // @[RegFile.scala 78:19:@43427.4]
  assign regs_121_io_enable = 1'h1; // @[RegFile.scala 74:20:@43421.4]
  assign regs_122_clock = clock; // @[:@43430.4]
  assign regs_122_reset = io_reset; // @[:@43431.4 RegFile.scala 76:16:@43438.4]
  assign regs_122_io_in = 64'h0; // @[RegFile.scala 75:16:@43437.4]
  assign regs_122_io_reset = reset; // @[RegFile.scala 78:19:@43441.4]
  assign regs_122_io_enable = 1'h1; // @[RegFile.scala 74:20:@43435.4]
  assign regs_123_clock = clock; // @[:@43444.4]
  assign regs_123_reset = io_reset; // @[:@43445.4 RegFile.scala 76:16:@43452.4]
  assign regs_123_io_in = 64'h0; // @[RegFile.scala 75:16:@43451.4]
  assign regs_123_io_reset = reset; // @[RegFile.scala 78:19:@43455.4]
  assign regs_123_io_enable = 1'h1; // @[RegFile.scala 74:20:@43449.4]
  assign regs_124_clock = clock; // @[:@43458.4]
  assign regs_124_reset = io_reset; // @[:@43459.4 RegFile.scala 76:16:@43466.4]
  assign regs_124_io_in = 64'h0; // @[RegFile.scala 75:16:@43465.4]
  assign regs_124_io_reset = reset; // @[RegFile.scala 78:19:@43469.4]
  assign regs_124_io_enable = 1'h1; // @[RegFile.scala 74:20:@43463.4]
  assign regs_125_clock = clock; // @[:@43472.4]
  assign regs_125_reset = io_reset; // @[:@43473.4 RegFile.scala 76:16:@43480.4]
  assign regs_125_io_in = 64'h0; // @[RegFile.scala 75:16:@43479.4]
  assign regs_125_io_reset = reset; // @[RegFile.scala 78:19:@43483.4]
  assign regs_125_io_enable = 1'h1; // @[RegFile.scala 74:20:@43477.4]
  assign regs_126_clock = clock; // @[:@43486.4]
  assign regs_126_reset = io_reset; // @[:@43487.4 RegFile.scala 76:16:@43494.4]
  assign regs_126_io_in = 64'h0; // @[RegFile.scala 75:16:@43493.4]
  assign regs_126_io_reset = reset; // @[RegFile.scala 78:19:@43497.4]
  assign regs_126_io_enable = 1'h1; // @[RegFile.scala 74:20:@43491.4]
  assign regs_127_clock = clock; // @[:@43500.4]
  assign regs_127_reset = io_reset; // @[:@43501.4 RegFile.scala 76:16:@43508.4]
  assign regs_127_io_in = 64'h0; // @[RegFile.scala 75:16:@43507.4]
  assign regs_127_io_reset = reset; // @[RegFile.scala 78:19:@43511.4]
  assign regs_127_io_enable = 1'h1; // @[RegFile.scala 74:20:@43505.4]
  assign regs_128_clock = clock; // @[:@43514.4]
  assign regs_128_reset = io_reset; // @[:@43515.4 RegFile.scala 76:16:@43522.4]
  assign regs_128_io_in = 64'h0; // @[RegFile.scala 75:16:@43521.4]
  assign regs_128_io_reset = reset; // @[RegFile.scala 78:19:@43525.4]
  assign regs_128_io_enable = 1'h1; // @[RegFile.scala 74:20:@43519.4]
  assign regs_129_clock = clock; // @[:@43528.4]
  assign regs_129_reset = io_reset; // @[:@43529.4 RegFile.scala 76:16:@43536.4]
  assign regs_129_io_in = 64'h0; // @[RegFile.scala 75:16:@43535.4]
  assign regs_129_io_reset = reset; // @[RegFile.scala 78:19:@43539.4]
  assign regs_129_io_enable = 1'h1; // @[RegFile.scala 74:20:@43533.4]
  assign regs_130_clock = clock; // @[:@43542.4]
  assign regs_130_reset = io_reset; // @[:@43543.4 RegFile.scala 76:16:@43550.4]
  assign regs_130_io_in = 64'h0; // @[RegFile.scala 75:16:@43549.4]
  assign regs_130_io_reset = reset; // @[RegFile.scala 78:19:@43553.4]
  assign regs_130_io_enable = 1'h1; // @[RegFile.scala 74:20:@43547.4]
  assign regs_131_clock = clock; // @[:@43556.4]
  assign regs_131_reset = io_reset; // @[:@43557.4 RegFile.scala 76:16:@43564.4]
  assign regs_131_io_in = 64'h0; // @[RegFile.scala 75:16:@43563.4]
  assign regs_131_io_reset = reset; // @[RegFile.scala 78:19:@43567.4]
  assign regs_131_io_enable = 1'h1; // @[RegFile.scala 74:20:@43561.4]
  assign regs_132_clock = clock; // @[:@43570.4]
  assign regs_132_reset = io_reset; // @[:@43571.4 RegFile.scala 76:16:@43578.4]
  assign regs_132_io_in = 64'h0; // @[RegFile.scala 75:16:@43577.4]
  assign regs_132_io_reset = reset; // @[RegFile.scala 78:19:@43581.4]
  assign regs_132_io_enable = 1'h1; // @[RegFile.scala 74:20:@43575.4]
  assign regs_133_clock = clock; // @[:@43584.4]
  assign regs_133_reset = io_reset; // @[:@43585.4 RegFile.scala 76:16:@43592.4]
  assign regs_133_io_in = 64'h0; // @[RegFile.scala 75:16:@43591.4]
  assign regs_133_io_reset = reset; // @[RegFile.scala 78:19:@43595.4]
  assign regs_133_io_enable = 1'h1; // @[RegFile.scala 74:20:@43589.4]
  assign regs_134_clock = clock; // @[:@43598.4]
  assign regs_134_reset = io_reset; // @[:@43599.4 RegFile.scala 76:16:@43606.4]
  assign regs_134_io_in = 64'h0; // @[RegFile.scala 75:16:@43605.4]
  assign regs_134_io_reset = reset; // @[RegFile.scala 78:19:@43609.4]
  assign regs_134_io_enable = 1'h1; // @[RegFile.scala 74:20:@43603.4]
  assign regs_135_clock = clock; // @[:@43612.4]
  assign regs_135_reset = io_reset; // @[:@43613.4 RegFile.scala 76:16:@43620.4]
  assign regs_135_io_in = 64'h0; // @[RegFile.scala 75:16:@43619.4]
  assign regs_135_io_reset = reset; // @[RegFile.scala 78:19:@43623.4]
  assign regs_135_io_enable = 1'h1; // @[RegFile.scala 74:20:@43617.4]
  assign regs_136_clock = clock; // @[:@43626.4]
  assign regs_136_reset = io_reset; // @[:@43627.4 RegFile.scala 76:16:@43634.4]
  assign regs_136_io_in = 64'h0; // @[RegFile.scala 75:16:@43633.4]
  assign regs_136_io_reset = reset; // @[RegFile.scala 78:19:@43637.4]
  assign regs_136_io_enable = 1'h1; // @[RegFile.scala 74:20:@43631.4]
  assign regs_137_clock = clock; // @[:@43640.4]
  assign regs_137_reset = io_reset; // @[:@43641.4 RegFile.scala 76:16:@43648.4]
  assign regs_137_io_in = 64'h0; // @[RegFile.scala 75:16:@43647.4]
  assign regs_137_io_reset = reset; // @[RegFile.scala 78:19:@43651.4]
  assign regs_137_io_enable = 1'h1; // @[RegFile.scala 74:20:@43645.4]
  assign regs_138_clock = clock; // @[:@43654.4]
  assign regs_138_reset = io_reset; // @[:@43655.4 RegFile.scala 76:16:@43662.4]
  assign regs_138_io_in = 64'h0; // @[RegFile.scala 75:16:@43661.4]
  assign regs_138_io_reset = reset; // @[RegFile.scala 78:19:@43665.4]
  assign regs_138_io_enable = 1'h1; // @[RegFile.scala 74:20:@43659.4]
  assign regs_139_clock = clock; // @[:@43668.4]
  assign regs_139_reset = io_reset; // @[:@43669.4 RegFile.scala 76:16:@43676.4]
  assign regs_139_io_in = 64'h0; // @[RegFile.scala 75:16:@43675.4]
  assign regs_139_io_reset = reset; // @[RegFile.scala 78:19:@43679.4]
  assign regs_139_io_enable = 1'h1; // @[RegFile.scala 74:20:@43673.4]
  assign regs_140_clock = clock; // @[:@43682.4]
  assign regs_140_reset = io_reset; // @[:@43683.4 RegFile.scala 76:16:@43690.4]
  assign regs_140_io_in = 64'h0; // @[RegFile.scala 75:16:@43689.4]
  assign regs_140_io_reset = reset; // @[RegFile.scala 78:19:@43693.4]
  assign regs_140_io_enable = 1'h1; // @[RegFile.scala 74:20:@43687.4]
  assign regs_141_clock = clock; // @[:@43696.4]
  assign regs_141_reset = io_reset; // @[:@43697.4 RegFile.scala 76:16:@43704.4]
  assign regs_141_io_in = 64'h0; // @[RegFile.scala 75:16:@43703.4]
  assign regs_141_io_reset = reset; // @[RegFile.scala 78:19:@43707.4]
  assign regs_141_io_enable = 1'h1; // @[RegFile.scala 74:20:@43701.4]
  assign regs_142_clock = clock; // @[:@43710.4]
  assign regs_142_reset = io_reset; // @[:@43711.4 RegFile.scala 76:16:@43718.4]
  assign regs_142_io_in = 64'h0; // @[RegFile.scala 75:16:@43717.4]
  assign regs_142_io_reset = reset; // @[RegFile.scala 78:19:@43721.4]
  assign regs_142_io_enable = 1'h1; // @[RegFile.scala 74:20:@43715.4]
  assign regs_143_clock = clock; // @[:@43724.4]
  assign regs_143_reset = io_reset; // @[:@43725.4 RegFile.scala 76:16:@43732.4]
  assign regs_143_io_in = 64'h0; // @[RegFile.scala 75:16:@43731.4]
  assign regs_143_io_reset = reset; // @[RegFile.scala 78:19:@43735.4]
  assign regs_143_io_enable = 1'h1; // @[RegFile.scala 74:20:@43729.4]
  assign regs_144_clock = clock; // @[:@43738.4]
  assign regs_144_reset = io_reset; // @[:@43739.4 RegFile.scala 76:16:@43746.4]
  assign regs_144_io_in = 64'h0; // @[RegFile.scala 75:16:@43745.4]
  assign regs_144_io_reset = reset; // @[RegFile.scala 78:19:@43749.4]
  assign regs_144_io_enable = 1'h1; // @[RegFile.scala 74:20:@43743.4]
  assign regs_145_clock = clock; // @[:@43752.4]
  assign regs_145_reset = io_reset; // @[:@43753.4 RegFile.scala 76:16:@43760.4]
  assign regs_145_io_in = 64'h0; // @[RegFile.scala 75:16:@43759.4]
  assign regs_145_io_reset = reset; // @[RegFile.scala 78:19:@43763.4]
  assign regs_145_io_enable = 1'h1; // @[RegFile.scala 74:20:@43757.4]
  assign regs_146_clock = clock; // @[:@43766.4]
  assign regs_146_reset = io_reset; // @[:@43767.4 RegFile.scala 76:16:@43774.4]
  assign regs_146_io_in = 64'h0; // @[RegFile.scala 75:16:@43773.4]
  assign regs_146_io_reset = reset; // @[RegFile.scala 78:19:@43777.4]
  assign regs_146_io_enable = 1'h1; // @[RegFile.scala 74:20:@43771.4]
  assign regs_147_clock = clock; // @[:@43780.4]
  assign regs_147_reset = io_reset; // @[:@43781.4 RegFile.scala 76:16:@43788.4]
  assign regs_147_io_in = 64'h0; // @[RegFile.scala 75:16:@43787.4]
  assign regs_147_io_reset = reset; // @[RegFile.scala 78:19:@43791.4]
  assign regs_147_io_enable = 1'h1; // @[RegFile.scala 74:20:@43785.4]
  assign regs_148_clock = clock; // @[:@43794.4]
  assign regs_148_reset = io_reset; // @[:@43795.4 RegFile.scala 76:16:@43802.4]
  assign regs_148_io_in = 64'h0; // @[RegFile.scala 75:16:@43801.4]
  assign regs_148_io_reset = reset; // @[RegFile.scala 78:19:@43805.4]
  assign regs_148_io_enable = 1'h1; // @[RegFile.scala 74:20:@43799.4]
  assign regs_149_clock = clock; // @[:@43808.4]
  assign regs_149_reset = io_reset; // @[:@43809.4 RegFile.scala 76:16:@43816.4]
  assign regs_149_io_in = 64'h0; // @[RegFile.scala 75:16:@43815.4]
  assign regs_149_io_reset = reset; // @[RegFile.scala 78:19:@43819.4]
  assign regs_149_io_enable = 1'h1; // @[RegFile.scala 74:20:@43813.4]
  assign regs_150_clock = clock; // @[:@43822.4]
  assign regs_150_reset = io_reset; // @[:@43823.4 RegFile.scala 76:16:@43830.4]
  assign regs_150_io_in = 64'h0; // @[RegFile.scala 75:16:@43829.4]
  assign regs_150_io_reset = reset; // @[RegFile.scala 78:19:@43833.4]
  assign regs_150_io_enable = 1'h1; // @[RegFile.scala 74:20:@43827.4]
  assign regs_151_clock = clock; // @[:@43836.4]
  assign regs_151_reset = io_reset; // @[:@43837.4 RegFile.scala 76:16:@43844.4]
  assign regs_151_io_in = 64'h0; // @[RegFile.scala 75:16:@43843.4]
  assign regs_151_io_reset = reset; // @[RegFile.scala 78:19:@43847.4]
  assign regs_151_io_enable = 1'h1; // @[RegFile.scala 74:20:@43841.4]
  assign regs_152_clock = clock; // @[:@43850.4]
  assign regs_152_reset = io_reset; // @[:@43851.4 RegFile.scala 76:16:@43858.4]
  assign regs_152_io_in = 64'h0; // @[RegFile.scala 75:16:@43857.4]
  assign regs_152_io_reset = reset; // @[RegFile.scala 78:19:@43861.4]
  assign regs_152_io_enable = 1'h1; // @[RegFile.scala 74:20:@43855.4]
  assign regs_153_clock = clock; // @[:@43864.4]
  assign regs_153_reset = io_reset; // @[:@43865.4 RegFile.scala 76:16:@43872.4]
  assign regs_153_io_in = 64'h0; // @[RegFile.scala 75:16:@43871.4]
  assign regs_153_io_reset = reset; // @[RegFile.scala 78:19:@43875.4]
  assign regs_153_io_enable = 1'h1; // @[RegFile.scala 74:20:@43869.4]
  assign regs_154_clock = clock; // @[:@43878.4]
  assign regs_154_reset = io_reset; // @[:@43879.4 RegFile.scala 76:16:@43886.4]
  assign regs_154_io_in = 64'h0; // @[RegFile.scala 75:16:@43885.4]
  assign regs_154_io_reset = reset; // @[RegFile.scala 78:19:@43889.4]
  assign regs_154_io_enable = 1'h1; // @[RegFile.scala 74:20:@43883.4]
  assign regs_155_clock = clock; // @[:@43892.4]
  assign regs_155_reset = io_reset; // @[:@43893.4 RegFile.scala 76:16:@43900.4]
  assign regs_155_io_in = 64'h0; // @[RegFile.scala 75:16:@43899.4]
  assign regs_155_io_reset = reset; // @[RegFile.scala 78:19:@43903.4]
  assign regs_155_io_enable = 1'h1; // @[RegFile.scala 74:20:@43897.4]
  assign regs_156_clock = clock; // @[:@43906.4]
  assign regs_156_reset = io_reset; // @[:@43907.4 RegFile.scala 76:16:@43914.4]
  assign regs_156_io_in = 64'h0; // @[RegFile.scala 75:16:@43913.4]
  assign regs_156_io_reset = reset; // @[RegFile.scala 78:19:@43917.4]
  assign regs_156_io_enable = 1'h1; // @[RegFile.scala 74:20:@43911.4]
  assign regs_157_clock = clock; // @[:@43920.4]
  assign regs_157_reset = io_reset; // @[:@43921.4 RegFile.scala 76:16:@43928.4]
  assign regs_157_io_in = 64'h0; // @[RegFile.scala 75:16:@43927.4]
  assign regs_157_io_reset = reset; // @[RegFile.scala 78:19:@43931.4]
  assign regs_157_io_enable = 1'h1; // @[RegFile.scala 74:20:@43925.4]
  assign regs_158_clock = clock; // @[:@43934.4]
  assign regs_158_reset = io_reset; // @[:@43935.4 RegFile.scala 76:16:@43942.4]
  assign regs_158_io_in = 64'h0; // @[RegFile.scala 75:16:@43941.4]
  assign regs_158_io_reset = reset; // @[RegFile.scala 78:19:@43945.4]
  assign regs_158_io_enable = 1'h1; // @[RegFile.scala 74:20:@43939.4]
  assign regs_159_clock = clock; // @[:@43948.4]
  assign regs_159_reset = io_reset; // @[:@43949.4 RegFile.scala 76:16:@43956.4]
  assign regs_159_io_in = 64'h0; // @[RegFile.scala 75:16:@43955.4]
  assign regs_159_io_reset = reset; // @[RegFile.scala 78:19:@43959.4]
  assign regs_159_io_enable = 1'h1; // @[RegFile.scala 74:20:@43953.4]
  assign regs_160_clock = clock; // @[:@43962.4]
  assign regs_160_reset = io_reset; // @[:@43963.4 RegFile.scala 76:16:@43970.4]
  assign regs_160_io_in = 64'h0; // @[RegFile.scala 75:16:@43969.4]
  assign regs_160_io_reset = reset; // @[RegFile.scala 78:19:@43973.4]
  assign regs_160_io_enable = 1'h1; // @[RegFile.scala 74:20:@43967.4]
  assign regs_161_clock = clock; // @[:@43976.4]
  assign regs_161_reset = io_reset; // @[:@43977.4 RegFile.scala 76:16:@43984.4]
  assign regs_161_io_in = 64'h0; // @[RegFile.scala 75:16:@43983.4]
  assign regs_161_io_reset = reset; // @[RegFile.scala 78:19:@43987.4]
  assign regs_161_io_enable = 1'h1; // @[RegFile.scala 74:20:@43981.4]
  assign regs_162_clock = clock; // @[:@43990.4]
  assign regs_162_reset = io_reset; // @[:@43991.4 RegFile.scala 76:16:@43998.4]
  assign regs_162_io_in = 64'h0; // @[RegFile.scala 75:16:@43997.4]
  assign regs_162_io_reset = reset; // @[RegFile.scala 78:19:@44001.4]
  assign regs_162_io_enable = 1'h1; // @[RegFile.scala 74:20:@43995.4]
  assign regs_163_clock = clock; // @[:@44004.4]
  assign regs_163_reset = io_reset; // @[:@44005.4 RegFile.scala 76:16:@44012.4]
  assign regs_163_io_in = 64'h0; // @[RegFile.scala 75:16:@44011.4]
  assign regs_163_io_reset = reset; // @[RegFile.scala 78:19:@44015.4]
  assign regs_163_io_enable = 1'h1; // @[RegFile.scala 74:20:@44009.4]
  assign regs_164_clock = clock; // @[:@44018.4]
  assign regs_164_reset = io_reset; // @[:@44019.4 RegFile.scala 76:16:@44026.4]
  assign regs_164_io_in = 64'h0; // @[RegFile.scala 75:16:@44025.4]
  assign regs_164_io_reset = reset; // @[RegFile.scala 78:19:@44029.4]
  assign regs_164_io_enable = 1'h1; // @[RegFile.scala 74:20:@44023.4]
  assign regs_165_clock = clock; // @[:@44032.4]
  assign regs_165_reset = io_reset; // @[:@44033.4 RegFile.scala 76:16:@44040.4]
  assign regs_165_io_in = 64'h0; // @[RegFile.scala 75:16:@44039.4]
  assign regs_165_io_reset = reset; // @[RegFile.scala 78:19:@44043.4]
  assign regs_165_io_enable = 1'h1; // @[RegFile.scala 74:20:@44037.4]
  assign regs_166_clock = clock; // @[:@44046.4]
  assign regs_166_reset = io_reset; // @[:@44047.4 RegFile.scala 76:16:@44054.4]
  assign regs_166_io_in = 64'h0; // @[RegFile.scala 75:16:@44053.4]
  assign regs_166_io_reset = reset; // @[RegFile.scala 78:19:@44057.4]
  assign regs_166_io_enable = 1'h1; // @[RegFile.scala 74:20:@44051.4]
  assign regs_167_clock = clock; // @[:@44060.4]
  assign regs_167_reset = io_reset; // @[:@44061.4 RegFile.scala 76:16:@44068.4]
  assign regs_167_io_in = 64'h0; // @[RegFile.scala 75:16:@44067.4]
  assign regs_167_io_reset = reset; // @[RegFile.scala 78:19:@44071.4]
  assign regs_167_io_enable = 1'h1; // @[RegFile.scala 74:20:@44065.4]
  assign regs_168_clock = clock; // @[:@44074.4]
  assign regs_168_reset = io_reset; // @[:@44075.4 RegFile.scala 76:16:@44082.4]
  assign regs_168_io_in = 64'h0; // @[RegFile.scala 75:16:@44081.4]
  assign regs_168_io_reset = reset; // @[RegFile.scala 78:19:@44085.4]
  assign regs_168_io_enable = 1'h1; // @[RegFile.scala 74:20:@44079.4]
  assign regs_169_clock = clock; // @[:@44088.4]
  assign regs_169_reset = io_reset; // @[:@44089.4 RegFile.scala 76:16:@44096.4]
  assign regs_169_io_in = 64'h0; // @[RegFile.scala 75:16:@44095.4]
  assign regs_169_io_reset = reset; // @[RegFile.scala 78:19:@44099.4]
  assign regs_169_io_enable = 1'h1; // @[RegFile.scala 74:20:@44093.4]
  assign regs_170_clock = clock; // @[:@44102.4]
  assign regs_170_reset = io_reset; // @[:@44103.4 RegFile.scala 76:16:@44110.4]
  assign regs_170_io_in = 64'h0; // @[RegFile.scala 75:16:@44109.4]
  assign regs_170_io_reset = reset; // @[RegFile.scala 78:19:@44113.4]
  assign regs_170_io_enable = 1'h1; // @[RegFile.scala 74:20:@44107.4]
  assign regs_171_clock = clock; // @[:@44116.4]
  assign regs_171_reset = io_reset; // @[:@44117.4 RegFile.scala 76:16:@44124.4]
  assign regs_171_io_in = 64'h0; // @[RegFile.scala 75:16:@44123.4]
  assign regs_171_io_reset = reset; // @[RegFile.scala 78:19:@44127.4]
  assign regs_171_io_enable = 1'h1; // @[RegFile.scala 74:20:@44121.4]
  assign regs_172_clock = clock; // @[:@44130.4]
  assign regs_172_reset = io_reset; // @[:@44131.4 RegFile.scala 76:16:@44138.4]
  assign regs_172_io_in = 64'h0; // @[RegFile.scala 75:16:@44137.4]
  assign regs_172_io_reset = reset; // @[RegFile.scala 78:19:@44141.4]
  assign regs_172_io_enable = 1'h1; // @[RegFile.scala 74:20:@44135.4]
  assign regs_173_clock = clock; // @[:@44144.4]
  assign regs_173_reset = io_reset; // @[:@44145.4 RegFile.scala 76:16:@44152.4]
  assign regs_173_io_in = 64'h0; // @[RegFile.scala 75:16:@44151.4]
  assign regs_173_io_reset = reset; // @[RegFile.scala 78:19:@44155.4]
  assign regs_173_io_enable = 1'h1; // @[RegFile.scala 74:20:@44149.4]
  assign regs_174_clock = clock; // @[:@44158.4]
  assign regs_174_reset = io_reset; // @[:@44159.4 RegFile.scala 76:16:@44166.4]
  assign regs_174_io_in = 64'h0; // @[RegFile.scala 75:16:@44165.4]
  assign regs_174_io_reset = reset; // @[RegFile.scala 78:19:@44169.4]
  assign regs_174_io_enable = 1'h1; // @[RegFile.scala 74:20:@44163.4]
  assign regs_175_clock = clock; // @[:@44172.4]
  assign regs_175_reset = io_reset; // @[:@44173.4 RegFile.scala 76:16:@44180.4]
  assign regs_175_io_in = 64'h0; // @[RegFile.scala 75:16:@44179.4]
  assign regs_175_io_reset = reset; // @[RegFile.scala 78:19:@44183.4]
  assign regs_175_io_enable = 1'h1; // @[RegFile.scala 74:20:@44177.4]
  assign regs_176_clock = clock; // @[:@44186.4]
  assign regs_176_reset = io_reset; // @[:@44187.4 RegFile.scala 76:16:@44194.4]
  assign regs_176_io_in = 64'h0; // @[RegFile.scala 75:16:@44193.4]
  assign regs_176_io_reset = reset; // @[RegFile.scala 78:19:@44197.4]
  assign regs_176_io_enable = 1'h1; // @[RegFile.scala 74:20:@44191.4]
  assign regs_177_clock = clock; // @[:@44200.4]
  assign regs_177_reset = io_reset; // @[:@44201.4 RegFile.scala 76:16:@44208.4]
  assign regs_177_io_in = 64'h0; // @[RegFile.scala 75:16:@44207.4]
  assign regs_177_io_reset = reset; // @[RegFile.scala 78:19:@44211.4]
  assign regs_177_io_enable = 1'h1; // @[RegFile.scala 74:20:@44205.4]
  assign regs_178_clock = clock; // @[:@44214.4]
  assign regs_178_reset = io_reset; // @[:@44215.4 RegFile.scala 76:16:@44222.4]
  assign regs_178_io_in = 64'h0; // @[RegFile.scala 75:16:@44221.4]
  assign regs_178_io_reset = reset; // @[RegFile.scala 78:19:@44225.4]
  assign regs_178_io_enable = 1'h1; // @[RegFile.scala 74:20:@44219.4]
  assign regs_179_clock = clock; // @[:@44228.4]
  assign regs_179_reset = io_reset; // @[:@44229.4 RegFile.scala 76:16:@44236.4]
  assign regs_179_io_in = 64'h0; // @[RegFile.scala 75:16:@44235.4]
  assign regs_179_io_reset = reset; // @[RegFile.scala 78:19:@44239.4]
  assign regs_179_io_enable = 1'h1; // @[RegFile.scala 74:20:@44233.4]
  assign regs_180_clock = clock; // @[:@44242.4]
  assign regs_180_reset = io_reset; // @[:@44243.4 RegFile.scala 76:16:@44250.4]
  assign regs_180_io_in = 64'h0; // @[RegFile.scala 75:16:@44249.4]
  assign regs_180_io_reset = reset; // @[RegFile.scala 78:19:@44253.4]
  assign regs_180_io_enable = 1'h1; // @[RegFile.scala 74:20:@44247.4]
  assign regs_181_clock = clock; // @[:@44256.4]
  assign regs_181_reset = io_reset; // @[:@44257.4 RegFile.scala 76:16:@44264.4]
  assign regs_181_io_in = 64'h0; // @[RegFile.scala 75:16:@44263.4]
  assign regs_181_io_reset = reset; // @[RegFile.scala 78:19:@44267.4]
  assign regs_181_io_enable = 1'h1; // @[RegFile.scala 74:20:@44261.4]
  assign regs_182_clock = clock; // @[:@44270.4]
  assign regs_182_reset = io_reset; // @[:@44271.4 RegFile.scala 76:16:@44278.4]
  assign regs_182_io_in = 64'h0; // @[RegFile.scala 75:16:@44277.4]
  assign regs_182_io_reset = reset; // @[RegFile.scala 78:19:@44281.4]
  assign regs_182_io_enable = 1'h1; // @[RegFile.scala 74:20:@44275.4]
  assign regs_183_clock = clock; // @[:@44284.4]
  assign regs_183_reset = io_reset; // @[:@44285.4 RegFile.scala 76:16:@44292.4]
  assign regs_183_io_in = 64'h0; // @[RegFile.scala 75:16:@44291.4]
  assign regs_183_io_reset = reset; // @[RegFile.scala 78:19:@44295.4]
  assign regs_183_io_enable = 1'h1; // @[RegFile.scala 74:20:@44289.4]
  assign regs_184_clock = clock; // @[:@44298.4]
  assign regs_184_reset = io_reset; // @[:@44299.4 RegFile.scala 76:16:@44306.4]
  assign regs_184_io_in = 64'h0; // @[RegFile.scala 75:16:@44305.4]
  assign regs_184_io_reset = reset; // @[RegFile.scala 78:19:@44309.4]
  assign regs_184_io_enable = 1'h1; // @[RegFile.scala 74:20:@44303.4]
  assign regs_185_clock = clock; // @[:@44312.4]
  assign regs_185_reset = io_reset; // @[:@44313.4 RegFile.scala 76:16:@44320.4]
  assign regs_185_io_in = 64'h0; // @[RegFile.scala 75:16:@44319.4]
  assign regs_185_io_reset = reset; // @[RegFile.scala 78:19:@44323.4]
  assign regs_185_io_enable = 1'h1; // @[RegFile.scala 74:20:@44317.4]
  assign regs_186_clock = clock; // @[:@44326.4]
  assign regs_186_reset = io_reset; // @[:@44327.4 RegFile.scala 76:16:@44334.4]
  assign regs_186_io_in = 64'h0; // @[RegFile.scala 75:16:@44333.4]
  assign regs_186_io_reset = reset; // @[RegFile.scala 78:19:@44337.4]
  assign regs_186_io_enable = 1'h1; // @[RegFile.scala 74:20:@44331.4]
  assign regs_187_clock = clock; // @[:@44340.4]
  assign regs_187_reset = io_reset; // @[:@44341.4 RegFile.scala 76:16:@44348.4]
  assign regs_187_io_in = 64'h0; // @[RegFile.scala 75:16:@44347.4]
  assign regs_187_io_reset = reset; // @[RegFile.scala 78:19:@44351.4]
  assign regs_187_io_enable = 1'h1; // @[RegFile.scala 74:20:@44345.4]
  assign regs_188_clock = clock; // @[:@44354.4]
  assign regs_188_reset = io_reset; // @[:@44355.4 RegFile.scala 76:16:@44362.4]
  assign regs_188_io_in = 64'h0; // @[RegFile.scala 75:16:@44361.4]
  assign regs_188_io_reset = reset; // @[RegFile.scala 78:19:@44365.4]
  assign regs_188_io_enable = 1'h1; // @[RegFile.scala 74:20:@44359.4]
  assign regs_189_clock = clock; // @[:@44368.4]
  assign regs_189_reset = io_reset; // @[:@44369.4 RegFile.scala 76:16:@44376.4]
  assign regs_189_io_in = 64'h0; // @[RegFile.scala 75:16:@44375.4]
  assign regs_189_io_reset = reset; // @[RegFile.scala 78:19:@44379.4]
  assign regs_189_io_enable = 1'h1; // @[RegFile.scala 74:20:@44373.4]
  assign regs_190_clock = clock; // @[:@44382.4]
  assign regs_190_reset = io_reset; // @[:@44383.4 RegFile.scala 76:16:@44390.4]
  assign regs_190_io_in = 64'h0; // @[RegFile.scala 75:16:@44389.4]
  assign regs_190_io_reset = reset; // @[RegFile.scala 78:19:@44393.4]
  assign regs_190_io_enable = 1'h1; // @[RegFile.scala 74:20:@44387.4]
  assign regs_191_clock = clock; // @[:@44396.4]
  assign regs_191_reset = io_reset; // @[:@44397.4 RegFile.scala 76:16:@44404.4]
  assign regs_191_io_in = 64'h0; // @[RegFile.scala 75:16:@44403.4]
  assign regs_191_io_reset = reset; // @[RegFile.scala 78:19:@44407.4]
  assign regs_191_io_enable = 1'h1; // @[RegFile.scala 74:20:@44401.4]
  assign regs_192_clock = clock; // @[:@44410.4]
  assign regs_192_reset = io_reset; // @[:@44411.4 RegFile.scala 76:16:@44418.4]
  assign regs_192_io_in = 64'h0; // @[RegFile.scala 75:16:@44417.4]
  assign regs_192_io_reset = reset; // @[RegFile.scala 78:19:@44421.4]
  assign regs_192_io_enable = 1'h1; // @[RegFile.scala 74:20:@44415.4]
  assign regs_193_clock = clock; // @[:@44424.4]
  assign regs_193_reset = io_reset; // @[:@44425.4 RegFile.scala 76:16:@44432.4]
  assign regs_193_io_in = 64'h0; // @[RegFile.scala 75:16:@44431.4]
  assign regs_193_io_reset = reset; // @[RegFile.scala 78:19:@44435.4]
  assign regs_193_io_enable = 1'h1; // @[RegFile.scala 74:20:@44429.4]
  assign regs_194_clock = clock; // @[:@44438.4]
  assign regs_194_reset = io_reset; // @[:@44439.4 RegFile.scala 76:16:@44446.4]
  assign regs_194_io_in = 64'h0; // @[RegFile.scala 75:16:@44445.4]
  assign regs_194_io_reset = reset; // @[RegFile.scala 78:19:@44449.4]
  assign regs_194_io_enable = 1'h1; // @[RegFile.scala 74:20:@44443.4]
  assign regs_195_clock = clock; // @[:@44452.4]
  assign regs_195_reset = io_reset; // @[:@44453.4 RegFile.scala 76:16:@44460.4]
  assign regs_195_io_in = 64'h0; // @[RegFile.scala 75:16:@44459.4]
  assign regs_195_io_reset = reset; // @[RegFile.scala 78:19:@44463.4]
  assign regs_195_io_enable = 1'h1; // @[RegFile.scala 74:20:@44457.4]
  assign regs_196_clock = clock; // @[:@44466.4]
  assign regs_196_reset = io_reset; // @[:@44467.4 RegFile.scala 76:16:@44474.4]
  assign regs_196_io_in = 64'h0; // @[RegFile.scala 75:16:@44473.4]
  assign regs_196_io_reset = reset; // @[RegFile.scala 78:19:@44477.4]
  assign regs_196_io_enable = 1'h1; // @[RegFile.scala 74:20:@44471.4]
  assign regs_197_clock = clock; // @[:@44480.4]
  assign regs_197_reset = io_reset; // @[:@44481.4 RegFile.scala 76:16:@44488.4]
  assign regs_197_io_in = 64'h0; // @[RegFile.scala 75:16:@44487.4]
  assign regs_197_io_reset = reset; // @[RegFile.scala 78:19:@44491.4]
  assign regs_197_io_enable = 1'h1; // @[RegFile.scala 74:20:@44485.4]
  assign regs_198_clock = clock; // @[:@44494.4]
  assign regs_198_reset = io_reset; // @[:@44495.4 RegFile.scala 76:16:@44502.4]
  assign regs_198_io_in = 64'h0; // @[RegFile.scala 75:16:@44501.4]
  assign regs_198_io_reset = reset; // @[RegFile.scala 78:19:@44505.4]
  assign regs_198_io_enable = 1'h1; // @[RegFile.scala 74:20:@44499.4]
  assign regs_199_clock = clock; // @[:@44508.4]
  assign regs_199_reset = io_reset; // @[:@44509.4 RegFile.scala 76:16:@44516.4]
  assign regs_199_io_in = 64'h0; // @[RegFile.scala 75:16:@44515.4]
  assign regs_199_io_reset = reset; // @[RegFile.scala 78:19:@44519.4]
  assign regs_199_io_enable = 1'h1; // @[RegFile.scala 74:20:@44513.4]
  assign regs_200_clock = clock; // @[:@44522.4]
  assign regs_200_reset = io_reset; // @[:@44523.4 RegFile.scala 76:16:@44530.4]
  assign regs_200_io_in = 64'h0; // @[RegFile.scala 75:16:@44529.4]
  assign regs_200_io_reset = reset; // @[RegFile.scala 78:19:@44533.4]
  assign regs_200_io_enable = 1'h1; // @[RegFile.scala 74:20:@44527.4]
  assign regs_201_clock = clock; // @[:@44536.4]
  assign regs_201_reset = io_reset; // @[:@44537.4 RegFile.scala 76:16:@44544.4]
  assign regs_201_io_in = 64'h0; // @[RegFile.scala 75:16:@44543.4]
  assign regs_201_io_reset = reset; // @[RegFile.scala 78:19:@44547.4]
  assign regs_201_io_enable = 1'h1; // @[RegFile.scala 74:20:@44541.4]
  assign regs_202_clock = clock; // @[:@44550.4]
  assign regs_202_reset = io_reset; // @[:@44551.4 RegFile.scala 76:16:@44558.4]
  assign regs_202_io_in = 64'h0; // @[RegFile.scala 75:16:@44557.4]
  assign regs_202_io_reset = reset; // @[RegFile.scala 78:19:@44561.4]
  assign regs_202_io_enable = 1'h1; // @[RegFile.scala 74:20:@44555.4]
  assign regs_203_clock = clock; // @[:@44564.4]
  assign regs_203_reset = io_reset; // @[:@44565.4 RegFile.scala 76:16:@44572.4]
  assign regs_203_io_in = 64'h0; // @[RegFile.scala 75:16:@44571.4]
  assign regs_203_io_reset = reset; // @[RegFile.scala 78:19:@44575.4]
  assign regs_203_io_enable = 1'h1; // @[RegFile.scala 74:20:@44569.4]
  assign regs_204_clock = clock; // @[:@44578.4]
  assign regs_204_reset = io_reset; // @[:@44579.4 RegFile.scala 76:16:@44586.4]
  assign regs_204_io_in = 64'h0; // @[RegFile.scala 75:16:@44585.4]
  assign regs_204_io_reset = reset; // @[RegFile.scala 78:19:@44589.4]
  assign regs_204_io_enable = 1'h1; // @[RegFile.scala 74:20:@44583.4]
  assign regs_205_clock = clock; // @[:@44592.4]
  assign regs_205_reset = io_reset; // @[:@44593.4 RegFile.scala 76:16:@44600.4]
  assign regs_205_io_in = 64'h0; // @[RegFile.scala 75:16:@44599.4]
  assign regs_205_io_reset = reset; // @[RegFile.scala 78:19:@44603.4]
  assign regs_205_io_enable = 1'h1; // @[RegFile.scala 74:20:@44597.4]
  assign regs_206_clock = clock; // @[:@44606.4]
  assign regs_206_reset = io_reset; // @[:@44607.4 RegFile.scala 76:16:@44614.4]
  assign regs_206_io_in = 64'h0; // @[RegFile.scala 75:16:@44613.4]
  assign regs_206_io_reset = reset; // @[RegFile.scala 78:19:@44617.4]
  assign regs_206_io_enable = 1'h1; // @[RegFile.scala 74:20:@44611.4]
  assign regs_207_clock = clock; // @[:@44620.4]
  assign regs_207_reset = io_reset; // @[:@44621.4 RegFile.scala 76:16:@44628.4]
  assign regs_207_io_in = 64'h0; // @[RegFile.scala 75:16:@44627.4]
  assign regs_207_io_reset = reset; // @[RegFile.scala 78:19:@44631.4]
  assign regs_207_io_enable = 1'h1; // @[RegFile.scala 74:20:@44625.4]
  assign regs_208_clock = clock; // @[:@44634.4]
  assign regs_208_reset = io_reset; // @[:@44635.4 RegFile.scala 76:16:@44642.4]
  assign regs_208_io_in = 64'h0; // @[RegFile.scala 75:16:@44641.4]
  assign regs_208_io_reset = reset; // @[RegFile.scala 78:19:@44645.4]
  assign regs_208_io_enable = 1'h1; // @[RegFile.scala 74:20:@44639.4]
  assign regs_209_clock = clock; // @[:@44648.4]
  assign regs_209_reset = io_reset; // @[:@44649.4 RegFile.scala 76:16:@44656.4]
  assign regs_209_io_in = 64'h0; // @[RegFile.scala 75:16:@44655.4]
  assign regs_209_io_reset = reset; // @[RegFile.scala 78:19:@44659.4]
  assign regs_209_io_enable = 1'h1; // @[RegFile.scala 74:20:@44653.4]
  assign regs_210_clock = clock; // @[:@44662.4]
  assign regs_210_reset = io_reset; // @[:@44663.4 RegFile.scala 76:16:@44670.4]
  assign regs_210_io_in = 64'h0; // @[RegFile.scala 75:16:@44669.4]
  assign regs_210_io_reset = reset; // @[RegFile.scala 78:19:@44673.4]
  assign regs_210_io_enable = 1'h1; // @[RegFile.scala 74:20:@44667.4]
  assign regs_211_clock = clock; // @[:@44676.4]
  assign regs_211_reset = io_reset; // @[:@44677.4 RegFile.scala 76:16:@44684.4]
  assign regs_211_io_in = 64'h0; // @[RegFile.scala 75:16:@44683.4]
  assign regs_211_io_reset = reset; // @[RegFile.scala 78:19:@44687.4]
  assign regs_211_io_enable = 1'h1; // @[RegFile.scala 74:20:@44681.4]
  assign regs_212_clock = clock; // @[:@44690.4]
  assign regs_212_reset = io_reset; // @[:@44691.4 RegFile.scala 76:16:@44698.4]
  assign regs_212_io_in = 64'h0; // @[RegFile.scala 75:16:@44697.4]
  assign regs_212_io_reset = reset; // @[RegFile.scala 78:19:@44701.4]
  assign regs_212_io_enable = 1'h1; // @[RegFile.scala 74:20:@44695.4]
  assign regs_213_clock = clock; // @[:@44704.4]
  assign regs_213_reset = io_reset; // @[:@44705.4 RegFile.scala 76:16:@44712.4]
  assign regs_213_io_in = 64'h0; // @[RegFile.scala 75:16:@44711.4]
  assign regs_213_io_reset = reset; // @[RegFile.scala 78:19:@44715.4]
  assign regs_213_io_enable = 1'h1; // @[RegFile.scala 74:20:@44709.4]
  assign regs_214_clock = clock; // @[:@44718.4]
  assign regs_214_reset = io_reset; // @[:@44719.4 RegFile.scala 76:16:@44726.4]
  assign regs_214_io_in = 64'h0; // @[RegFile.scala 75:16:@44725.4]
  assign regs_214_io_reset = reset; // @[RegFile.scala 78:19:@44729.4]
  assign regs_214_io_enable = 1'h1; // @[RegFile.scala 74:20:@44723.4]
  assign regs_215_clock = clock; // @[:@44732.4]
  assign regs_215_reset = io_reset; // @[:@44733.4 RegFile.scala 76:16:@44740.4]
  assign regs_215_io_in = 64'h0; // @[RegFile.scala 75:16:@44739.4]
  assign regs_215_io_reset = reset; // @[RegFile.scala 78:19:@44743.4]
  assign regs_215_io_enable = 1'h1; // @[RegFile.scala 74:20:@44737.4]
  assign regs_216_clock = clock; // @[:@44746.4]
  assign regs_216_reset = io_reset; // @[:@44747.4 RegFile.scala 76:16:@44754.4]
  assign regs_216_io_in = 64'h0; // @[RegFile.scala 75:16:@44753.4]
  assign regs_216_io_reset = reset; // @[RegFile.scala 78:19:@44757.4]
  assign regs_216_io_enable = 1'h1; // @[RegFile.scala 74:20:@44751.4]
  assign regs_217_clock = clock; // @[:@44760.4]
  assign regs_217_reset = io_reset; // @[:@44761.4 RegFile.scala 76:16:@44768.4]
  assign regs_217_io_in = 64'h0; // @[RegFile.scala 75:16:@44767.4]
  assign regs_217_io_reset = reset; // @[RegFile.scala 78:19:@44771.4]
  assign regs_217_io_enable = 1'h1; // @[RegFile.scala 74:20:@44765.4]
  assign regs_218_clock = clock; // @[:@44774.4]
  assign regs_218_reset = io_reset; // @[:@44775.4 RegFile.scala 76:16:@44782.4]
  assign regs_218_io_in = 64'h0; // @[RegFile.scala 75:16:@44781.4]
  assign regs_218_io_reset = reset; // @[RegFile.scala 78:19:@44785.4]
  assign regs_218_io_enable = 1'h1; // @[RegFile.scala 74:20:@44779.4]
  assign regs_219_clock = clock; // @[:@44788.4]
  assign regs_219_reset = io_reset; // @[:@44789.4 RegFile.scala 76:16:@44796.4]
  assign regs_219_io_in = 64'h0; // @[RegFile.scala 75:16:@44795.4]
  assign regs_219_io_reset = reset; // @[RegFile.scala 78:19:@44799.4]
  assign regs_219_io_enable = 1'h1; // @[RegFile.scala 74:20:@44793.4]
  assign regs_220_clock = clock; // @[:@44802.4]
  assign regs_220_reset = io_reset; // @[:@44803.4 RegFile.scala 76:16:@44810.4]
  assign regs_220_io_in = 64'h0; // @[RegFile.scala 75:16:@44809.4]
  assign regs_220_io_reset = reset; // @[RegFile.scala 78:19:@44813.4]
  assign regs_220_io_enable = 1'h1; // @[RegFile.scala 74:20:@44807.4]
  assign regs_221_clock = clock; // @[:@44816.4]
  assign regs_221_reset = io_reset; // @[:@44817.4 RegFile.scala 76:16:@44824.4]
  assign regs_221_io_in = 64'h0; // @[RegFile.scala 75:16:@44823.4]
  assign regs_221_io_reset = reset; // @[RegFile.scala 78:19:@44827.4]
  assign regs_221_io_enable = 1'h1; // @[RegFile.scala 74:20:@44821.4]
  assign regs_222_clock = clock; // @[:@44830.4]
  assign regs_222_reset = io_reset; // @[:@44831.4 RegFile.scala 76:16:@44838.4]
  assign regs_222_io_in = 64'h0; // @[RegFile.scala 75:16:@44837.4]
  assign regs_222_io_reset = reset; // @[RegFile.scala 78:19:@44841.4]
  assign regs_222_io_enable = 1'h1; // @[RegFile.scala 74:20:@44835.4]
  assign regs_223_clock = clock; // @[:@44844.4]
  assign regs_223_reset = io_reset; // @[:@44845.4 RegFile.scala 76:16:@44852.4]
  assign regs_223_io_in = 64'h0; // @[RegFile.scala 75:16:@44851.4]
  assign regs_223_io_reset = reset; // @[RegFile.scala 78:19:@44855.4]
  assign regs_223_io_enable = 1'h1; // @[RegFile.scala 74:20:@44849.4]
  assign regs_224_clock = clock; // @[:@44858.4]
  assign regs_224_reset = io_reset; // @[:@44859.4 RegFile.scala 76:16:@44866.4]
  assign regs_224_io_in = 64'h0; // @[RegFile.scala 75:16:@44865.4]
  assign regs_224_io_reset = reset; // @[RegFile.scala 78:19:@44869.4]
  assign regs_224_io_enable = 1'h1; // @[RegFile.scala 74:20:@44863.4]
  assign regs_225_clock = clock; // @[:@44872.4]
  assign regs_225_reset = io_reset; // @[:@44873.4 RegFile.scala 76:16:@44880.4]
  assign regs_225_io_in = 64'h0; // @[RegFile.scala 75:16:@44879.4]
  assign regs_225_io_reset = reset; // @[RegFile.scala 78:19:@44883.4]
  assign regs_225_io_enable = 1'h1; // @[RegFile.scala 74:20:@44877.4]
  assign regs_226_clock = clock; // @[:@44886.4]
  assign regs_226_reset = io_reset; // @[:@44887.4 RegFile.scala 76:16:@44894.4]
  assign regs_226_io_in = 64'h0; // @[RegFile.scala 75:16:@44893.4]
  assign regs_226_io_reset = reset; // @[RegFile.scala 78:19:@44897.4]
  assign regs_226_io_enable = 1'h1; // @[RegFile.scala 74:20:@44891.4]
  assign regs_227_clock = clock; // @[:@44900.4]
  assign regs_227_reset = io_reset; // @[:@44901.4 RegFile.scala 76:16:@44908.4]
  assign regs_227_io_in = 64'h0; // @[RegFile.scala 75:16:@44907.4]
  assign regs_227_io_reset = reset; // @[RegFile.scala 78:19:@44911.4]
  assign regs_227_io_enable = 1'h1; // @[RegFile.scala 74:20:@44905.4]
  assign regs_228_clock = clock; // @[:@44914.4]
  assign regs_228_reset = io_reset; // @[:@44915.4 RegFile.scala 76:16:@44922.4]
  assign regs_228_io_in = 64'h0; // @[RegFile.scala 75:16:@44921.4]
  assign regs_228_io_reset = reset; // @[RegFile.scala 78:19:@44925.4]
  assign regs_228_io_enable = 1'h1; // @[RegFile.scala 74:20:@44919.4]
  assign regs_229_clock = clock; // @[:@44928.4]
  assign regs_229_reset = io_reset; // @[:@44929.4 RegFile.scala 76:16:@44936.4]
  assign regs_229_io_in = 64'h0; // @[RegFile.scala 75:16:@44935.4]
  assign regs_229_io_reset = reset; // @[RegFile.scala 78:19:@44939.4]
  assign regs_229_io_enable = 1'h1; // @[RegFile.scala 74:20:@44933.4]
  assign regs_230_clock = clock; // @[:@44942.4]
  assign regs_230_reset = io_reset; // @[:@44943.4 RegFile.scala 76:16:@44950.4]
  assign regs_230_io_in = 64'h0; // @[RegFile.scala 75:16:@44949.4]
  assign regs_230_io_reset = reset; // @[RegFile.scala 78:19:@44953.4]
  assign regs_230_io_enable = 1'h1; // @[RegFile.scala 74:20:@44947.4]
  assign regs_231_clock = clock; // @[:@44956.4]
  assign regs_231_reset = io_reset; // @[:@44957.4 RegFile.scala 76:16:@44964.4]
  assign regs_231_io_in = 64'h0; // @[RegFile.scala 75:16:@44963.4]
  assign regs_231_io_reset = reset; // @[RegFile.scala 78:19:@44967.4]
  assign regs_231_io_enable = 1'h1; // @[RegFile.scala 74:20:@44961.4]
  assign regs_232_clock = clock; // @[:@44970.4]
  assign regs_232_reset = io_reset; // @[:@44971.4 RegFile.scala 76:16:@44978.4]
  assign regs_232_io_in = 64'h0; // @[RegFile.scala 75:16:@44977.4]
  assign regs_232_io_reset = reset; // @[RegFile.scala 78:19:@44981.4]
  assign regs_232_io_enable = 1'h1; // @[RegFile.scala 74:20:@44975.4]
  assign regs_233_clock = clock; // @[:@44984.4]
  assign regs_233_reset = io_reset; // @[:@44985.4 RegFile.scala 76:16:@44992.4]
  assign regs_233_io_in = 64'h0; // @[RegFile.scala 75:16:@44991.4]
  assign regs_233_io_reset = reset; // @[RegFile.scala 78:19:@44995.4]
  assign regs_233_io_enable = 1'h1; // @[RegFile.scala 74:20:@44989.4]
  assign regs_234_clock = clock; // @[:@44998.4]
  assign regs_234_reset = io_reset; // @[:@44999.4 RegFile.scala 76:16:@45006.4]
  assign regs_234_io_in = 64'h0; // @[RegFile.scala 75:16:@45005.4]
  assign regs_234_io_reset = reset; // @[RegFile.scala 78:19:@45009.4]
  assign regs_234_io_enable = 1'h1; // @[RegFile.scala 74:20:@45003.4]
  assign regs_235_clock = clock; // @[:@45012.4]
  assign regs_235_reset = io_reset; // @[:@45013.4 RegFile.scala 76:16:@45020.4]
  assign regs_235_io_in = 64'h0; // @[RegFile.scala 75:16:@45019.4]
  assign regs_235_io_reset = reset; // @[RegFile.scala 78:19:@45023.4]
  assign regs_235_io_enable = 1'h1; // @[RegFile.scala 74:20:@45017.4]
  assign regs_236_clock = clock; // @[:@45026.4]
  assign regs_236_reset = io_reset; // @[:@45027.4 RegFile.scala 76:16:@45034.4]
  assign regs_236_io_in = 64'h0; // @[RegFile.scala 75:16:@45033.4]
  assign regs_236_io_reset = reset; // @[RegFile.scala 78:19:@45037.4]
  assign regs_236_io_enable = 1'h1; // @[RegFile.scala 74:20:@45031.4]
  assign regs_237_clock = clock; // @[:@45040.4]
  assign regs_237_reset = io_reset; // @[:@45041.4 RegFile.scala 76:16:@45048.4]
  assign regs_237_io_in = 64'h0; // @[RegFile.scala 75:16:@45047.4]
  assign regs_237_io_reset = reset; // @[RegFile.scala 78:19:@45051.4]
  assign regs_237_io_enable = 1'h1; // @[RegFile.scala 74:20:@45045.4]
  assign regs_238_clock = clock; // @[:@45054.4]
  assign regs_238_reset = io_reset; // @[:@45055.4 RegFile.scala 76:16:@45062.4]
  assign regs_238_io_in = 64'h0; // @[RegFile.scala 75:16:@45061.4]
  assign regs_238_io_reset = reset; // @[RegFile.scala 78:19:@45065.4]
  assign regs_238_io_enable = 1'h1; // @[RegFile.scala 74:20:@45059.4]
  assign regs_239_clock = clock; // @[:@45068.4]
  assign regs_239_reset = io_reset; // @[:@45069.4 RegFile.scala 76:16:@45076.4]
  assign regs_239_io_in = 64'h0; // @[RegFile.scala 75:16:@45075.4]
  assign regs_239_io_reset = reset; // @[RegFile.scala 78:19:@45079.4]
  assign regs_239_io_enable = 1'h1; // @[RegFile.scala 74:20:@45073.4]
  assign regs_240_clock = clock; // @[:@45082.4]
  assign regs_240_reset = io_reset; // @[:@45083.4 RegFile.scala 76:16:@45090.4]
  assign regs_240_io_in = 64'h0; // @[RegFile.scala 75:16:@45089.4]
  assign regs_240_io_reset = reset; // @[RegFile.scala 78:19:@45093.4]
  assign regs_240_io_enable = 1'h1; // @[RegFile.scala 74:20:@45087.4]
  assign regs_241_clock = clock; // @[:@45096.4]
  assign regs_241_reset = io_reset; // @[:@45097.4 RegFile.scala 76:16:@45104.4]
  assign regs_241_io_in = 64'h0; // @[RegFile.scala 75:16:@45103.4]
  assign regs_241_io_reset = reset; // @[RegFile.scala 78:19:@45107.4]
  assign regs_241_io_enable = 1'h1; // @[RegFile.scala 74:20:@45101.4]
  assign regs_242_clock = clock; // @[:@45110.4]
  assign regs_242_reset = io_reset; // @[:@45111.4 RegFile.scala 76:16:@45118.4]
  assign regs_242_io_in = 64'h0; // @[RegFile.scala 75:16:@45117.4]
  assign regs_242_io_reset = reset; // @[RegFile.scala 78:19:@45121.4]
  assign regs_242_io_enable = 1'h1; // @[RegFile.scala 74:20:@45115.4]
  assign regs_243_clock = clock; // @[:@45124.4]
  assign regs_243_reset = io_reset; // @[:@45125.4 RegFile.scala 76:16:@45132.4]
  assign regs_243_io_in = 64'h0; // @[RegFile.scala 75:16:@45131.4]
  assign regs_243_io_reset = reset; // @[RegFile.scala 78:19:@45135.4]
  assign regs_243_io_enable = 1'h1; // @[RegFile.scala 74:20:@45129.4]
  assign regs_244_clock = clock; // @[:@45138.4]
  assign regs_244_reset = io_reset; // @[:@45139.4 RegFile.scala 76:16:@45146.4]
  assign regs_244_io_in = 64'h0; // @[RegFile.scala 75:16:@45145.4]
  assign regs_244_io_reset = reset; // @[RegFile.scala 78:19:@45149.4]
  assign regs_244_io_enable = 1'h1; // @[RegFile.scala 74:20:@45143.4]
  assign regs_245_clock = clock; // @[:@45152.4]
  assign regs_245_reset = io_reset; // @[:@45153.4 RegFile.scala 76:16:@45160.4]
  assign regs_245_io_in = 64'h0; // @[RegFile.scala 75:16:@45159.4]
  assign regs_245_io_reset = reset; // @[RegFile.scala 78:19:@45163.4]
  assign regs_245_io_enable = 1'h1; // @[RegFile.scala 74:20:@45157.4]
  assign regs_246_clock = clock; // @[:@45166.4]
  assign regs_246_reset = io_reset; // @[:@45167.4 RegFile.scala 76:16:@45174.4]
  assign regs_246_io_in = 64'h0; // @[RegFile.scala 75:16:@45173.4]
  assign regs_246_io_reset = reset; // @[RegFile.scala 78:19:@45177.4]
  assign regs_246_io_enable = 1'h1; // @[RegFile.scala 74:20:@45171.4]
  assign regs_247_clock = clock; // @[:@45180.4]
  assign regs_247_reset = io_reset; // @[:@45181.4 RegFile.scala 76:16:@45188.4]
  assign regs_247_io_in = 64'h0; // @[RegFile.scala 75:16:@45187.4]
  assign regs_247_io_reset = reset; // @[RegFile.scala 78:19:@45191.4]
  assign regs_247_io_enable = 1'h1; // @[RegFile.scala 74:20:@45185.4]
  assign regs_248_clock = clock; // @[:@45194.4]
  assign regs_248_reset = io_reset; // @[:@45195.4 RegFile.scala 76:16:@45202.4]
  assign regs_248_io_in = 64'h0; // @[RegFile.scala 75:16:@45201.4]
  assign regs_248_io_reset = reset; // @[RegFile.scala 78:19:@45205.4]
  assign regs_248_io_enable = 1'h1; // @[RegFile.scala 74:20:@45199.4]
  assign regs_249_clock = clock; // @[:@45208.4]
  assign regs_249_reset = io_reset; // @[:@45209.4 RegFile.scala 76:16:@45216.4]
  assign regs_249_io_in = 64'h0; // @[RegFile.scala 75:16:@45215.4]
  assign regs_249_io_reset = reset; // @[RegFile.scala 78:19:@45219.4]
  assign regs_249_io_enable = 1'h1; // @[RegFile.scala 74:20:@45213.4]
  assign regs_250_clock = clock; // @[:@45222.4]
  assign regs_250_reset = io_reset; // @[:@45223.4 RegFile.scala 76:16:@45230.4]
  assign regs_250_io_in = 64'h0; // @[RegFile.scala 75:16:@45229.4]
  assign regs_250_io_reset = reset; // @[RegFile.scala 78:19:@45233.4]
  assign regs_250_io_enable = 1'h1; // @[RegFile.scala 74:20:@45227.4]
  assign regs_251_clock = clock; // @[:@45236.4]
  assign regs_251_reset = io_reset; // @[:@45237.4 RegFile.scala 76:16:@45244.4]
  assign regs_251_io_in = 64'h0; // @[RegFile.scala 75:16:@45243.4]
  assign regs_251_io_reset = reset; // @[RegFile.scala 78:19:@45247.4]
  assign regs_251_io_enable = 1'h1; // @[RegFile.scala 74:20:@45241.4]
  assign regs_252_clock = clock; // @[:@45250.4]
  assign regs_252_reset = io_reset; // @[:@45251.4 RegFile.scala 76:16:@45258.4]
  assign regs_252_io_in = 64'h0; // @[RegFile.scala 75:16:@45257.4]
  assign regs_252_io_reset = reset; // @[RegFile.scala 78:19:@45261.4]
  assign regs_252_io_enable = 1'h1; // @[RegFile.scala 74:20:@45255.4]
  assign regs_253_clock = clock; // @[:@45264.4]
  assign regs_253_reset = io_reset; // @[:@45265.4 RegFile.scala 76:16:@45272.4]
  assign regs_253_io_in = 64'h0; // @[RegFile.scala 75:16:@45271.4]
  assign regs_253_io_reset = reset; // @[RegFile.scala 78:19:@45275.4]
  assign regs_253_io_enable = 1'h1; // @[RegFile.scala 74:20:@45269.4]
  assign regs_254_clock = clock; // @[:@45278.4]
  assign regs_254_reset = io_reset; // @[:@45279.4 RegFile.scala 76:16:@45286.4]
  assign regs_254_io_in = 64'h0; // @[RegFile.scala 75:16:@45285.4]
  assign regs_254_io_reset = reset; // @[RegFile.scala 78:19:@45289.4]
  assign regs_254_io_enable = 1'h1; // @[RegFile.scala 74:20:@45283.4]
  assign regs_255_clock = clock; // @[:@45292.4]
  assign regs_255_reset = io_reset; // @[:@45293.4 RegFile.scala 76:16:@45300.4]
  assign regs_255_io_in = 64'h0; // @[RegFile.scala 75:16:@45299.4]
  assign regs_255_io_reset = reset; // @[RegFile.scala 78:19:@45303.4]
  assign regs_255_io_enable = 1'h1; // @[RegFile.scala 74:20:@45297.4]
  assign regs_256_clock = clock; // @[:@45306.4]
  assign regs_256_reset = io_reset; // @[:@45307.4 RegFile.scala 76:16:@45314.4]
  assign regs_256_io_in = 64'h0; // @[RegFile.scala 75:16:@45313.4]
  assign regs_256_io_reset = reset; // @[RegFile.scala 78:19:@45317.4]
  assign regs_256_io_enable = 1'h1; // @[RegFile.scala 74:20:@45311.4]
  assign regs_257_clock = clock; // @[:@45320.4]
  assign regs_257_reset = io_reset; // @[:@45321.4 RegFile.scala 76:16:@45328.4]
  assign regs_257_io_in = 64'h0; // @[RegFile.scala 75:16:@45327.4]
  assign regs_257_io_reset = reset; // @[RegFile.scala 78:19:@45331.4]
  assign regs_257_io_enable = 1'h1; // @[RegFile.scala 74:20:@45325.4]
  assign regs_258_clock = clock; // @[:@45334.4]
  assign regs_258_reset = io_reset; // @[:@45335.4 RegFile.scala 76:16:@45342.4]
  assign regs_258_io_in = 64'h0; // @[RegFile.scala 75:16:@45341.4]
  assign regs_258_io_reset = reset; // @[RegFile.scala 78:19:@45345.4]
  assign regs_258_io_enable = 1'h1; // @[RegFile.scala 74:20:@45339.4]
  assign regs_259_clock = clock; // @[:@45348.4]
  assign regs_259_reset = io_reset; // @[:@45349.4 RegFile.scala 76:16:@45356.4]
  assign regs_259_io_in = 64'h0; // @[RegFile.scala 75:16:@45355.4]
  assign regs_259_io_reset = reset; // @[RegFile.scala 78:19:@45359.4]
  assign regs_259_io_enable = 1'h1; // @[RegFile.scala 74:20:@45353.4]
  assign regs_260_clock = clock; // @[:@45362.4]
  assign regs_260_reset = io_reset; // @[:@45363.4 RegFile.scala 76:16:@45370.4]
  assign regs_260_io_in = 64'h0; // @[RegFile.scala 75:16:@45369.4]
  assign regs_260_io_reset = reset; // @[RegFile.scala 78:19:@45373.4]
  assign regs_260_io_enable = 1'h1; // @[RegFile.scala 74:20:@45367.4]
  assign regs_261_clock = clock; // @[:@45376.4]
  assign regs_261_reset = io_reset; // @[:@45377.4 RegFile.scala 76:16:@45384.4]
  assign regs_261_io_in = 64'h0; // @[RegFile.scala 75:16:@45383.4]
  assign regs_261_io_reset = reset; // @[RegFile.scala 78:19:@45387.4]
  assign regs_261_io_enable = 1'h1; // @[RegFile.scala 74:20:@45381.4]
  assign regs_262_clock = clock; // @[:@45390.4]
  assign regs_262_reset = io_reset; // @[:@45391.4 RegFile.scala 76:16:@45398.4]
  assign regs_262_io_in = 64'h0; // @[RegFile.scala 75:16:@45397.4]
  assign regs_262_io_reset = reset; // @[RegFile.scala 78:19:@45401.4]
  assign regs_262_io_enable = 1'h1; // @[RegFile.scala 74:20:@45395.4]
  assign regs_263_clock = clock; // @[:@45404.4]
  assign regs_263_reset = io_reset; // @[:@45405.4 RegFile.scala 76:16:@45412.4]
  assign regs_263_io_in = 64'h0; // @[RegFile.scala 75:16:@45411.4]
  assign regs_263_io_reset = reset; // @[RegFile.scala 78:19:@45415.4]
  assign regs_263_io_enable = 1'h1; // @[RegFile.scala 74:20:@45409.4]
  assign regs_264_clock = clock; // @[:@45418.4]
  assign regs_264_reset = io_reset; // @[:@45419.4 RegFile.scala 76:16:@45426.4]
  assign regs_264_io_in = 64'h0; // @[RegFile.scala 75:16:@45425.4]
  assign regs_264_io_reset = reset; // @[RegFile.scala 78:19:@45429.4]
  assign regs_264_io_enable = 1'h1; // @[RegFile.scala 74:20:@45423.4]
  assign regs_265_clock = clock; // @[:@45432.4]
  assign regs_265_reset = io_reset; // @[:@45433.4 RegFile.scala 76:16:@45440.4]
  assign regs_265_io_in = 64'h0; // @[RegFile.scala 75:16:@45439.4]
  assign regs_265_io_reset = reset; // @[RegFile.scala 78:19:@45443.4]
  assign regs_265_io_enable = 1'h1; // @[RegFile.scala 74:20:@45437.4]
  assign regs_266_clock = clock; // @[:@45446.4]
  assign regs_266_reset = io_reset; // @[:@45447.4 RegFile.scala 76:16:@45454.4]
  assign regs_266_io_in = 64'h0; // @[RegFile.scala 75:16:@45453.4]
  assign regs_266_io_reset = reset; // @[RegFile.scala 78:19:@45457.4]
  assign regs_266_io_enable = 1'h1; // @[RegFile.scala 74:20:@45451.4]
  assign regs_267_clock = clock; // @[:@45460.4]
  assign regs_267_reset = io_reset; // @[:@45461.4 RegFile.scala 76:16:@45468.4]
  assign regs_267_io_in = 64'h0; // @[RegFile.scala 75:16:@45467.4]
  assign regs_267_io_reset = reset; // @[RegFile.scala 78:19:@45471.4]
  assign regs_267_io_enable = 1'h1; // @[RegFile.scala 74:20:@45465.4]
  assign regs_268_clock = clock; // @[:@45474.4]
  assign regs_268_reset = io_reset; // @[:@45475.4 RegFile.scala 76:16:@45482.4]
  assign regs_268_io_in = 64'h0; // @[RegFile.scala 75:16:@45481.4]
  assign regs_268_io_reset = reset; // @[RegFile.scala 78:19:@45485.4]
  assign regs_268_io_enable = 1'h1; // @[RegFile.scala 74:20:@45479.4]
  assign regs_269_clock = clock; // @[:@45488.4]
  assign regs_269_reset = io_reset; // @[:@45489.4 RegFile.scala 76:16:@45496.4]
  assign regs_269_io_in = 64'h0; // @[RegFile.scala 75:16:@45495.4]
  assign regs_269_io_reset = reset; // @[RegFile.scala 78:19:@45499.4]
  assign regs_269_io_enable = 1'h1; // @[RegFile.scala 74:20:@45493.4]
  assign regs_270_clock = clock; // @[:@45502.4]
  assign regs_270_reset = io_reset; // @[:@45503.4 RegFile.scala 76:16:@45510.4]
  assign regs_270_io_in = 64'h0; // @[RegFile.scala 75:16:@45509.4]
  assign regs_270_io_reset = reset; // @[RegFile.scala 78:19:@45513.4]
  assign regs_270_io_enable = 1'h1; // @[RegFile.scala 74:20:@45507.4]
  assign regs_271_clock = clock; // @[:@45516.4]
  assign regs_271_reset = io_reset; // @[:@45517.4 RegFile.scala 76:16:@45524.4]
  assign regs_271_io_in = 64'h0; // @[RegFile.scala 75:16:@45523.4]
  assign regs_271_io_reset = reset; // @[RegFile.scala 78:19:@45527.4]
  assign regs_271_io_enable = 1'h1; // @[RegFile.scala 74:20:@45521.4]
  assign regs_272_clock = clock; // @[:@45530.4]
  assign regs_272_reset = io_reset; // @[:@45531.4 RegFile.scala 76:16:@45538.4]
  assign regs_272_io_in = 64'h0; // @[RegFile.scala 75:16:@45537.4]
  assign regs_272_io_reset = reset; // @[RegFile.scala 78:19:@45541.4]
  assign regs_272_io_enable = 1'h1; // @[RegFile.scala 74:20:@45535.4]
  assign regs_273_clock = clock; // @[:@45544.4]
  assign regs_273_reset = io_reset; // @[:@45545.4 RegFile.scala 76:16:@45552.4]
  assign regs_273_io_in = 64'h0; // @[RegFile.scala 75:16:@45551.4]
  assign regs_273_io_reset = reset; // @[RegFile.scala 78:19:@45555.4]
  assign regs_273_io_enable = 1'h1; // @[RegFile.scala 74:20:@45549.4]
  assign regs_274_clock = clock; // @[:@45558.4]
  assign regs_274_reset = io_reset; // @[:@45559.4 RegFile.scala 76:16:@45566.4]
  assign regs_274_io_in = 64'h0; // @[RegFile.scala 75:16:@45565.4]
  assign regs_274_io_reset = reset; // @[RegFile.scala 78:19:@45569.4]
  assign regs_274_io_enable = 1'h1; // @[RegFile.scala 74:20:@45563.4]
  assign regs_275_clock = clock; // @[:@45572.4]
  assign regs_275_reset = io_reset; // @[:@45573.4 RegFile.scala 76:16:@45580.4]
  assign regs_275_io_in = 64'h0; // @[RegFile.scala 75:16:@45579.4]
  assign regs_275_io_reset = reset; // @[RegFile.scala 78:19:@45583.4]
  assign regs_275_io_enable = 1'h1; // @[RegFile.scala 74:20:@45577.4]
  assign regs_276_clock = clock; // @[:@45586.4]
  assign regs_276_reset = io_reset; // @[:@45587.4 RegFile.scala 76:16:@45594.4]
  assign regs_276_io_in = 64'h0; // @[RegFile.scala 75:16:@45593.4]
  assign regs_276_io_reset = reset; // @[RegFile.scala 78:19:@45597.4]
  assign regs_276_io_enable = 1'h1; // @[RegFile.scala 74:20:@45591.4]
  assign regs_277_clock = clock; // @[:@45600.4]
  assign regs_277_reset = io_reset; // @[:@45601.4 RegFile.scala 76:16:@45608.4]
  assign regs_277_io_in = 64'h0; // @[RegFile.scala 75:16:@45607.4]
  assign regs_277_io_reset = reset; // @[RegFile.scala 78:19:@45611.4]
  assign regs_277_io_enable = 1'h1; // @[RegFile.scala 74:20:@45605.4]
  assign regs_278_clock = clock; // @[:@45614.4]
  assign regs_278_reset = io_reset; // @[:@45615.4 RegFile.scala 76:16:@45622.4]
  assign regs_278_io_in = 64'h0; // @[RegFile.scala 75:16:@45621.4]
  assign regs_278_io_reset = reset; // @[RegFile.scala 78:19:@45625.4]
  assign regs_278_io_enable = 1'h1; // @[RegFile.scala 74:20:@45619.4]
  assign regs_279_clock = clock; // @[:@45628.4]
  assign regs_279_reset = io_reset; // @[:@45629.4 RegFile.scala 76:16:@45636.4]
  assign regs_279_io_in = 64'h0; // @[RegFile.scala 75:16:@45635.4]
  assign regs_279_io_reset = reset; // @[RegFile.scala 78:19:@45639.4]
  assign regs_279_io_enable = 1'h1; // @[RegFile.scala 74:20:@45633.4]
  assign regs_280_clock = clock; // @[:@45642.4]
  assign regs_280_reset = io_reset; // @[:@45643.4 RegFile.scala 76:16:@45650.4]
  assign regs_280_io_in = 64'h0; // @[RegFile.scala 75:16:@45649.4]
  assign regs_280_io_reset = reset; // @[RegFile.scala 78:19:@45653.4]
  assign regs_280_io_enable = 1'h1; // @[RegFile.scala 74:20:@45647.4]
  assign regs_281_clock = clock; // @[:@45656.4]
  assign regs_281_reset = io_reset; // @[:@45657.4 RegFile.scala 76:16:@45664.4]
  assign regs_281_io_in = 64'h0; // @[RegFile.scala 75:16:@45663.4]
  assign regs_281_io_reset = reset; // @[RegFile.scala 78:19:@45667.4]
  assign regs_281_io_enable = 1'h1; // @[RegFile.scala 74:20:@45661.4]
  assign regs_282_clock = clock; // @[:@45670.4]
  assign regs_282_reset = io_reset; // @[:@45671.4 RegFile.scala 76:16:@45678.4]
  assign regs_282_io_in = 64'h0; // @[RegFile.scala 75:16:@45677.4]
  assign regs_282_io_reset = reset; // @[RegFile.scala 78:19:@45681.4]
  assign regs_282_io_enable = 1'h1; // @[RegFile.scala 74:20:@45675.4]
  assign regs_283_clock = clock; // @[:@45684.4]
  assign regs_283_reset = io_reset; // @[:@45685.4 RegFile.scala 76:16:@45692.4]
  assign regs_283_io_in = 64'h0; // @[RegFile.scala 75:16:@45691.4]
  assign regs_283_io_reset = reset; // @[RegFile.scala 78:19:@45695.4]
  assign regs_283_io_enable = 1'h1; // @[RegFile.scala 74:20:@45689.4]
  assign regs_284_clock = clock; // @[:@45698.4]
  assign regs_284_reset = io_reset; // @[:@45699.4 RegFile.scala 76:16:@45706.4]
  assign regs_284_io_in = 64'h0; // @[RegFile.scala 75:16:@45705.4]
  assign regs_284_io_reset = reset; // @[RegFile.scala 78:19:@45709.4]
  assign regs_284_io_enable = 1'h1; // @[RegFile.scala 74:20:@45703.4]
  assign regs_285_clock = clock; // @[:@45712.4]
  assign regs_285_reset = io_reset; // @[:@45713.4 RegFile.scala 76:16:@45720.4]
  assign regs_285_io_in = 64'h0; // @[RegFile.scala 75:16:@45719.4]
  assign regs_285_io_reset = reset; // @[RegFile.scala 78:19:@45723.4]
  assign regs_285_io_enable = 1'h1; // @[RegFile.scala 74:20:@45717.4]
  assign regs_286_clock = clock; // @[:@45726.4]
  assign regs_286_reset = io_reset; // @[:@45727.4 RegFile.scala 76:16:@45734.4]
  assign regs_286_io_in = 64'h0; // @[RegFile.scala 75:16:@45733.4]
  assign regs_286_io_reset = reset; // @[RegFile.scala 78:19:@45737.4]
  assign regs_286_io_enable = 1'h1; // @[RegFile.scala 74:20:@45731.4]
  assign regs_287_clock = clock; // @[:@45740.4]
  assign regs_287_reset = io_reset; // @[:@45741.4 RegFile.scala 76:16:@45748.4]
  assign regs_287_io_in = 64'h0; // @[RegFile.scala 75:16:@45747.4]
  assign regs_287_io_reset = reset; // @[RegFile.scala 78:19:@45751.4]
  assign regs_287_io_enable = 1'h1; // @[RegFile.scala 74:20:@45745.4]
  assign regs_288_clock = clock; // @[:@45754.4]
  assign regs_288_reset = io_reset; // @[:@45755.4 RegFile.scala 76:16:@45762.4]
  assign regs_288_io_in = 64'h0; // @[RegFile.scala 75:16:@45761.4]
  assign regs_288_io_reset = reset; // @[RegFile.scala 78:19:@45765.4]
  assign regs_288_io_enable = 1'h1; // @[RegFile.scala 74:20:@45759.4]
  assign regs_289_clock = clock; // @[:@45768.4]
  assign regs_289_reset = io_reset; // @[:@45769.4 RegFile.scala 76:16:@45776.4]
  assign regs_289_io_in = 64'h0; // @[RegFile.scala 75:16:@45775.4]
  assign regs_289_io_reset = reset; // @[RegFile.scala 78:19:@45779.4]
  assign regs_289_io_enable = 1'h1; // @[RegFile.scala 74:20:@45773.4]
  assign regs_290_clock = clock; // @[:@45782.4]
  assign regs_290_reset = io_reset; // @[:@45783.4 RegFile.scala 76:16:@45790.4]
  assign regs_290_io_in = 64'h0; // @[RegFile.scala 75:16:@45789.4]
  assign regs_290_io_reset = reset; // @[RegFile.scala 78:19:@45793.4]
  assign regs_290_io_enable = 1'h1; // @[RegFile.scala 74:20:@45787.4]
  assign regs_291_clock = clock; // @[:@45796.4]
  assign regs_291_reset = io_reset; // @[:@45797.4 RegFile.scala 76:16:@45804.4]
  assign regs_291_io_in = 64'h0; // @[RegFile.scala 75:16:@45803.4]
  assign regs_291_io_reset = reset; // @[RegFile.scala 78:19:@45807.4]
  assign regs_291_io_enable = 1'h1; // @[RegFile.scala 74:20:@45801.4]
  assign regs_292_clock = clock; // @[:@45810.4]
  assign regs_292_reset = io_reset; // @[:@45811.4 RegFile.scala 76:16:@45818.4]
  assign regs_292_io_in = 64'h0; // @[RegFile.scala 75:16:@45817.4]
  assign regs_292_io_reset = reset; // @[RegFile.scala 78:19:@45821.4]
  assign regs_292_io_enable = 1'h1; // @[RegFile.scala 74:20:@45815.4]
  assign regs_293_clock = clock; // @[:@45824.4]
  assign regs_293_reset = io_reset; // @[:@45825.4 RegFile.scala 76:16:@45832.4]
  assign regs_293_io_in = 64'h0; // @[RegFile.scala 75:16:@45831.4]
  assign regs_293_io_reset = reset; // @[RegFile.scala 78:19:@45835.4]
  assign regs_293_io_enable = 1'h1; // @[RegFile.scala 74:20:@45829.4]
  assign regs_294_clock = clock; // @[:@45838.4]
  assign regs_294_reset = io_reset; // @[:@45839.4 RegFile.scala 76:16:@45846.4]
  assign regs_294_io_in = 64'h0; // @[RegFile.scala 75:16:@45845.4]
  assign regs_294_io_reset = reset; // @[RegFile.scala 78:19:@45849.4]
  assign regs_294_io_enable = 1'h1; // @[RegFile.scala 74:20:@45843.4]
  assign regs_295_clock = clock; // @[:@45852.4]
  assign regs_295_reset = io_reset; // @[:@45853.4 RegFile.scala 76:16:@45860.4]
  assign regs_295_io_in = 64'h0; // @[RegFile.scala 75:16:@45859.4]
  assign regs_295_io_reset = reset; // @[RegFile.scala 78:19:@45863.4]
  assign regs_295_io_enable = 1'h1; // @[RegFile.scala 74:20:@45857.4]
  assign regs_296_clock = clock; // @[:@45866.4]
  assign regs_296_reset = io_reset; // @[:@45867.4 RegFile.scala 76:16:@45874.4]
  assign regs_296_io_in = 64'h0; // @[RegFile.scala 75:16:@45873.4]
  assign regs_296_io_reset = reset; // @[RegFile.scala 78:19:@45877.4]
  assign regs_296_io_enable = 1'h1; // @[RegFile.scala 74:20:@45871.4]
  assign regs_297_clock = clock; // @[:@45880.4]
  assign regs_297_reset = io_reset; // @[:@45881.4 RegFile.scala 76:16:@45888.4]
  assign regs_297_io_in = 64'h0; // @[RegFile.scala 75:16:@45887.4]
  assign regs_297_io_reset = reset; // @[RegFile.scala 78:19:@45891.4]
  assign regs_297_io_enable = 1'h1; // @[RegFile.scala 74:20:@45885.4]
  assign regs_298_clock = clock; // @[:@45894.4]
  assign regs_298_reset = io_reset; // @[:@45895.4 RegFile.scala 76:16:@45902.4]
  assign regs_298_io_in = 64'h0; // @[RegFile.scala 75:16:@45901.4]
  assign regs_298_io_reset = reset; // @[RegFile.scala 78:19:@45905.4]
  assign regs_298_io_enable = 1'h1; // @[RegFile.scala 74:20:@45899.4]
  assign regs_299_clock = clock; // @[:@45908.4]
  assign regs_299_reset = io_reset; // @[:@45909.4 RegFile.scala 76:16:@45916.4]
  assign regs_299_io_in = 64'h0; // @[RegFile.scala 75:16:@45915.4]
  assign regs_299_io_reset = reset; // @[RegFile.scala 78:19:@45919.4]
  assign regs_299_io_enable = 1'h1; // @[RegFile.scala 74:20:@45913.4]
  assign regs_300_clock = clock; // @[:@45922.4]
  assign regs_300_reset = io_reset; // @[:@45923.4 RegFile.scala 76:16:@45930.4]
  assign regs_300_io_in = 64'h0; // @[RegFile.scala 75:16:@45929.4]
  assign regs_300_io_reset = reset; // @[RegFile.scala 78:19:@45933.4]
  assign regs_300_io_enable = 1'h1; // @[RegFile.scala 74:20:@45927.4]
  assign regs_301_clock = clock; // @[:@45936.4]
  assign regs_301_reset = io_reset; // @[:@45937.4 RegFile.scala 76:16:@45944.4]
  assign regs_301_io_in = 64'h0; // @[RegFile.scala 75:16:@45943.4]
  assign regs_301_io_reset = reset; // @[RegFile.scala 78:19:@45947.4]
  assign regs_301_io_enable = 1'h1; // @[RegFile.scala 74:20:@45941.4]
  assign regs_302_clock = clock; // @[:@45950.4]
  assign regs_302_reset = io_reset; // @[:@45951.4 RegFile.scala 76:16:@45958.4]
  assign regs_302_io_in = 64'h0; // @[RegFile.scala 75:16:@45957.4]
  assign regs_302_io_reset = reset; // @[RegFile.scala 78:19:@45961.4]
  assign regs_302_io_enable = 1'h1; // @[RegFile.scala 74:20:@45955.4]
  assign regs_303_clock = clock; // @[:@45964.4]
  assign regs_303_reset = io_reset; // @[:@45965.4 RegFile.scala 76:16:@45972.4]
  assign regs_303_io_in = 64'h0; // @[RegFile.scala 75:16:@45971.4]
  assign regs_303_io_reset = reset; // @[RegFile.scala 78:19:@45975.4]
  assign regs_303_io_enable = 1'h1; // @[RegFile.scala 74:20:@45969.4]
  assign regs_304_clock = clock; // @[:@45978.4]
  assign regs_304_reset = io_reset; // @[:@45979.4 RegFile.scala 76:16:@45986.4]
  assign regs_304_io_in = 64'h0; // @[RegFile.scala 75:16:@45985.4]
  assign regs_304_io_reset = reset; // @[RegFile.scala 78:19:@45989.4]
  assign regs_304_io_enable = 1'h1; // @[RegFile.scala 74:20:@45983.4]
  assign regs_305_clock = clock; // @[:@45992.4]
  assign regs_305_reset = io_reset; // @[:@45993.4 RegFile.scala 76:16:@46000.4]
  assign regs_305_io_in = 64'h0; // @[RegFile.scala 75:16:@45999.4]
  assign regs_305_io_reset = reset; // @[RegFile.scala 78:19:@46003.4]
  assign regs_305_io_enable = 1'h1; // @[RegFile.scala 74:20:@45997.4]
  assign regs_306_clock = clock; // @[:@46006.4]
  assign regs_306_reset = io_reset; // @[:@46007.4 RegFile.scala 76:16:@46014.4]
  assign regs_306_io_in = 64'h0; // @[RegFile.scala 75:16:@46013.4]
  assign regs_306_io_reset = reset; // @[RegFile.scala 78:19:@46017.4]
  assign regs_306_io_enable = 1'h1; // @[RegFile.scala 74:20:@46011.4]
  assign regs_307_clock = clock; // @[:@46020.4]
  assign regs_307_reset = io_reset; // @[:@46021.4 RegFile.scala 76:16:@46028.4]
  assign regs_307_io_in = 64'h0; // @[RegFile.scala 75:16:@46027.4]
  assign regs_307_io_reset = reset; // @[RegFile.scala 78:19:@46031.4]
  assign regs_307_io_enable = 1'h1; // @[RegFile.scala 74:20:@46025.4]
  assign regs_308_clock = clock; // @[:@46034.4]
  assign regs_308_reset = io_reset; // @[:@46035.4 RegFile.scala 76:16:@46042.4]
  assign regs_308_io_in = 64'h0; // @[RegFile.scala 75:16:@46041.4]
  assign regs_308_io_reset = reset; // @[RegFile.scala 78:19:@46045.4]
  assign regs_308_io_enable = 1'h1; // @[RegFile.scala 74:20:@46039.4]
  assign regs_309_clock = clock; // @[:@46048.4]
  assign regs_309_reset = io_reset; // @[:@46049.4 RegFile.scala 76:16:@46056.4]
  assign regs_309_io_in = 64'h0; // @[RegFile.scala 75:16:@46055.4]
  assign regs_309_io_reset = reset; // @[RegFile.scala 78:19:@46059.4]
  assign regs_309_io_enable = 1'h1; // @[RegFile.scala 74:20:@46053.4]
  assign regs_310_clock = clock; // @[:@46062.4]
  assign regs_310_reset = io_reset; // @[:@46063.4 RegFile.scala 76:16:@46070.4]
  assign regs_310_io_in = 64'h0; // @[RegFile.scala 75:16:@46069.4]
  assign regs_310_io_reset = reset; // @[RegFile.scala 78:19:@46073.4]
  assign regs_310_io_enable = 1'h1; // @[RegFile.scala 74:20:@46067.4]
  assign regs_311_clock = clock; // @[:@46076.4]
  assign regs_311_reset = io_reset; // @[:@46077.4 RegFile.scala 76:16:@46084.4]
  assign regs_311_io_in = 64'h0; // @[RegFile.scala 75:16:@46083.4]
  assign regs_311_io_reset = reset; // @[RegFile.scala 78:19:@46087.4]
  assign regs_311_io_enable = 1'h1; // @[RegFile.scala 74:20:@46081.4]
  assign regs_312_clock = clock; // @[:@46090.4]
  assign regs_312_reset = io_reset; // @[:@46091.4 RegFile.scala 76:16:@46098.4]
  assign regs_312_io_in = 64'h0; // @[RegFile.scala 75:16:@46097.4]
  assign regs_312_io_reset = reset; // @[RegFile.scala 78:19:@46101.4]
  assign regs_312_io_enable = 1'h1; // @[RegFile.scala 74:20:@46095.4]
  assign regs_313_clock = clock; // @[:@46104.4]
  assign regs_313_reset = io_reset; // @[:@46105.4 RegFile.scala 76:16:@46112.4]
  assign regs_313_io_in = 64'h0; // @[RegFile.scala 75:16:@46111.4]
  assign regs_313_io_reset = reset; // @[RegFile.scala 78:19:@46115.4]
  assign regs_313_io_enable = 1'h1; // @[RegFile.scala 74:20:@46109.4]
  assign regs_314_clock = clock; // @[:@46118.4]
  assign regs_314_reset = io_reset; // @[:@46119.4 RegFile.scala 76:16:@46126.4]
  assign regs_314_io_in = 64'h0; // @[RegFile.scala 75:16:@46125.4]
  assign regs_314_io_reset = reset; // @[RegFile.scala 78:19:@46129.4]
  assign regs_314_io_enable = 1'h1; // @[RegFile.scala 74:20:@46123.4]
  assign regs_315_clock = clock; // @[:@46132.4]
  assign regs_315_reset = io_reset; // @[:@46133.4 RegFile.scala 76:16:@46140.4]
  assign regs_315_io_in = 64'h0; // @[RegFile.scala 75:16:@46139.4]
  assign regs_315_io_reset = reset; // @[RegFile.scala 78:19:@46143.4]
  assign regs_315_io_enable = 1'h1; // @[RegFile.scala 74:20:@46137.4]
  assign regs_316_clock = clock; // @[:@46146.4]
  assign regs_316_reset = io_reset; // @[:@46147.4 RegFile.scala 76:16:@46154.4]
  assign regs_316_io_in = 64'h0; // @[RegFile.scala 75:16:@46153.4]
  assign regs_316_io_reset = reset; // @[RegFile.scala 78:19:@46157.4]
  assign regs_316_io_enable = 1'h1; // @[RegFile.scala 74:20:@46151.4]
  assign regs_317_clock = clock; // @[:@46160.4]
  assign regs_317_reset = io_reset; // @[:@46161.4 RegFile.scala 76:16:@46168.4]
  assign regs_317_io_in = 64'h0; // @[RegFile.scala 75:16:@46167.4]
  assign regs_317_io_reset = reset; // @[RegFile.scala 78:19:@46171.4]
  assign regs_317_io_enable = 1'h1; // @[RegFile.scala 74:20:@46165.4]
  assign regs_318_clock = clock; // @[:@46174.4]
  assign regs_318_reset = io_reset; // @[:@46175.4 RegFile.scala 76:16:@46182.4]
  assign regs_318_io_in = 64'h0; // @[RegFile.scala 75:16:@46181.4]
  assign regs_318_io_reset = reset; // @[RegFile.scala 78:19:@46185.4]
  assign regs_318_io_enable = 1'h1; // @[RegFile.scala 74:20:@46179.4]
  assign regs_319_clock = clock; // @[:@46188.4]
  assign regs_319_reset = io_reset; // @[:@46189.4 RegFile.scala 76:16:@46196.4]
  assign regs_319_io_in = 64'h0; // @[RegFile.scala 75:16:@46195.4]
  assign regs_319_io_reset = reset; // @[RegFile.scala 78:19:@46199.4]
  assign regs_319_io_enable = 1'h1; // @[RegFile.scala 74:20:@46193.4]
  assign regs_320_clock = clock; // @[:@46202.4]
  assign regs_320_reset = io_reset; // @[:@46203.4 RegFile.scala 76:16:@46210.4]
  assign regs_320_io_in = 64'h0; // @[RegFile.scala 75:16:@46209.4]
  assign regs_320_io_reset = reset; // @[RegFile.scala 78:19:@46213.4]
  assign regs_320_io_enable = 1'h1; // @[RegFile.scala 74:20:@46207.4]
  assign regs_321_clock = clock; // @[:@46216.4]
  assign regs_321_reset = io_reset; // @[:@46217.4 RegFile.scala 76:16:@46224.4]
  assign regs_321_io_in = 64'h0; // @[RegFile.scala 75:16:@46223.4]
  assign regs_321_io_reset = reset; // @[RegFile.scala 78:19:@46227.4]
  assign regs_321_io_enable = 1'h1; // @[RegFile.scala 74:20:@46221.4]
  assign regs_322_clock = clock; // @[:@46230.4]
  assign regs_322_reset = io_reset; // @[:@46231.4 RegFile.scala 76:16:@46238.4]
  assign regs_322_io_in = 64'h0; // @[RegFile.scala 75:16:@46237.4]
  assign regs_322_io_reset = reset; // @[RegFile.scala 78:19:@46241.4]
  assign regs_322_io_enable = 1'h1; // @[RegFile.scala 74:20:@46235.4]
  assign regs_323_clock = clock; // @[:@46244.4]
  assign regs_323_reset = io_reset; // @[:@46245.4 RegFile.scala 76:16:@46252.4]
  assign regs_323_io_in = 64'h0; // @[RegFile.scala 75:16:@46251.4]
  assign regs_323_io_reset = reset; // @[RegFile.scala 78:19:@46255.4]
  assign regs_323_io_enable = 1'h1; // @[RegFile.scala 74:20:@46249.4]
  assign regs_324_clock = clock; // @[:@46258.4]
  assign regs_324_reset = io_reset; // @[:@46259.4 RegFile.scala 76:16:@46266.4]
  assign regs_324_io_in = 64'h0; // @[RegFile.scala 75:16:@46265.4]
  assign regs_324_io_reset = reset; // @[RegFile.scala 78:19:@46269.4]
  assign regs_324_io_enable = 1'h1; // @[RegFile.scala 74:20:@46263.4]
  assign regs_325_clock = clock; // @[:@46272.4]
  assign regs_325_reset = io_reset; // @[:@46273.4 RegFile.scala 76:16:@46280.4]
  assign regs_325_io_in = 64'h0; // @[RegFile.scala 75:16:@46279.4]
  assign regs_325_io_reset = reset; // @[RegFile.scala 78:19:@46283.4]
  assign regs_325_io_enable = 1'h1; // @[RegFile.scala 74:20:@46277.4]
  assign regs_326_clock = clock; // @[:@46286.4]
  assign regs_326_reset = io_reset; // @[:@46287.4 RegFile.scala 76:16:@46294.4]
  assign regs_326_io_in = 64'h0; // @[RegFile.scala 75:16:@46293.4]
  assign regs_326_io_reset = reset; // @[RegFile.scala 78:19:@46297.4]
  assign regs_326_io_enable = 1'h1; // @[RegFile.scala 74:20:@46291.4]
  assign regs_327_clock = clock; // @[:@46300.4]
  assign regs_327_reset = io_reset; // @[:@46301.4 RegFile.scala 76:16:@46308.4]
  assign regs_327_io_in = 64'h0; // @[RegFile.scala 75:16:@46307.4]
  assign regs_327_io_reset = reset; // @[RegFile.scala 78:19:@46311.4]
  assign regs_327_io_enable = 1'h1; // @[RegFile.scala 74:20:@46305.4]
  assign regs_328_clock = clock; // @[:@46314.4]
  assign regs_328_reset = io_reset; // @[:@46315.4 RegFile.scala 76:16:@46322.4]
  assign regs_328_io_in = 64'h0; // @[RegFile.scala 75:16:@46321.4]
  assign regs_328_io_reset = reset; // @[RegFile.scala 78:19:@46325.4]
  assign regs_328_io_enable = 1'h1; // @[RegFile.scala 74:20:@46319.4]
  assign regs_329_clock = clock; // @[:@46328.4]
  assign regs_329_reset = io_reset; // @[:@46329.4 RegFile.scala 76:16:@46336.4]
  assign regs_329_io_in = 64'h0; // @[RegFile.scala 75:16:@46335.4]
  assign regs_329_io_reset = reset; // @[RegFile.scala 78:19:@46339.4]
  assign regs_329_io_enable = 1'h1; // @[RegFile.scala 74:20:@46333.4]
  assign regs_330_clock = clock; // @[:@46342.4]
  assign regs_330_reset = io_reset; // @[:@46343.4 RegFile.scala 76:16:@46350.4]
  assign regs_330_io_in = 64'h0; // @[RegFile.scala 75:16:@46349.4]
  assign regs_330_io_reset = reset; // @[RegFile.scala 78:19:@46353.4]
  assign regs_330_io_enable = 1'h1; // @[RegFile.scala 74:20:@46347.4]
  assign regs_331_clock = clock; // @[:@46356.4]
  assign regs_331_reset = io_reset; // @[:@46357.4 RegFile.scala 76:16:@46364.4]
  assign regs_331_io_in = 64'h0; // @[RegFile.scala 75:16:@46363.4]
  assign regs_331_io_reset = reset; // @[RegFile.scala 78:19:@46367.4]
  assign regs_331_io_enable = 1'h1; // @[RegFile.scala 74:20:@46361.4]
  assign regs_332_clock = clock; // @[:@46370.4]
  assign regs_332_reset = io_reset; // @[:@46371.4 RegFile.scala 76:16:@46378.4]
  assign regs_332_io_in = 64'h0; // @[RegFile.scala 75:16:@46377.4]
  assign regs_332_io_reset = reset; // @[RegFile.scala 78:19:@46381.4]
  assign regs_332_io_enable = 1'h1; // @[RegFile.scala 74:20:@46375.4]
  assign regs_333_clock = clock; // @[:@46384.4]
  assign regs_333_reset = io_reset; // @[:@46385.4 RegFile.scala 76:16:@46392.4]
  assign regs_333_io_in = 64'h0; // @[RegFile.scala 75:16:@46391.4]
  assign regs_333_io_reset = reset; // @[RegFile.scala 78:19:@46395.4]
  assign regs_333_io_enable = 1'h1; // @[RegFile.scala 74:20:@46389.4]
  assign regs_334_clock = clock; // @[:@46398.4]
  assign regs_334_reset = io_reset; // @[:@46399.4 RegFile.scala 76:16:@46406.4]
  assign regs_334_io_in = 64'h0; // @[RegFile.scala 75:16:@46405.4]
  assign regs_334_io_reset = reset; // @[RegFile.scala 78:19:@46409.4]
  assign regs_334_io_enable = 1'h1; // @[RegFile.scala 74:20:@46403.4]
  assign regs_335_clock = clock; // @[:@46412.4]
  assign regs_335_reset = io_reset; // @[:@46413.4 RegFile.scala 76:16:@46420.4]
  assign regs_335_io_in = 64'h0; // @[RegFile.scala 75:16:@46419.4]
  assign regs_335_io_reset = reset; // @[RegFile.scala 78:19:@46423.4]
  assign regs_335_io_enable = 1'h1; // @[RegFile.scala 74:20:@46417.4]
  assign regs_336_clock = clock; // @[:@46426.4]
  assign regs_336_reset = io_reset; // @[:@46427.4 RegFile.scala 76:16:@46434.4]
  assign regs_336_io_in = 64'h0; // @[RegFile.scala 75:16:@46433.4]
  assign regs_336_io_reset = reset; // @[RegFile.scala 78:19:@46437.4]
  assign regs_336_io_enable = 1'h1; // @[RegFile.scala 74:20:@46431.4]
  assign regs_337_clock = clock; // @[:@46440.4]
  assign regs_337_reset = io_reset; // @[:@46441.4 RegFile.scala 76:16:@46448.4]
  assign regs_337_io_in = 64'h0; // @[RegFile.scala 75:16:@46447.4]
  assign regs_337_io_reset = reset; // @[RegFile.scala 78:19:@46451.4]
  assign regs_337_io_enable = 1'h1; // @[RegFile.scala 74:20:@46445.4]
  assign regs_338_clock = clock; // @[:@46454.4]
  assign regs_338_reset = io_reset; // @[:@46455.4 RegFile.scala 76:16:@46462.4]
  assign regs_338_io_in = 64'h0; // @[RegFile.scala 75:16:@46461.4]
  assign regs_338_io_reset = reset; // @[RegFile.scala 78:19:@46465.4]
  assign regs_338_io_enable = 1'h1; // @[RegFile.scala 74:20:@46459.4]
  assign regs_339_clock = clock; // @[:@46468.4]
  assign regs_339_reset = io_reset; // @[:@46469.4 RegFile.scala 76:16:@46476.4]
  assign regs_339_io_in = 64'h0; // @[RegFile.scala 75:16:@46475.4]
  assign regs_339_io_reset = reset; // @[RegFile.scala 78:19:@46479.4]
  assign regs_339_io_enable = 1'h1; // @[RegFile.scala 74:20:@46473.4]
  assign regs_340_clock = clock; // @[:@46482.4]
  assign regs_340_reset = io_reset; // @[:@46483.4 RegFile.scala 76:16:@46490.4]
  assign regs_340_io_in = 64'h0; // @[RegFile.scala 75:16:@46489.4]
  assign regs_340_io_reset = reset; // @[RegFile.scala 78:19:@46493.4]
  assign regs_340_io_enable = 1'h1; // @[RegFile.scala 74:20:@46487.4]
  assign regs_341_clock = clock; // @[:@46496.4]
  assign regs_341_reset = io_reset; // @[:@46497.4 RegFile.scala 76:16:@46504.4]
  assign regs_341_io_in = 64'h0; // @[RegFile.scala 75:16:@46503.4]
  assign regs_341_io_reset = reset; // @[RegFile.scala 78:19:@46507.4]
  assign regs_341_io_enable = 1'h1; // @[RegFile.scala 74:20:@46501.4]
  assign regs_342_clock = clock; // @[:@46510.4]
  assign regs_342_reset = io_reset; // @[:@46511.4 RegFile.scala 76:16:@46518.4]
  assign regs_342_io_in = 64'h0; // @[RegFile.scala 75:16:@46517.4]
  assign regs_342_io_reset = reset; // @[RegFile.scala 78:19:@46521.4]
  assign regs_342_io_enable = 1'h1; // @[RegFile.scala 74:20:@46515.4]
  assign regs_343_clock = clock; // @[:@46524.4]
  assign regs_343_reset = io_reset; // @[:@46525.4 RegFile.scala 76:16:@46532.4]
  assign regs_343_io_in = 64'h0; // @[RegFile.scala 75:16:@46531.4]
  assign regs_343_io_reset = reset; // @[RegFile.scala 78:19:@46535.4]
  assign regs_343_io_enable = 1'h1; // @[RegFile.scala 74:20:@46529.4]
  assign regs_344_clock = clock; // @[:@46538.4]
  assign regs_344_reset = io_reset; // @[:@46539.4 RegFile.scala 76:16:@46546.4]
  assign regs_344_io_in = 64'h0; // @[RegFile.scala 75:16:@46545.4]
  assign regs_344_io_reset = reset; // @[RegFile.scala 78:19:@46549.4]
  assign regs_344_io_enable = 1'h1; // @[RegFile.scala 74:20:@46543.4]
  assign regs_345_clock = clock; // @[:@46552.4]
  assign regs_345_reset = io_reset; // @[:@46553.4 RegFile.scala 76:16:@46560.4]
  assign regs_345_io_in = 64'h0; // @[RegFile.scala 75:16:@46559.4]
  assign regs_345_io_reset = reset; // @[RegFile.scala 78:19:@46563.4]
  assign regs_345_io_enable = 1'h1; // @[RegFile.scala 74:20:@46557.4]
  assign regs_346_clock = clock; // @[:@46566.4]
  assign regs_346_reset = io_reset; // @[:@46567.4 RegFile.scala 76:16:@46574.4]
  assign regs_346_io_in = 64'h0; // @[RegFile.scala 75:16:@46573.4]
  assign regs_346_io_reset = reset; // @[RegFile.scala 78:19:@46577.4]
  assign regs_346_io_enable = 1'h1; // @[RegFile.scala 74:20:@46571.4]
  assign regs_347_clock = clock; // @[:@46580.4]
  assign regs_347_reset = io_reset; // @[:@46581.4 RegFile.scala 76:16:@46588.4]
  assign regs_347_io_in = 64'h0; // @[RegFile.scala 75:16:@46587.4]
  assign regs_347_io_reset = reset; // @[RegFile.scala 78:19:@46591.4]
  assign regs_347_io_enable = 1'h1; // @[RegFile.scala 74:20:@46585.4]
  assign regs_348_clock = clock; // @[:@46594.4]
  assign regs_348_reset = io_reset; // @[:@46595.4 RegFile.scala 76:16:@46602.4]
  assign regs_348_io_in = 64'h0; // @[RegFile.scala 75:16:@46601.4]
  assign regs_348_io_reset = reset; // @[RegFile.scala 78:19:@46605.4]
  assign regs_348_io_enable = 1'h1; // @[RegFile.scala 74:20:@46599.4]
  assign regs_349_clock = clock; // @[:@46608.4]
  assign regs_349_reset = io_reset; // @[:@46609.4 RegFile.scala 76:16:@46616.4]
  assign regs_349_io_in = 64'h0; // @[RegFile.scala 75:16:@46615.4]
  assign regs_349_io_reset = reset; // @[RegFile.scala 78:19:@46619.4]
  assign regs_349_io_enable = 1'h1; // @[RegFile.scala 74:20:@46613.4]
  assign regs_350_clock = clock; // @[:@46622.4]
  assign regs_350_reset = io_reset; // @[:@46623.4 RegFile.scala 76:16:@46630.4]
  assign regs_350_io_in = 64'h0; // @[RegFile.scala 75:16:@46629.4]
  assign regs_350_io_reset = reset; // @[RegFile.scala 78:19:@46633.4]
  assign regs_350_io_enable = 1'h1; // @[RegFile.scala 74:20:@46627.4]
  assign regs_351_clock = clock; // @[:@46636.4]
  assign regs_351_reset = io_reset; // @[:@46637.4 RegFile.scala 76:16:@46644.4]
  assign regs_351_io_in = 64'h0; // @[RegFile.scala 75:16:@46643.4]
  assign regs_351_io_reset = reset; // @[RegFile.scala 78:19:@46647.4]
  assign regs_351_io_enable = 1'h1; // @[RegFile.scala 74:20:@46641.4]
  assign regs_352_clock = clock; // @[:@46650.4]
  assign regs_352_reset = io_reset; // @[:@46651.4 RegFile.scala 76:16:@46658.4]
  assign regs_352_io_in = 64'h0; // @[RegFile.scala 75:16:@46657.4]
  assign regs_352_io_reset = reset; // @[RegFile.scala 78:19:@46661.4]
  assign regs_352_io_enable = 1'h1; // @[RegFile.scala 74:20:@46655.4]
  assign regs_353_clock = clock; // @[:@46664.4]
  assign regs_353_reset = io_reset; // @[:@46665.4 RegFile.scala 76:16:@46672.4]
  assign regs_353_io_in = 64'h0; // @[RegFile.scala 75:16:@46671.4]
  assign regs_353_io_reset = reset; // @[RegFile.scala 78:19:@46675.4]
  assign regs_353_io_enable = 1'h1; // @[RegFile.scala 74:20:@46669.4]
  assign regs_354_clock = clock; // @[:@46678.4]
  assign regs_354_reset = io_reset; // @[:@46679.4 RegFile.scala 76:16:@46686.4]
  assign regs_354_io_in = 64'h0; // @[RegFile.scala 75:16:@46685.4]
  assign regs_354_io_reset = reset; // @[RegFile.scala 78:19:@46689.4]
  assign regs_354_io_enable = 1'h1; // @[RegFile.scala 74:20:@46683.4]
  assign regs_355_clock = clock; // @[:@46692.4]
  assign regs_355_reset = io_reset; // @[:@46693.4 RegFile.scala 76:16:@46700.4]
  assign regs_355_io_in = 64'h0; // @[RegFile.scala 75:16:@46699.4]
  assign regs_355_io_reset = reset; // @[RegFile.scala 78:19:@46703.4]
  assign regs_355_io_enable = 1'h1; // @[RegFile.scala 74:20:@46697.4]
  assign regs_356_clock = clock; // @[:@46706.4]
  assign regs_356_reset = io_reset; // @[:@46707.4 RegFile.scala 76:16:@46714.4]
  assign regs_356_io_in = 64'h0; // @[RegFile.scala 75:16:@46713.4]
  assign regs_356_io_reset = reset; // @[RegFile.scala 78:19:@46717.4]
  assign regs_356_io_enable = 1'h1; // @[RegFile.scala 74:20:@46711.4]
  assign regs_357_clock = clock; // @[:@46720.4]
  assign regs_357_reset = io_reset; // @[:@46721.4 RegFile.scala 76:16:@46728.4]
  assign regs_357_io_in = 64'h0; // @[RegFile.scala 75:16:@46727.4]
  assign regs_357_io_reset = reset; // @[RegFile.scala 78:19:@46731.4]
  assign regs_357_io_enable = 1'h1; // @[RegFile.scala 74:20:@46725.4]
  assign regs_358_clock = clock; // @[:@46734.4]
  assign regs_358_reset = io_reset; // @[:@46735.4 RegFile.scala 76:16:@46742.4]
  assign regs_358_io_in = 64'h0; // @[RegFile.scala 75:16:@46741.4]
  assign regs_358_io_reset = reset; // @[RegFile.scala 78:19:@46745.4]
  assign regs_358_io_enable = 1'h1; // @[RegFile.scala 74:20:@46739.4]
  assign regs_359_clock = clock; // @[:@46748.4]
  assign regs_359_reset = io_reset; // @[:@46749.4 RegFile.scala 76:16:@46756.4]
  assign regs_359_io_in = 64'h0; // @[RegFile.scala 75:16:@46755.4]
  assign regs_359_io_reset = reset; // @[RegFile.scala 78:19:@46759.4]
  assign regs_359_io_enable = 1'h1; // @[RegFile.scala 74:20:@46753.4]
  assign regs_360_clock = clock; // @[:@46762.4]
  assign regs_360_reset = io_reset; // @[:@46763.4 RegFile.scala 76:16:@46770.4]
  assign regs_360_io_in = 64'h0; // @[RegFile.scala 75:16:@46769.4]
  assign regs_360_io_reset = reset; // @[RegFile.scala 78:19:@46773.4]
  assign regs_360_io_enable = 1'h1; // @[RegFile.scala 74:20:@46767.4]
  assign regs_361_clock = clock; // @[:@46776.4]
  assign regs_361_reset = io_reset; // @[:@46777.4 RegFile.scala 76:16:@46784.4]
  assign regs_361_io_in = 64'h0; // @[RegFile.scala 75:16:@46783.4]
  assign regs_361_io_reset = reset; // @[RegFile.scala 78:19:@46787.4]
  assign regs_361_io_enable = 1'h1; // @[RegFile.scala 74:20:@46781.4]
  assign regs_362_clock = clock; // @[:@46790.4]
  assign regs_362_reset = io_reset; // @[:@46791.4 RegFile.scala 76:16:@46798.4]
  assign regs_362_io_in = 64'h0; // @[RegFile.scala 75:16:@46797.4]
  assign regs_362_io_reset = reset; // @[RegFile.scala 78:19:@46801.4]
  assign regs_362_io_enable = 1'h1; // @[RegFile.scala 74:20:@46795.4]
  assign regs_363_clock = clock; // @[:@46804.4]
  assign regs_363_reset = io_reset; // @[:@46805.4 RegFile.scala 76:16:@46812.4]
  assign regs_363_io_in = 64'h0; // @[RegFile.scala 75:16:@46811.4]
  assign regs_363_io_reset = reset; // @[RegFile.scala 78:19:@46815.4]
  assign regs_363_io_enable = 1'h1; // @[RegFile.scala 74:20:@46809.4]
  assign regs_364_clock = clock; // @[:@46818.4]
  assign regs_364_reset = io_reset; // @[:@46819.4 RegFile.scala 76:16:@46826.4]
  assign regs_364_io_in = 64'h0; // @[RegFile.scala 75:16:@46825.4]
  assign regs_364_io_reset = reset; // @[RegFile.scala 78:19:@46829.4]
  assign regs_364_io_enable = 1'h1; // @[RegFile.scala 74:20:@46823.4]
  assign regs_365_clock = clock; // @[:@46832.4]
  assign regs_365_reset = io_reset; // @[:@46833.4 RegFile.scala 76:16:@46840.4]
  assign regs_365_io_in = 64'h0; // @[RegFile.scala 75:16:@46839.4]
  assign regs_365_io_reset = reset; // @[RegFile.scala 78:19:@46843.4]
  assign regs_365_io_enable = 1'h1; // @[RegFile.scala 74:20:@46837.4]
  assign regs_366_clock = clock; // @[:@46846.4]
  assign regs_366_reset = io_reset; // @[:@46847.4 RegFile.scala 76:16:@46854.4]
  assign regs_366_io_in = 64'h0; // @[RegFile.scala 75:16:@46853.4]
  assign regs_366_io_reset = reset; // @[RegFile.scala 78:19:@46857.4]
  assign regs_366_io_enable = 1'h1; // @[RegFile.scala 74:20:@46851.4]
  assign regs_367_clock = clock; // @[:@46860.4]
  assign regs_367_reset = io_reset; // @[:@46861.4 RegFile.scala 76:16:@46868.4]
  assign regs_367_io_in = 64'h0; // @[RegFile.scala 75:16:@46867.4]
  assign regs_367_io_reset = reset; // @[RegFile.scala 78:19:@46871.4]
  assign regs_367_io_enable = 1'h1; // @[RegFile.scala 74:20:@46865.4]
  assign regs_368_clock = clock; // @[:@46874.4]
  assign regs_368_reset = io_reset; // @[:@46875.4 RegFile.scala 76:16:@46882.4]
  assign regs_368_io_in = 64'h0; // @[RegFile.scala 75:16:@46881.4]
  assign regs_368_io_reset = reset; // @[RegFile.scala 78:19:@46885.4]
  assign regs_368_io_enable = 1'h1; // @[RegFile.scala 74:20:@46879.4]
  assign regs_369_clock = clock; // @[:@46888.4]
  assign regs_369_reset = io_reset; // @[:@46889.4 RegFile.scala 76:16:@46896.4]
  assign regs_369_io_in = 64'h0; // @[RegFile.scala 75:16:@46895.4]
  assign regs_369_io_reset = reset; // @[RegFile.scala 78:19:@46899.4]
  assign regs_369_io_enable = 1'h1; // @[RegFile.scala 74:20:@46893.4]
  assign regs_370_clock = clock; // @[:@46902.4]
  assign regs_370_reset = io_reset; // @[:@46903.4 RegFile.scala 76:16:@46910.4]
  assign regs_370_io_in = 64'h0; // @[RegFile.scala 75:16:@46909.4]
  assign regs_370_io_reset = reset; // @[RegFile.scala 78:19:@46913.4]
  assign regs_370_io_enable = 1'h1; // @[RegFile.scala 74:20:@46907.4]
  assign regs_371_clock = clock; // @[:@46916.4]
  assign regs_371_reset = io_reset; // @[:@46917.4 RegFile.scala 76:16:@46924.4]
  assign regs_371_io_in = 64'h0; // @[RegFile.scala 75:16:@46923.4]
  assign regs_371_io_reset = reset; // @[RegFile.scala 78:19:@46927.4]
  assign regs_371_io_enable = 1'h1; // @[RegFile.scala 74:20:@46921.4]
  assign regs_372_clock = clock; // @[:@46930.4]
  assign regs_372_reset = io_reset; // @[:@46931.4 RegFile.scala 76:16:@46938.4]
  assign regs_372_io_in = 64'h0; // @[RegFile.scala 75:16:@46937.4]
  assign regs_372_io_reset = reset; // @[RegFile.scala 78:19:@46941.4]
  assign regs_372_io_enable = 1'h1; // @[RegFile.scala 74:20:@46935.4]
  assign regs_373_clock = clock; // @[:@46944.4]
  assign regs_373_reset = io_reset; // @[:@46945.4 RegFile.scala 76:16:@46952.4]
  assign regs_373_io_in = 64'h0; // @[RegFile.scala 75:16:@46951.4]
  assign regs_373_io_reset = reset; // @[RegFile.scala 78:19:@46955.4]
  assign regs_373_io_enable = 1'h1; // @[RegFile.scala 74:20:@46949.4]
  assign regs_374_clock = clock; // @[:@46958.4]
  assign regs_374_reset = io_reset; // @[:@46959.4 RegFile.scala 76:16:@46966.4]
  assign regs_374_io_in = 64'h0; // @[RegFile.scala 75:16:@46965.4]
  assign regs_374_io_reset = reset; // @[RegFile.scala 78:19:@46969.4]
  assign regs_374_io_enable = 1'h1; // @[RegFile.scala 74:20:@46963.4]
  assign regs_375_clock = clock; // @[:@46972.4]
  assign regs_375_reset = io_reset; // @[:@46973.4 RegFile.scala 76:16:@46980.4]
  assign regs_375_io_in = 64'h0; // @[RegFile.scala 75:16:@46979.4]
  assign regs_375_io_reset = reset; // @[RegFile.scala 78:19:@46983.4]
  assign regs_375_io_enable = 1'h1; // @[RegFile.scala 74:20:@46977.4]
  assign regs_376_clock = clock; // @[:@46986.4]
  assign regs_376_reset = io_reset; // @[:@46987.4 RegFile.scala 76:16:@46994.4]
  assign regs_376_io_in = 64'h0; // @[RegFile.scala 75:16:@46993.4]
  assign regs_376_io_reset = reset; // @[RegFile.scala 78:19:@46997.4]
  assign regs_376_io_enable = 1'h1; // @[RegFile.scala 74:20:@46991.4]
  assign regs_377_clock = clock; // @[:@47000.4]
  assign regs_377_reset = io_reset; // @[:@47001.4 RegFile.scala 76:16:@47008.4]
  assign regs_377_io_in = 64'h0; // @[RegFile.scala 75:16:@47007.4]
  assign regs_377_io_reset = reset; // @[RegFile.scala 78:19:@47011.4]
  assign regs_377_io_enable = 1'h1; // @[RegFile.scala 74:20:@47005.4]
  assign regs_378_clock = clock; // @[:@47014.4]
  assign regs_378_reset = io_reset; // @[:@47015.4 RegFile.scala 76:16:@47022.4]
  assign regs_378_io_in = 64'h0; // @[RegFile.scala 75:16:@47021.4]
  assign regs_378_io_reset = reset; // @[RegFile.scala 78:19:@47025.4]
  assign regs_378_io_enable = 1'h1; // @[RegFile.scala 74:20:@47019.4]
  assign regs_379_clock = clock; // @[:@47028.4]
  assign regs_379_reset = io_reset; // @[:@47029.4 RegFile.scala 76:16:@47036.4]
  assign regs_379_io_in = 64'h0; // @[RegFile.scala 75:16:@47035.4]
  assign regs_379_io_reset = reset; // @[RegFile.scala 78:19:@47039.4]
  assign regs_379_io_enable = 1'h1; // @[RegFile.scala 74:20:@47033.4]
  assign regs_380_clock = clock; // @[:@47042.4]
  assign regs_380_reset = io_reset; // @[:@47043.4 RegFile.scala 76:16:@47050.4]
  assign regs_380_io_in = 64'h0; // @[RegFile.scala 75:16:@47049.4]
  assign regs_380_io_reset = reset; // @[RegFile.scala 78:19:@47053.4]
  assign regs_380_io_enable = 1'h1; // @[RegFile.scala 74:20:@47047.4]
  assign regs_381_clock = clock; // @[:@47056.4]
  assign regs_381_reset = io_reset; // @[:@47057.4 RegFile.scala 76:16:@47064.4]
  assign regs_381_io_in = 64'h0; // @[RegFile.scala 75:16:@47063.4]
  assign regs_381_io_reset = reset; // @[RegFile.scala 78:19:@47067.4]
  assign regs_381_io_enable = 1'h1; // @[RegFile.scala 74:20:@47061.4]
  assign regs_382_clock = clock; // @[:@47070.4]
  assign regs_382_reset = io_reset; // @[:@47071.4 RegFile.scala 76:16:@47078.4]
  assign regs_382_io_in = 64'h0; // @[RegFile.scala 75:16:@47077.4]
  assign regs_382_io_reset = reset; // @[RegFile.scala 78:19:@47081.4]
  assign regs_382_io_enable = 1'h1; // @[RegFile.scala 74:20:@47075.4]
  assign regs_383_clock = clock; // @[:@47084.4]
  assign regs_383_reset = io_reset; // @[:@47085.4 RegFile.scala 76:16:@47092.4]
  assign regs_383_io_in = 64'h0; // @[RegFile.scala 75:16:@47091.4]
  assign regs_383_io_reset = reset; // @[RegFile.scala 78:19:@47095.4]
  assign regs_383_io_enable = 1'h1; // @[RegFile.scala 74:20:@47089.4]
  assign regs_384_clock = clock; // @[:@47098.4]
  assign regs_384_reset = io_reset; // @[:@47099.4 RegFile.scala 76:16:@47106.4]
  assign regs_384_io_in = 64'h0; // @[RegFile.scala 75:16:@47105.4]
  assign regs_384_io_reset = reset; // @[RegFile.scala 78:19:@47109.4]
  assign regs_384_io_enable = 1'h1; // @[RegFile.scala 74:20:@47103.4]
  assign regs_385_clock = clock; // @[:@47112.4]
  assign regs_385_reset = io_reset; // @[:@47113.4 RegFile.scala 76:16:@47120.4]
  assign regs_385_io_in = 64'h0; // @[RegFile.scala 75:16:@47119.4]
  assign regs_385_io_reset = reset; // @[RegFile.scala 78:19:@47123.4]
  assign regs_385_io_enable = 1'h1; // @[RegFile.scala 74:20:@47117.4]
  assign regs_386_clock = clock; // @[:@47126.4]
  assign regs_386_reset = io_reset; // @[:@47127.4 RegFile.scala 76:16:@47134.4]
  assign regs_386_io_in = 64'h0; // @[RegFile.scala 75:16:@47133.4]
  assign regs_386_io_reset = reset; // @[RegFile.scala 78:19:@47137.4]
  assign regs_386_io_enable = 1'h1; // @[RegFile.scala 74:20:@47131.4]
  assign regs_387_clock = clock; // @[:@47140.4]
  assign regs_387_reset = io_reset; // @[:@47141.4 RegFile.scala 76:16:@47148.4]
  assign regs_387_io_in = 64'h0; // @[RegFile.scala 75:16:@47147.4]
  assign regs_387_io_reset = reset; // @[RegFile.scala 78:19:@47151.4]
  assign regs_387_io_enable = 1'h1; // @[RegFile.scala 74:20:@47145.4]
  assign regs_388_clock = clock; // @[:@47154.4]
  assign regs_388_reset = io_reset; // @[:@47155.4 RegFile.scala 76:16:@47162.4]
  assign regs_388_io_in = 64'h0; // @[RegFile.scala 75:16:@47161.4]
  assign regs_388_io_reset = reset; // @[RegFile.scala 78:19:@47165.4]
  assign regs_388_io_enable = 1'h1; // @[RegFile.scala 74:20:@47159.4]
  assign regs_389_clock = clock; // @[:@47168.4]
  assign regs_389_reset = io_reset; // @[:@47169.4 RegFile.scala 76:16:@47176.4]
  assign regs_389_io_in = 64'h0; // @[RegFile.scala 75:16:@47175.4]
  assign regs_389_io_reset = reset; // @[RegFile.scala 78:19:@47179.4]
  assign regs_389_io_enable = 1'h1; // @[RegFile.scala 74:20:@47173.4]
  assign regs_390_clock = clock; // @[:@47182.4]
  assign regs_390_reset = io_reset; // @[:@47183.4 RegFile.scala 76:16:@47190.4]
  assign regs_390_io_in = 64'h0; // @[RegFile.scala 75:16:@47189.4]
  assign regs_390_io_reset = reset; // @[RegFile.scala 78:19:@47193.4]
  assign regs_390_io_enable = 1'h1; // @[RegFile.scala 74:20:@47187.4]
  assign regs_391_clock = clock; // @[:@47196.4]
  assign regs_391_reset = io_reset; // @[:@47197.4 RegFile.scala 76:16:@47204.4]
  assign regs_391_io_in = 64'h0; // @[RegFile.scala 75:16:@47203.4]
  assign regs_391_io_reset = reset; // @[RegFile.scala 78:19:@47207.4]
  assign regs_391_io_enable = 1'h1; // @[RegFile.scala 74:20:@47201.4]
  assign regs_392_clock = clock; // @[:@47210.4]
  assign regs_392_reset = io_reset; // @[:@47211.4 RegFile.scala 76:16:@47218.4]
  assign regs_392_io_in = 64'h0; // @[RegFile.scala 75:16:@47217.4]
  assign regs_392_io_reset = reset; // @[RegFile.scala 78:19:@47221.4]
  assign regs_392_io_enable = 1'h1; // @[RegFile.scala 74:20:@47215.4]
  assign regs_393_clock = clock; // @[:@47224.4]
  assign regs_393_reset = io_reset; // @[:@47225.4 RegFile.scala 76:16:@47232.4]
  assign regs_393_io_in = 64'h0; // @[RegFile.scala 75:16:@47231.4]
  assign regs_393_io_reset = reset; // @[RegFile.scala 78:19:@47235.4]
  assign regs_393_io_enable = 1'h1; // @[RegFile.scala 74:20:@47229.4]
  assign regs_394_clock = clock; // @[:@47238.4]
  assign regs_394_reset = io_reset; // @[:@47239.4 RegFile.scala 76:16:@47246.4]
  assign regs_394_io_in = 64'h0; // @[RegFile.scala 75:16:@47245.4]
  assign regs_394_io_reset = reset; // @[RegFile.scala 78:19:@47249.4]
  assign regs_394_io_enable = 1'h1; // @[RegFile.scala 74:20:@47243.4]
  assign regs_395_clock = clock; // @[:@47252.4]
  assign regs_395_reset = io_reset; // @[:@47253.4 RegFile.scala 76:16:@47260.4]
  assign regs_395_io_in = 64'h0; // @[RegFile.scala 75:16:@47259.4]
  assign regs_395_io_reset = reset; // @[RegFile.scala 78:19:@47263.4]
  assign regs_395_io_enable = 1'h1; // @[RegFile.scala 74:20:@47257.4]
  assign regs_396_clock = clock; // @[:@47266.4]
  assign regs_396_reset = io_reset; // @[:@47267.4 RegFile.scala 76:16:@47274.4]
  assign regs_396_io_in = 64'h0; // @[RegFile.scala 75:16:@47273.4]
  assign regs_396_io_reset = reset; // @[RegFile.scala 78:19:@47277.4]
  assign regs_396_io_enable = 1'h1; // @[RegFile.scala 74:20:@47271.4]
  assign regs_397_clock = clock; // @[:@47280.4]
  assign regs_397_reset = io_reset; // @[:@47281.4 RegFile.scala 76:16:@47288.4]
  assign regs_397_io_in = 64'h0; // @[RegFile.scala 75:16:@47287.4]
  assign regs_397_io_reset = reset; // @[RegFile.scala 78:19:@47291.4]
  assign regs_397_io_enable = 1'h1; // @[RegFile.scala 74:20:@47285.4]
  assign regs_398_clock = clock; // @[:@47294.4]
  assign regs_398_reset = io_reset; // @[:@47295.4 RegFile.scala 76:16:@47302.4]
  assign regs_398_io_in = 64'h0; // @[RegFile.scala 75:16:@47301.4]
  assign regs_398_io_reset = reset; // @[RegFile.scala 78:19:@47305.4]
  assign regs_398_io_enable = 1'h1; // @[RegFile.scala 74:20:@47299.4]
  assign regs_399_clock = clock; // @[:@47308.4]
  assign regs_399_reset = io_reset; // @[:@47309.4 RegFile.scala 76:16:@47316.4]
  assign regs_399_io_in = 64'h0; // @[RegFile.scala 75:16:@47315.4]
  assign regs_399_io_reset = reset; // @[RegFile.scala 78:19:@47319.4]
  assign regs_399_io_enable = 1'h1; // @[RegFile.scala 74:20:@47313.4]
  assign regs_400_clock = clock; // @[:@47322.4]
  assign regs_400_reset = io_reset; // @[:@47323.4 RegFile.scala 76:16:@47330.4]
  assign regs_400_io_in = 64'h0; // @[RegFile.scala 75:16:@47329.4]
  assign regs_400_io_reset = reset; // @[RegFile.scala 78:19:@47333.4]
  assign regs_400_io_enable = 1'h1; // @[RegFile.scala 74:20:@47327.4]
  assign regs_401_clock = clock; // @[:@47336.4]
  assign regs_401_reset = io_reset; // @[:@47337.4 RegFile.scala 76:16:@47344.4]
  assign regs_401_io_in = 64'h0; // @[RegFile.scala 75:16:@47343.4]
  assign regs_401_io_reset = reset; // @[RegFile.scala 78:19:@47347.4]
  assign regs_401_io_enable = 1'h1; // @[RegFile.scala 74:20:@47341.4]
  assign regs_402_clock = clock; // @[:@47350.4]
  assign regs_402_reset = io_reset; // @[:@47351.4 RegFile.scala 76:16:@47358.4]
  assign regs_402_io_in = 64'h0; // @[RegFile.scala 75:16:@47357.4]
  assign regs_402_io_reset = reset; // @[RegFile.scala 78:19:@47361.4]
  assign regs_402_io_enable = 1'h1; // @[RegFile.scala 74:20:@47355.4]
  assign regs_403_clock = clock; // @[:@47364.4]
  assign regs_403_reset = io_reset; // @[:@47365.4 RegFile.scala 76:16:@47372.4]
  assign regs_403_io_in = 64'h0; // @[RegFile.scala 75:16:@47371.4]
  assign regs_403_io_reset = reset; // @[RegFile.scala 78:19:@47375.4]
  assign regs_403_io_enable = 1'h1; // @[RegFile.scala 74:20:@47369.4]
  assign regs_404_clock = clock; // @[:@47378.4]
  assign regs_404_reset = io_reset; // @[:@47379.4 RegFile.scala 76:16:@47386.4]
  assign regs_404_io_in = 64'h0; // @[RegFile.scala 75:16:@47385.4]
  assign regs_404_io_reset = reset; // @[RegFile.scala 78:19:@47389.4]
  assign regs_404_io_enable = 1'h1; // @[RegFile.scala 74:20:@47383.4]
  assign regs_405_clock = clock; // @[:@47392.4]
  assign regs_405_reset = io_reset; // @[:@47393.4 RegFile.scala 76:16:@47400.4]
  assign regs_405_io_in = 64'h0; // @[RegFile.scala 75:16:@47399.4]
  assign regs_405_io_reset = reset; // @[RegFile.scala 78:19:@47403.4]
  assign regs_405_io_enable = 1'h1; // @[RegFile.scala 74:20:@47397.4]
  assign regs_406_clock = clock; // @[:@47406.4]
  assign regs_406_reset = io_reset; // @[:@47407.4 RegFile.scala 76:16:@47414.4]
  assign regs_406_io_in = 64'h0; // @[RegFile.scala 75:16:@47413.4]
  assign regs_406_io_reset = reset; // @[RegFile.scala 78:19:@47417.4]
  assign regs_406_io_enable = 1'h1; // @[RegFile.scala 74:20:@47411.4]
  assign regs_407_clock = clock; // @[:@47420.4]
  assign regs_407_reset = io_reset; // @[:@47421.4 RegFile.scala 76:16:@47428.4]
  assign regs_407_io_in = 64'h0; // @[RegFile.scala 75:16:@47427.4]
  assign regs_407_io_reset = reset; // @[RegFile.scala 78:19:@47431.4]
  assign regs_407_io_enable = 1'h1; // @[RegFile.scala 74:20:@47425.4]
  assign regs_408_clock = clock; // @[:@47434.4]
  assign regs_408_reset = io_reset; // @[:@47435.4 RegFile.scala 76:16:@47442.4]
  assign regs_408_io_in = 64'h0; // @[RegFile.scala 75:16:@47441.4]
  assign regs_408_io_reset = reset; // @[RegFile.scala 78:19:@47445.4]
  assign regs_408_io_enable = 1'h1; // @[RegFile.scala 74:20:@47439.4]
  assign regs_409_clock = clock; // @[:@47448.4]
  assign regs_409_reset = io_reset; // @[:@47449.4 RegFile.scala 76:16:@47456.4]
  assign regs_409_io_in = 64'h0; // @[RegFile.scala 75:16:@47455.4]
  assign regs_409_io_reset = reset; // @[RegFile.scala 78:19:@47459.4]
  assign regs_409_io_enable = 1'h1; // @[RegFile.scala 74:20:@47453.4]
  assign regs_410_clock = clock; // @[:@47462.4]
  assign regs_410_reset = io_reset; // @[:@47463.4 RegFile.scala 76:16:@47470.4]
  assign regs_410_io_in = 64'h0; // @[RegFile.scala 75:16:@47469.4]
  assign regs_410_io_reset = reset; // @[RegFile.scala 78:19:@47473.4]
  assign regs_410_io_enable = 1'h1; // @[RegFile.scala 74:20:@47467.4]
  assign regs_411_clock = clock; // @[:@47476.4]
  assign regs_411_reset = io_reset; // @[:@47477.4 RegFile.scala 76:16:@47484.4]
  assign regs_411_io_in = 64'h0; // @[RegFile.scala 75:16:@47483.4]
  assign regs_411_io_reset = reset; // @[RegFile.scala 78:19:@47487.4]
  assign regs_411_io_enable = 1'h1; // @[RegFile.scala 74:20:@47481.4]
  assign regs_412_clock = clock; // @[:@47490.4]
  assign regs_412_reset = io_reset; // @[:@47491.4 RegFile.scala 76:16:@47498.4]
  assign regs_412_io_in = 64'h0; // @[RegFile.scala 75:16:@47497.4]
  assign regs_412_io_reset = reset; // @[RegFile.scala 78:19:@47501.4]
  assign regs_412_io_enable = 1'h1; // @[RegFile.scala 74:20:@47495.4]
  assign regs_413_clock = clock; // @[:@47504.4]
  assign regs_413_reset = io_reset; // @[:@47505.4 RegFile.scala 76:16:@47512.4]
  assign regs_413_io_in = 64'h0; // @[RegFile.scala 75:16:@47511.4]
  assign regs_413_io_reset = reset; // @[RegFile.scala 78:19:@47515.4]
  assign regs_413_io_enable = 1'h1; // @[RegFile.scala 74:20:@47509.4]
  assign regs_414_clock = clock; // @[:@47518.4]
  assign regs_414_reset = io_reset; // @[:@47519.4 RegFile.scala 76:16:@47526.4]
  assign regs_414_io_in = 64'h0; // @[RegFile.scala 75:16:@47525.4]
  assign regs_414_io_reset = reset; // @[RegFile.scala 78:19:@47529.4]
  assign regs_414_io_enable = 1'h1; // @[RegFile.scala 74:20:@47523.4]
  assign regs_415_clock = clock; // @[:@47532.4]
  assign regs_415_reset = io_reset; // @[:@47533.4 RegFile.scala 76:16:@47540.4]
  assign regs_415_io_in = 64'h0; // @[RegFile.scala 75:16:@47539.4]
  assign regs_415_io_reset = reset; // @[RegFile.scala 78:19:@47543.4]
  assign regs_415_io_enable = 1'h1; // @[RegFile.scala 74:20:@47537.4]
  assign regs_416_clock = clock; // @[:@47546.4]
  assign regs_416_reset = io_reset; // @[:@47547.4 RegFile.scala 76:16:@47554.4]
  assign regs_416_io_in = 64'h0; // @[RegFile.scala 75:16:@47553.4]
  assign regs_416_io_reset = reset; // @[RegFile.scala 78:19:@47557.4]
  assign regs_416_io_enable = 1'h1; // @[RegFile.scala 74:20:@47551.4]
  assign regs_417_clock = clock; // @[:@47560.4]
  assign regs_417_reset = io_reset; // @[:@47561.4 RegFile.scala 76:16:@47568.4]
  assign regs_417_io_in = 64'h0; // @[RegFile.scala 75:16:@47567.4]
  assign regs_417_io_reset = reset; // @[RegFile.scala 78:19:@47571.4]
  assign regs_417_io_enable = 1'h1; // @[RegFile.scala 74:20:@47565.4]
  assign regs_418_clock = clock; // @[:@47574.4]
  assign regs_418_reset = io_reset; // @[:@47575.4 RegFile.scala 76:16:@47582.4]
  assign regs_418_io_in = 64'h0; // @[RegFile.scala 75:16:@47581.4]
  assign regs_418_io_reset = reset; // @[RegFile.scala 78:19:@47585.4]
  assign regs_418_io_enable = 1'h1; // @[RegFile.scala 74:20:@47579.4]
  assign regs_419_clock = clock; // @[:@47588.4]
  assign regs_419_reset = io_reset; // @[:@47589.4 RegFile.scala 76:16:@47596.4]
  assign regs_419_io_in = 64'h0; // @[RegFile.scala 75:16:@47595.4]
  assign regs_419_io_reset = reset; // @[RegFile.scala 78:19:@47599.4]
  assign regs_419_io_enable = 1'h1; // @[RegFile.scala 74:20:@47593.4]
  assign regs_420_clock = clock; // @[:@47602.4]
  assign regs_420_reset = io_reset; // @[:@47603.4 RegFile.scala 76:16:@47610.4]
  assign regs_420_io_in = 64'h0; // @[RegFile.scala 75:16:@47609.4]
  assign regs_420_io_reset = reset; // @[RegFile.scala 78:19:@47613.4]
  assign regs_420_io_enable = 1'h1; // @[RegFile.scala 74:20:@47607.4]
  assign regs_421_clock = clock; // @[:@47616.4]
  assign regs_421_reset = io_reset; // @[:@47617.4 RegFile.scala 76:16:@47624.4]
  assign regs_421_io_in = 64'h0; // @[RegFile.scala 75:16:@47623.4]
  assign regs_421_io_reset = reset; // @[RegFile.scala 78:19:@47627.4]
  assign regs_421_io_enable = 1'h1; // @[RegFile.scala 74:20:@47621.4]
  assign regs_422_clock = clock; // @[:@47630.4]
  assign regs_422_reset = io_reset; // @[:@47631.4 RegFile.scala 76:16:@47638.4]
  assign regs_422_io_in = 64'h0; // @[RegFile.scala 75:16:@47637.4]
  assign regs_422_io_reset = reset; // @[RegFile.scala 78:19:@47641.4]
  assign regs_422_io_enable = 1'h1; // @[RegFile.scala 74:20:@47635.4]
  assign regs_423_clock = clock; // @[:@47644.4]
  assign regs_423_reset = io_reset; // @[:@47645.4 RegFile.scala 76:16:@47652.4]
  assign regs_423_io_in = 64'h0; // @[RegFile.scala 75:16:@47651.4]
  assign regs_423_io_reset = reset; // @[RegFile.scala 78:19:@47655.4]
  assign regs_423_io_enable = 1'h1; // @[RegFile.scala 74:20:@47649.4]
  assign regs_424_clock = clock; // @[:@47658.4]
  assign regs_424_reset = io_reset; // @[:@47659.4 RegFile.scala 76:16:@47666.4]
  assign regs_424_io_in = 64'h0; // @[RegFile.scala 75:16:@47665.4]
  assign regs_424_io_reset = reset; // @[RegFile.scala 78:19:@47669.4]
  assign regs_424_io_enable = 1'h1; // @[RegFile.scala 74:20:@47663.4]
  assign regs_425_clock = clock; // @[:@47672.4]
  assign regs_425_reset = io_reset; // @[:@47673.4 RegFile.scala 76:16:@47680.4]
  assign regs_425_io_in = 64'h0; // @[RegFile.scala 75:16:@47679.4]
  assign regs_425_io_reset = reset; // @[RegFile.scala 78:19:@47683.4]
  assign regs_425_io_enable = 1'h1; // @[RegFile.scala 74:20:@47677.4]
  assign regs_426_clock = clock; // @[:@47686.4]
  assign regs_426_reset = io_reset; // @[:@47687.4 RegFile.scala 76:16:@47694.4]
  assign regs_426_io_in = 64'h0; // @[RegFile.scala 75:16:@47693.4]
  assign regs_426_io_reset = reset; // @[RegFile.scala 78:19:@47697.4]
  assign regs_426_io_enable = 1'h1; // @[RegFile.scala 74:20:@47691.4]
  assign regs_427_clock = clock; // @[:@47700.4]
  assign regs_427_reset = io_reset; // @[:@47701.4 RegFile.scala 76:16:@47708.4]
  assign regs_427_io_in = 64'h0; // @[RegFile.scala 75:16:@47707.4]
  assign regs_427_io_reset = reset; // @[RegFile.scala 78:19:@47711.4]
  assign regs_427_io_enable = 1'h1; // @[RegFile.scala 74:20:@47705.4]
  assign regs_428_clock = clock; // @[:@47714.4]
  assign regs_428_reset = io_reset; // @[:@47715.4 RegFile.scala 76:16:@47722.4]
  assign regs_428_io_in = 64'h0; // @[RegFile.scala 75:16:@47721.4]
  assign regs_428_io_reset = reset; // @[RegFile.scala 78:19:@47725.4]
  assign regs_428_io_enable = 1'h1; // @[RegFile.scala 74:20:@47719.4]
  assign regs_429_clock = clock; // @[:@47728.4]
  assign regs_429_reset = io_reset; // @[:@47729.4 RegFile.scala 76:16:@47736.4]
  assign regs_429_io_in = 64'h0; // @[RegFile.scala 75:16:@47735.4]
  assign regs_429_io_reset = reset; // @[RegFile.scala 78:19:@47739.4]
  assign regs_429_io_enable = 1'h1; // @[RegFile.scala 74:20:@47733.4]
  assign regs_430_clock = clock; // @[:@47742.4]
  assign regs_430_reset = io_reset; // @[:@47743.4 RegFile.scala 76:16:@47750.4]
  assign regs_430_io_in = 64'h0; // @[RegFile.scala 75:16:@47749.4]
  assign regs_430_io_reset = reset; // @[RegFile.scala 78:19:@47753.4]
  assign regs_430_io_enable = 1'h1; // @[RegFile.scala 74:20:@47747.4]
  assign regs_431_clock = clock; // @[:@47756.4]
  assign regs_431_reset = io_reset; // @[:@47757.4 RegFile.scala 76:16:@47764.4]
  assign regs_431_io_in = 64'h0; // @[RegFile.scala 75:16:@47763.4]
  assign regs_431_io_reset = reset; // @[RegFile.scala 78:19:@47767.4]
  assign regs_431_io_enable = 1'h1; // @[RegFile.scala 74:20:@47761.4]
  assign regs_432_clock = clock; // @[:@47770.4]
  assign regs_432_reset = io_reset; // @[:@47771.4 RegFile.scala 76:16:@47778.4]
  assign regs_432_io_in = 64'h0; // @[RegFile.scala 75:16:@47777.4]
  assign regs_432_io_reset = reset; // @[RegFile.scala 78:19:@47781.4]
  assign regs_432_io_enable = 1'h1; // @[RegFile.scala 74:20:@47775.4]
  assign regs_433_clock = clock; // @[:@47784.4]
  assign regs_433_reset = io_reset; // @[:@47785.4 RegFile.scala 76:16:@47792.4]
  assign regs_433_io_in = 64'h0; // @[RegFile.scala 75:16:@47791.4]
  assign regs_433_io_reset = reset; // @[RegFile.scala 78:19:@47795.4]
  assign regs_433_io_enable = 1'h1; // @[RegFile.scala 74:20:@47789.4]
  assign regs_434_clock = clock; // @[:@47798.4]
  assign regs_434_reset = io_reset; // @[:@47799.4 RegFile.scala 76:16:@47806.4]
  assign regs_434_io_in = 64'h0; // @[RegFile.scala 75:16:@47805.4]
  assign regs_434_io_reset = reset; // @[RegFile.scala 78:19:@47809.4]
  assign regs_434_io_enable = 1'h1; // @[RegFile.scala 74:20:@47803.4]
  assign regs_435_clock = clock; // @[:@47812.4]
  assign regs_435_reset = io_reset; // @[:@47813.4 RegFile.scala 76:16:@47820.4]
  assign regs_435_io_in = 64'h0; // @[RegFile.scala 75:16:@47819.4]
  assign regs_435_io_reset = reset; // @[RegFile.scala 78:19:@47823.4]
  assign regs_435_io_enable = 1'h1; // @[RegFile.scala 74:20:@47817.4]
  assign regs_436_clock = clock; // @[:@47826.4]
  assign regs_436_reset = io_reset; // @[:@47827.4 RegFile.scala 76:16:@47834.4]
  assign regs_436_io_in = 64'h0; // @[RegFile.scala 75:16:@47833.4]
  assign regs_436_io_reset = reset; // @[RegFile.scala 78:19:@47837.4]
  assign regs_436_io_enable = 1'h1; // @[RegFile.scala 74:20:@47831.4]
  assign regs_437_clock = clock; // @[:@47840.4]
  assign regs_437_reset = io_reset; // @[:@47841.4 RegFile.scala 76:16:@47848.4]
  assign regs_437_io_in = 64'h0; // @[RegFile.scala 75:16:@47847.4]
  assign regs_437_io_reset = reset; // @[RegFile.scala 78:19:@47851.4]
  assign regs_437_io_enable = 1'h1; // @[RegFile.scala 74:20:@47845.4]
  assign regs_438_clock = clock; // @[:@47854.4]
  assign regs_438_reset = io_reset; // @[:@47855.4 RegFile.scala 76:16:@47862.4]
  assign regs_438_io_in = 64'h0; // @[RegFile.scala 75:16:@47861.4]
  assign regs_438_io_reset = reset; // @[RegFile.scala 78:19:@47865.4]
  assign regs_438_io_enable = 1'h1; // @[RegFile.scala 74:20:@47859.4]
  assign regs_439_clock = clock; // @[:@47868.4]
  assign regs_439_reset = io_reset; // @[:@47869.4 RegFile.scala 76:16:@47876.4]
  assign regs_439_io_in = 64'h0; // @[RegFile.scala 75:16:@47875.4]
  assign regs_439_io_reset = reset; // @[RegFile.scala 78:19:@47879.4]
  assign regs_439_io_enable = 1'h1; // @[RegFile.scala 74:20:@47873.4]
  assign regs_440_clock = clock; // @[:@47882.4]
  assign regs_440_reset = io_reset; // @[:@47883.4 RegFile.scala 76:16:@47890.4]
  assign regs_440_io_in = 64'h0; // @[RegFile.scala 75:16:@47889.4]
  assign regs_440_io_reset = reset; // @[RegFile.scala 78:19:@47893.4]
  assign regs_440_io_enable = 1'h1; // @[RegFile.scala 74:20:@47887.4]
  assign regs_441_clock = clock; // @[:@47896.4]
  assign regs_441_reset = io_reset; // @[:@47897.4 RegFile.scala 76:16:@47904.4]
  assign regs_441_io_in = 64'h0; // @[RegFile.scala 75:16:@47903.4]
  assign regs_441_io_reset = reset; // @[RegFile.scala 78:19:@47907.4]
  assign regs_441_io_enable = 1'h1; // @[RegFile.scala 74:20:@47901.4]
  assign regs_442_clock = clock; // @[:@47910.4]
  assign regs_442_reset = io_reset; // @[:@47911.4 RegFile.scala 76:16:@47918.4]
  assign regs_442_io_in = 64'h0; // @[RegFile.scala 75:16:@47917.4]
  assign regs_442_io_reset = reset; // @[RegFile.scala 78:19:@47921.4]
  assign regs_442_io_enable = 1'h1; // @[RegFile.scala 74:20:@47915.4]
  assign regs_443_clock = clock; // @[:@47924.4]
  assign regs_443_reset = io_reset; // @[:@47925.4 RegFile.scala 76:16:@47932.4]
  assign regs_443_io_in = 64'h0; // @[RegFile.scala 75:16:@47931.4]
  assign regs_443_io_reset = reset; // @[RegFile.scala 78:19:@47935.4]
  assign regs_443_io_enable = 1'h1; // @[RegFile.scala 74:20:@47929.4]
  assign regs_444_clock = clock; // @[:@47938.4]
  assign regs_444_reset = io_reset; // @[:@47939.4 RegFile.scala 76:16:@47946.4]
  assign regs_444_io_in = 64'h0; // @[RegFile.scala 75:16:@47945.4]
  assign regs_444_io_reset = reset; // @[RegFile.scala 78:19:@47949.4]
  assign regs_444_io_enable = 1'h1; // @[RegFile.scala 74:20:@47943.4]
  assign regs_445_clock = clock; // @[:@47952.4]
  assign regs_445_reset = io_reset; // @[:@47953.4 RegFile.scala 76:16:@47960.4]
  assign regs_445_io_in = 64'h0; // @[RegFile.scala 75:16:@47959.4]
  assign regs_445_io_reset = reset; // @[RegFile.scala 78:19:@47963.4]
  assign regs_445_io_enable = 1'h1; // @[RegFile.scala 74:20:@47957.4]
  assign regs_446_clock = clock; // @[:@47966.4]
  assign regs_446_reset = io_reset; // @[:@47967.4 RegFile.scala 76:16:@47974.4]
  assign regs_446_io_in = 64'h0; // @[RegFile.scala 75:16:@47973.4]
  assign regs_446_io_reset = reset; // @[RegFile.scala 78:19:@47977.4]
  assign regs_446_io_enable = 1'h1; // @[RegFile.scala 74:20:@47971.4]
  assign regs_447_clock = clock; // @[:@47980.4]
  assign regs_447_reset = io_reset; // @[:@47981.4 RegFile.scala 76:16:@47988.4]
  assign regs_447_io_in = 64'h0; // @[RegFile.scala 75:16:@47987.4]
  assign regs_447_io_reset = reset; // @[RegFile.scala 78:19:@47991.4]
  assign regs_447_io_enable = 1'h1; // @[RegFile.scala 74:20:@47985.4]
  assign regs_448_clock = clock; // @[:@47994.4]
  assign regs_448_reset = io_reset; // @[:@47995.4 RegFile.scala 76:16:@48002.4]
  assign regs_448_io_in = 64'h0; // @[RegFile.scala 75:16:@48001.4]
  assign regs_448_io_reset = reset; // @[RegFile.scala 78:19:@48005.4]
  assign regs_448_io_enable = 1'h1; // @[RegFile.scala 74:20:@47999.4]
  assign regs_449_clock = clock; // @[:@48008.4]
  assign regs_449_reset = io_reset; // @[:@48009.4 RegFile.scala 76:16:@48016.4]
  assign regs_449_io_in = 64'h0; // @[RegFile.scala 75:16:@48015.4]
  assign regs_449_io_reset = reset; // @[RegFile.scala 78:19:@48019.4]
  assign regs_449_io_enable = 1'h1; // @[RegFile.scala 74:20:@48013.4]
  assign regs_450_clock = clock; // @[:@48022.4]
  assign regs_450_reset = io_reset; // @[:@48023.4 RegFile.scala 76:16:@48030.4]
  assign regs_450_io_in = 64'h0; // @[RegFile.scala 75:16:@48029.4]
  assign regs_450_io_reset = reset; // @[RegFile.scala 78:19:@48033.4]
  assign regs_450_io_enable = 1'h1; // @[RegFile.scala 74:20:@48027.4]
  assign regs_451_clock = clock; // @[:@48036.4]
  assign regs_451_reset = io_reset; // @[:@48037.4 RegFile.scala 76:16:@48044.4]
  assign regs_451_io_in = 64'h0; // @[RegFile.scala 75:16:@48043.4]
  assign regs_451_io_reset = reset; // @[RegFile.scala 78:19:@48047.4]
  assign regs_451_io_enable = 1'h1; // @[RegFile.scala 74:20:@48041.4]
  assign regs_452_clock = clock; // @[:@48050.4]
  assign regs_452_reset = io_reset; // @[:@48051.4 RegFile.scala 76:16:@48058.4]
  assign regs_452_io_in = 64'h0; // @[RegFile.scala 75:16:@48057.4]
  assign regs_452_io_reset = reset; // @[RegFile.scala 78:19:@48061.4]
  assign regs_452_io_enable = 1'h1; // @[RegFile.scala 74:20:@48055.4]
  assign regs_453_clock = clock; // @[:@48064.4]
  assign regs_453_reset = io_reset; // @[:@48065.4 RegFile.scala 76:16:@48072.4]
  assign regs_453_io_in = 64'h0; // @[RegFile.scala 75:16:@48071.4]
  assign regs_453_io_reset = reset; // @[RegFile.scala 78:19:@48075.4]
  assign regs_453_io_enable = 1'h1; // @[RegFile.scala 74:20:@48069.4]
  assign regs_454_clock = clock; // @[:@48078.4]
  assign regs_454_reset = io_reset; // @[:@48079.4 RegFile.scala 76:16:@48086.4]
  assign regs_454_io_in = 64'h0; // @[RegFile.scala 75:16:@48085.4]
  assign regs_454_io_reset = reset; // @[RegFile.scala 78:19:@48089.4]
  assign regs_454_io_enable = 1'h1; // @[RegFile.scala 74:20:@48083.4]
  assign regs_455_clock = clock; // @[:@48092.4]
  assign regs_455_reset = io_reset; // @[:@48093.4 RegFile.scala 76:16:@48100.4]
  assign regs_455_io_in = 64'h0; // @[RegFile.scala 75:16:@48099.4]
  assign regs_455_io_reset = reset; // @[RegFile.scala 78:19:@48103.4]
  assign regs_455_io_enable = 1'h1; // @[RegFile.scala 74:20:@48097.4]
  assign regs_456_clock = clock; // @[:@48106.4]
  assign regs_456_reset = io_reset; // @[:@48107.4 RegFile.scala 76:16:@48114.4]
  assign regs_456_io_in = 64'h0; // @[RegFile.scala 75:16:@48113.4]
  assign regs_456_io_reset = reset; // @[RegFile.scala 78:19:@48117.4]
  assign regs_456_io_enable = 1'h1; // @[RegFile.scala 74:20:@48111.4]
  assign regs_457_clock = clock; // @[:@48120.4]
  assign regs_457_reset = io_reset; // @[:@48121.4 RegFile.scala 76:16:@48128.4]
  assign regs_457_io_in = 64'h0; // @[RegFile.scala 75:16:@48127.4]
  assign regs_457_io_reset = reset; // @[RegFile.scala 78:19:@48131.4]
  assign regs_457_io_enable = 1'h1; // @[RegFile.scala 74:20:@48125.4]
  assign regs_458_clock = clock; // @[:@48134.4]
  assign regs_458_reset = io_reset; // @[:@48135.4 RegFile.scala 76:16:@48142.4]
  assign regs_458_io_in = 64'h0; // @[RegFile.scala 75:16:@48141.4]
  assign regs_458_io_reset = reset; // @[RegFile.scala 78:19:@48145.4]
  assign regs_458_io_enable = 1'h1; // @[RegFile.scala 74:20:@48139.4]
  assign regs_459_clock = clock; // @[:@48148.4]
  assign regs_459_reset = io_reset; // @[:@48149.4 RegFile.scala 76:16:@48156.4]
  assign regs_459_io_in = 64'h0; // @[RegFile.scala 75:16:@48155.4]
  assign regs_459_io_reset = reset; // @[RegFile.scala 78:19:@48159.4]
  assign regs_459_io_enable = 1'h1; // @[RegFile.scala 74:20:@48153.4]
  assign regs_460_clock = clock; // @[:@48162.4]
  assign regs_460_reset = io_reset; // @[:@48163.4 RegFile.scala 76:16:@48170.4]
  assign regs_460_io_in = 64'h0; // @[RegFile.scala 75:16:@48169.4]
  assign regs_460_io_reset = reset; // @[RegFile.scala 78:19:@48173.4]
  assign regs_460_io_enable = 1'h1; // @[RegFile.scala 74:20:@48167.4]
  assign regs_461_clock = clock; // @[:@48176.4]
  assign regs_461_reset = io_reset; // @[:@48177.4 RegFile.scala 76:16:@48184.4]
  assign regs_461_io_in = 64'h0; // @[RegFile.scala 75:16:@48183.4]
  assign regs_461_io_reset = reset; // @[RegFile.scala 78:19:@48187.4]
  assign regs_461_io_enable = 1'h1; // @[RegFile.scala 74:20:@48181.4]
  assign regs_462_clock = clock; // @[:@48190.4]
  assign regs_462_reset = io_reset; // @[:@48191.4 RegFile.scala 76:16:@48198.4]
  assign regs_462_io_in = 64'h0; // @[RegFile.scala 75:16:@48197.4]
  assign regs_462_io_reset = reset; // @[RegFile.scala 78:19:@48201.4]
  assign regs_462_io_enable = 1'h1; // @[RegFile.scala 74:20:@48195.4]
  assign regs_463_clock = clock; // @[:@48204.4]
  assign regs_463_reset = io_reset; // @[:@48205.4 RegFile.scala 76:16:@48212.4]
  assign regs_463_io_in = 64'h0; // @[RegFile.scala 75:16:@48211.4]
  assign regs_463_io_reset = reset; // @[RegFile.scala 78:19:@48215.4]
  assign regs_463_io_enable = 1'h1; // @[RegFile.scala 74:20:@48209.4]
  assign regs_464_clock = clock; // @[:@48218.4]
  assign regs_464_reset = io_reset; // @[:@48219.4 RegFile.scala 76:16:@48226.4]
  assign regs_464_io_in = 64'h0; // @[RegFile.scala 75:16:@48225.4]
  assign regs_464_io_reset = reset; // @[RegFile.scala 78:19:@48229.4]
  assign regs_464_io_enable = 1'h1; // @[RegFile.scala 74:20:@48223.4]
  assign regs_465_clock = clock; // @[:@48232.4]
  assign regs_465_reset = io_reset; // @[:@48233.4 RegFile.scala 76:16:@48240.4]
  assign regs_465_io_in = 64'h0; // @[RegFile.scala 75:16:@48239.4]
  assign regs_465_io_reset = reset; // @[RegFile.scala 78:19:@48243.4]
  assign regs_465_io_enable = 1'h1; // @[RegFile.scala 74:20:@48237.4]
  assign regs_466_clock = clock; // @[:@48246.4]
  assign regs_466_reset = io_reset; // @[:@48247.4 RegFile.scala 76:16:@48254.4]
  assign regs_466_io_in = 64'h0; // @[RegFile.scala 75:16:@48253.4]
  assign regs_466_io_reset = reset; // @[RegFile.scala 78:19:@48257.4]
  assign regs_466_io_enable = 1'h1; // @[RegFile.scala 74:20:@48251.4]
  assign regs_467_clock = clock; // @[:@48260.4]
  assign regs_467_reset = io_reset; // @[:@48261.4 RegFile.scala 76:16:@48268.4]
  assign regs_467_io_in = 64'h0; // @[RegFile.scala 75:16:@48267.4]
  assign regs_467_io_reset = reset; // @[RegFile.scala 78:19:@48271.4]
  assign regs_467_io_enable = 1'h1; // @[RegFile.scala 74:20:@48265.4]
  assign regs_468_clock = clock; // @[:@48274.4]
  assign regs_468_reset = io_reset; // @[:@48275.4 RegFile.scala 76:16:@48282.4]
  assign regs_468_io_in = 64'h0; // @[RegFile.scala 75:16:@48281.4]
  assign regs_468_io_reset = reset; // @[RegFile.scala 78:19:@48285.4]
  assign regs_468_io_enable = 1'h1; // @[RegFile.scala 74:20:@48279.4]
  assign regs_469_clock = clock; // @[:@48288.4]
  assign regs_469_reset = io_reset; // @[:@48289.4 RegFile.scala 76:16:@48296.4]
  assign regs_469_io_in = 64'h0; // @[RegFile.scala 75:16:@48295.4]
  assign regs_469_io_reset = reset; // @[RegFile.scala 78:19:@48299.4]
  assign regs_469_io_enable = 1'h1; // @[RegFile.scala 74:20:@48293.4]
  assign regs_470_clock = clock; // @[:@48302.4]
  assign regs_470_reset = io_reset; // @[:@48303.4 RegFile.scala 76:16:@48310.4]
  assign regs_470_io_in = 64'h0; // @[RegFile.scala 75:16:@48309.4]
  assign regs_470_io_reset = reset; // @[RegFile.scala 78:19:@48313.4]
  assign regs_470_io_enable = 1'h1; // @[RegFile.scala 74:20:@48307.4]
  assign regs_471_clock = clock; // @[:@48316.4]
  assign regs_471_reset = io_reset; // @[:@48317.4 RegFile.scala 76:16:@48324.4]
  assign regs_471_io_in = 64'h0; // @[RegFile.scala 75:16:@48323.4]
  assign regs_471_io_reset = reset; // @[RegFile.scala 78:19:@48327.4]
  assign regs_471_io_enable = 1'h1; // @[RegFile.scala 74:20:@48321.4]
  assign regs_472_clock = clock; // @[:@48330.4]
  assign regs_472_reset = io_reset; // @[:@48331.4 RegFile.scala 76:16:@48338.4]
  assign regs_472_io_in = 64'h0; // @[RegFile.scala 75:16:@48337.4]
  assign regs_472_io_reset = reset; // @[RegFile.scala 78:19:@48341.4]
  assign regs_472_io_enable = 1'h1; // @[RegFile.scala 74:20:@48335.4]
  assign regs_473_clock = clock; // @[:@48344.4]
  assign regs_473_reset = io_reset; // @[:@48345.4 RegFile.scala 76:16:@48352.4]
  assign regs_473_io_in = 64'h0; // @[RegFile.scala 75:16:@48351.4]
  assign regs_473_io_reset = reset; // @[RegFile.scala 78:19:@48355.4]
  assign regs_473_io_enable = 1'h1; // @[RegFile.scala 74:20:@48349.4]
  assign regs_474_clock = clock; // @[:@48358.4]
  assign regs_474_reset = io_reset; // @[:@48359.4 RegFile.scala 76:16:@48366.4]
  assign regs_474_io_in = 64'h0; // @[RegFile.scala 75:16:@48365.4]
  assign regs_474_io_reset = reset; // @[RegFile.scala 78:19:@48369.4]
  assign regs_474_io_enable = 1'h1; // @[RegFile.scala 74:20:@48363.4]
  assign regs_475_clock = clock; // @[:@48372.4]
  assign regs_475_reset = io_reset; // @[:@48373.4 RegFile.scala 76:16:@48380.4]
  assign regs_475_io_in = 64'h0; // @[RegFile.scala 75:16:@48379.4]
  assign regs_475_io_reset = reset; // @[RegFile.scala 78:19:@48383.4]
  assign regs_475_io_enable = 1'h1; // @[RegFile.scala 74:20:@48377.4]
  assign regs_476_clock = clock; // @[:@48386.4]
  assign regs_476_reset = io_reset; // @[:@48387.4 RegFile.scala 76:16:@48394.4]
  assign regs_476_io_in = 64'h0; // @[RegFile.scala 75:16:@48393.4]
  assign regs_476_io_reset = reset; // @[RegFile.scala 78:19:@48397.4]
  assign regs_476_io_enable = 1'h1; // @[RegFile.scala 74:20:@48391.4]
  assign regs_477_clock = clock; // @[:@48400.4]
  assign regs_477_reset = io_reset; // @[:@48401.4 RegFile.scala 76:16:@48408.4]
  assign regs_477_io_in = 64'h0; // @[RegFile.scala 75:16:@48407.4]
  assign regs_477_io_reset = reset; // @[RegFile.scala 78:19:@48411.4]
  assign regs_477_io_enable = 1'h1; // @[RegFile.scala 74:20:@48405.4]
  assign regs_478_clock = clock; // @[:@48414.4]
  assign regs_478_reset = io_reset; // @[:@48415.4 RegFile.scala 76:16:@48422.4]
  assign regs_478_io_in = 64'h0; // @[RegFile.scala 75:16:@48421.4]
  assign regs_478_io_reset = reset; // @[RegFile.scala 78:19:@48425.4]
  assign regs_478_io_enable = 1'h1; // @[RegFile.scala 74:20:@48419.4]
  assign regs_479_clock = clock; // @[:@48428.4]
  assign regs_479_reset = io_reset; // @[:@48429.4 RegFile.scala 76:16:@48436.4]
  assign regs_479_io_in = 64'h0; // @[RegFile.scala 75:16:@48435.4]
  assign regs_479_io_reset = reset; // @[RegFile.scala 78:19:@48439.4]
  assign regs_479_io_enable = 1'h1; // @[RegFile.scala 74:20:@48433.4]
  assign regs_480_clock = clock; // @[:@48442.4]
  assign regs_480_reset = io_reset; // @[:@48443.4 RegFile.scala 76:16:@48450.4]
  assign regs_480_io_in = 64'h0; // @[RegFile.scala 75:16:@48449.4]
  assign regs_480_io_reset = reset; // @[RegFile.scala 78:19:@48453.4]
  assign regs_480_io_enable = 1'h1; // @[RegFile.scala 74:20:@48447.4]
  assign regs_481_clock = clock; // @[:@48456.4]
  assign regs_481_reset = io_reset; // @[:@48457.4 RegFile.scala 76:16:@48464.4]
  assign regs_481_io_in = 64'h0; // @[RegFile.scala 75:16:@48463.4]
  assign regs_481_io_reset = reset; // @[RegFile.scala 78:19:@48467.4]
  assign regs_481_io_enable = 1'h1; // @[RegFile.scala 74:20:@48461.4]
  assign regs_482_clock = clock; // @[:@48470.4]
  assign regs_482_reset = io_reset; // @[:@48471.4 RegFile.scala 76:16:@48478.4]
  assign regs_482_io_in = 64'h0; // @[RegFile.scala 75:16:@48477.4]
  assign regs_482_io_reset = reset; // @[RegFile.scala 78:19:@48481.4]
  assign regs_482_io_enable = 1'h1; // @[RegFile.scala 74:20:@48475.4]
  assign regs_483_clock = clock; // @[:@48484.4]
  assign regs_483_reset = io_reset; // @[:@48485.4 RegFile.scala 76:16:@48492.4]
  assign regs_483_io_in = 64'h0; // @[RegFile.scala 75:16:@48491.4]
  assign regs_483_io_reset = reset; // @[RegFile.scala 78:19:@48495.4]
  assign regs_483_io_enable = 1'h1; // @[RegFile.scala 74:20:@48489.4]
  assign regs_484_clock = clock; // @[:@48498.4]
  assign regs_484_reset = io_reset; // @[:@48499.4 RegFile.scala 76:16:@48506.4]
  assign regs_484_io_in = 64'h0; // @[RegFile.scala 75:16:@48505.4]
  assign regs_484_io_reset = reset; // @[RegFile.scala 78:19:@48509.4]
  assign regs_484_io_enable = 1'h1; // @[RegFile.scala 74:20:@48503.4]
  assign regs_485_clock = clock; // @[:@48512.4]
  assign regs_485_reset = io_reset; // @[:@48513.4 RegFile.scala 76:16:@48520.4]
  assign regs_485_io_in = 64'h0; // @[RegFile.scala 75:16:@48519.4]
  assign regs_485_io_reset = reset; // @[RegFile.scala 78:19:@48523.4]
  assign regs_485_io_enable = 1'h1; // @[RegFile.scala 74:20:@48517.4]
  assign regs_486_clock = clock; // @[:@48526.4]
  assign regs_486_reset = io_reset; // @[:@48527.4 RegFile.scala 76:16:@48534.4]
  assign regs_486_io_in = 64'h0; // @[RegFile.scala 75:16:@48533.4]
  assign regs_486_io_reset = reset; // @[RegFile.scala 78:19:@48537.4]
  assign regs_486_io_enable = 1'h1; // @[RegFile.scala 74:20:@48531.4]
  assign regs_487_clock = clock; // @[:@48540.4]
  assign regs_487_reset = io_reset; // @[:@48541.4 RegFile.scala 76:16:@48548.4]
  assign regs_487_io_in = 64'h0; // @[RegFile.scala 75:16:@48547.4]
  assign regs_487_io_reset = reset; // @[RegFile.scala 78:19:@48551.4]
  assign regs_487_io_enable = 1'h1; // @[RegFile.scala 74:20:@48545.4]
  assign regs_488_clock = clock; // @[:@48554.4]
  assign regs_488_reset = io_reset; // @[:@48555.4 RegFile.scala 76:16:@48562.4]
  assign regs_488_io_in = 64'h0; // @[RegFile.scala 75:16:@48561.4]
  assign regs_488_io_reset = reset; // @[RegFile.scala 78:19:@48565.4]
  assign regs_488_io_enable = 1'h1; // @[RegFile.scala 74:20:@48559.4]
  assign regs_489_clock = clock; // @[:@48568.4]
  assign regs_489_reset = io_reset; // @[:@48569.4 RegFile.scala 76:16:@48576.4]
  assign regs_489_io_in = 64'h0; // @[RegFile.scala 75:16:@48575.4]
  assign regs_489_io_reset = reset; // @[RegFile.scala 78:19:@48579.4]
  assign regs_489_io_enable = 1'h1; // @[RegFile.scala 74:20:@48573.4]
  assign regs_490_clock = clock; // @[:@48582.4]
  assign regs_490_reset = io_reset; // @[:@48583.4 RegFile.scala 76:16:@48590.4]
  assign regs_490_io_in = 64'h0; // @[RegFile.scala 75:16:@48589.4]
  assign regs_490_io_reset = reset; // @[RegFile.scala 78:19:@48593.4]
  assign regs_490_io_enable = 1'h1; // @[RegFile.scala 74:20:@48587.4]
  assign regs_491_clock = clock; // @[:@48596.4]
  assign regs_491_reset = io_reset; // @[:@48597.4 RegFile.scala 76:16:@48604.4]
  assign regs_491_io_in = 64'h0; // @[RegFile.scala 75:16:@48603.4]
  assign regs_491_io_reset = reset; // @[RegFile.scala 78:19:@48607.4]
  assign regs_491_io_enable = 1'h1; // @[RegFile.scala 74:20:@48601.4]
  assign regs_492_clock = clock; // @[:@48610.4]
  assign regs_492_reset = io_reset; // @[:@48611.4 RegFile.scala 76:16:@48618.4]
  assign regs_492_io_in = 64'h0; // @[RegFile.scala 75:16:@48617.4]
  assign regs_492_io_reset = reset; // @[RegFile.scala 78:19:@48621.4]
  assign regs_492_io_enable = 1'h1; // @[RegFile.scala 74:20:@48615.4]
  assign regs_493_clock = clock; // @[:@48624.4]
  assign regs_493_reset = io_reset; // @[:@48625.4 RegFile.scala 76:16:@48632.4]
  assign regs_493_io_in = 64'h0; // @[RegFile.scala 75:16:@48631.4]
  assign regs_493_io_reset = reset; // @[RegFile.scala 78:19:@48635.4]
  assign regs_493_io_enable = 1'h1; // @[RegFile.scala 74:20:@48629.4]
  assign regs_494_clock = clock; // @[:@48638.4]
  assign regs_494_reset = io_reset; // @[:@48639.4 RegFile.scala 76:16:@48646.4]
  assign regs_494_io_in = 64'h0; // @[RegFile.scala 75:16:@48645.4]
  assign regs_494_io_reset = reset; // @[RegFile.scala 78:19:@48649.4]
  assign regs_494_io_enable = 1'h1; // @[RegFile.scala 74:20:@48643.4]
  assign regs_495_clock = clock; // @[:@48652.4]
  assign regs_495_reset = io_reset; // @[:@48653.4 RegFile.scala 76:16:@48660.4]
  assign regs_495_io_in = 64'h0; // @[RegFile.scala 75:16:@48659.4]
  assign regs_495_io_reset = reset; // @[RegFile.scala 78:19:@48663.4]
  assign regs_495_io_enable = 1'h1; // @[RegFile.scala 74:20:@48657.4]
  assign regs_496_clock = clock; // @[:@48666.4]
  assign regs_496_reset = io_reset; // @[:@48667.4 RegFile.scala 76:16:@48674.4]
  assign regs_496_io_in = 64'h0; // @[RegFile.scala 75:16:@48673.4]
  assign regs_496_io_reset = reset; // @[RegFile.scala 78:19:@48677.4]
  assign regs_496_io_enable = 1'h1; // @[RegFile.scala 74:20:@48671.4]
  assign regs_497_clock = clock; // @[:@48680.4]
  assign regs_497_reset = io_reset; // @[:@48681.4 RegFile.scala 76:16:@48688.4]
  assign regs_497_io_in = 64'h0; // @[RegFile.scala 75:16:@48687.4]
  assign regs_497_io_reset = reset; // @[RegFile.scala 78:19:@48691.4]
  assign regs_497_io_enable = 1'h1; // @[RegFile.scala 74:20:@48685.4]
  assign regs_498_clock = clock; // @[:@48694.4]
  assign regs_498_reset = io_reset; // @[:@48695.4 RegFile.scala 76:16:@48702.4]
  assign regs_498_io_in = 64'h0; // @[RegFile.scala 75:16:@48701.4]
  assign regs_498_io_reset = reset; // @[RegFile.scala 78:19:@48705.4]
  assign regs_498_io_enable = 1'h1; // @[RegFile.scala 74:20:@48699.4]
  assign regs_499_clock = clock; // @[:@48708.4]
  assign regs_499_reset = io_reset; // @[:@48709.4 RegFile.scala 76:16:@48716.4]
  assign regs_499_io_in = 64'h0; // @[RegFile.scala 75:16:@48715.4]
  assign regs_499_io_reset = reset; // @[RegFile.scala 78:19:@48719.4]
  assign regs_499_io_enable = 1'h1; // @[RegFile.scala 74:20:@48713.4]
  assign regs_500_clock = clock; // @[:@48722.4]
  assign regs_500_reset = io_reset; // @[:@48723.4 RegFile.scala 76:16:@48730.4]
  assign regs_500_io_in = 64'h0; // @[RegFile.scala 75:16:@48729.4]
  assign regs_500_io_reset = reset; // @[RegFile.scala 78:19:@48733.4]
  assign regs_500_io_enable = 1'h1; // @[RegFile.scala 74:20:@48727.4]
  assign regs_501_clock = clock; // @[:@48736.4]
  assign regs_501_reset = io_reset; // @[:@48737.4 RegFile.scala 76:16:@48744.4]
  assign regs_501_io_in = 64'h0; // @[RegFile.scala 75:16:@48743.4]
  assign regs_501_io_reset = reset; // @[RegFile.scala 78:19:@48747.4]
  assign regs_501_io_enable = 1'h1; // @[RegFile.scala 74:20:@48741.4]
  assign regs_502_clock = clock; // @[:@48750.4]
  assign regs_502_reset = io_reset; // @[:@48751.4 RegFile.scala 76:16:@48758.4]
  assign regs_502_io_in = 64'h0; // @[RegFile.scala 75:16:@48757.4]
  assign regs_502_io_reset = reset; // @[RegFile.scala 78:19:@48761.4]
  assign regs_502_io_enable = 1'h1; // @[RegFile.scala 74:20:@48755.4]
  assign regs_503_clock = clock; // @[:@48764.4]
  assign regs_503_reset = io_reset; // @[:@48765.4 RegFile.scala 76:16:@48772.4]
  assign regs_503_io_in = 64'h0; // @[RegFile.scala 75:16:@48771.4]
  assign regs_503_io_reset = reset; // @[RegFile.scala 78:19:@48775.4]
  assign regs_503_io_enable = 1'h1; // @[RegFile.scala 74:20:@48769.4]
  assign regs_504_clock = clock; // @[:@48778.4]
  assign regs_504_reset = io_reset; // @[:@48779.4 RegFile.scala 76:16:@48786.4]
  assign regs_504_io_in = 64'h0; // @[RegFile.scala 75:16:@48785.4]
  assign regs_504_io_reset = reset; // @[RegFile.scala 78:19:@48789.4]
  assign regs_504_io_enable = 1'h1; // @[RegFile.scala 74:20:@48783.4]
  assign regs_505_clock = clock; // @[:@48792.4]
  assign regs_505_reset = io_reset; // @[:@48793.4 RegFile.scala 76:16:@48800.4]
  assign regs_505_io_in = 64'h0; // @[RegFile.scala 75:16:@48799.4]
  assign regs_505_io_reset = reset; // @[RegFile.scala 78:19:@48803.4]
  assign regs_505_io_enable = 1'h1; // @[RegFile.scala 74:20:@48797.4]
  assign regs_506_clock = clock; // @[:@48806.4]
  assign regs_506_reset = io_reset; // @[:@48807.4 RegFile.scala 76:16:@48814.4]
  assign regs_506_io_in = 64'h0; // @[RegFile.scala 75:16:@48813.4]
  assign regs_506_io_reset = reset; // @[RegFile.scala 78:19:@48817.4]
  assign regs_506_io_enable = 1'h1; // @[RegFile.scala 74:20:@48811.4]
  assign regs_507_clock = clock; // @[:@48820.4]
  assign regs_507_reset = io_reset; // @[:@48821.4 RegFile.scala 76:16:@48828.4]
  assign regs_507_io_in = 64'h0; // @[RegFile.scala 75:16:@48827.4]
  assign regs_507_io_reset = reset; // @[RegFile.scala 78:19:@48831.4]
  assign regs_507_io_enable = 1'h1; // @[RegFile.scala 74:20:@48825.4]
  assign regs_508_clock = clock; // @[:@48834.4]
  assign regs_508_reset = io_reset; // @[:@48835.4 RegFile.scala 76:16:@48842.4]
  assign regs_508_io_in = 64'h0; // @[RegFile.scala 75:16:@48841.4]
  assign regs_508_io_reset = reset; // @[RegFile.scala 78:19:@48845.4]
  assign regs_508_io_enable = 1'h1; // @[RegFile.scala 74:20:@48839.4]
  assign regs_509_clock = clock; // @[:@48848.4]
  assign regs_509_reset = io_reset; // @[:@48849.4 RegFile.scala 76:16:@48856.4]
  assign regs_509_io_in = 64'h0; // @[RegFile.scala 75:16:@48855.4]
  assign regs_509_io_reset = reset; // @[RegFile.scala 78:19:@48859.4]
  assign regs_509_io_enable = 1'h1; // @[RegFile.scala 74:20:@48853.4]
  assign regs_510_clock = clock; // @[:@48862.4]
  assign regs_510_reset = io_reset; // @[:@48863.4 RegFile.scala 76:16:@48870.4]
  assign regs_510_io_in = 64'h0; // @[RegFile.scala 75:16:@48869.4]
  assign regs_510_io_reset = reset; // @[RegFile.scala 78:19:@48873.4]
  assign regs_510_io_enable = 1'h1; // @[RegFile.scala 74:20:@48867.4]
  assign regs_511_clock = clock; // @[:@48876.4]
  assign regs_511_reset = io_reset; // @[:@48877.4 RegFile.scala 76:16:@48884.4]
  assign regs_511_io_in = 64'h0; // @[RegFile.scala 75:16:@48883.4]
  assign regs_511_io_reset = reset; // @[RegFile.scala 78:19:@48887.4]
  assign regs_511_io_enable = 1'h1; // @[RegFile.scala 74:20:@48881.4]
  assign regs_512_clock = clock; // @[:@48890.4]
  assign regs_512_reset = io_reset; // @[:@48891.4 RegFile.scala 76:16:@48898.4]
  assign regs_512_io_in = 64'h0; // @[RegFile.scala 75:16:@48897.4]
  assign regs_512_io_reset = reset; // @[RegFile.scala 78:19:@48901.4]
  assign regs_512_io_enable = 1'h1; // @[RegFile.scala 74:20:@48895.4]
  assign regs_513_clock = clock; // @[:@48904.4]
  assign regs_513_reset = io_reset; // @[:@48905.4 RegFile.scala 76:16:@48912.4]
  assign regs_513_io_in = 64'h0; // @[RegFile.scala 75:16:@48911.4]
  assign regs_513_io_reset = reset; // @[RegFile.scala 78:19:@48915.4]
  assign regs_513_io_enable = 1'h1; // @[RegFile.scala 74:20:@48909.4]
  assign regs_514_clock = clock; // @[:@48918.4]
  assign regs_514_reset = io_reset; // @[:@48919.4 RegFile.scala 76:16:@48926.4]
  assign regs_514_io_in = 64'h0; // @[RegFile.scala 75:16:@48925.4]
  assign regs_514_io_reset = reset; // @[RegFile.scala 78:19:@48929.4]
  assign regs_514_io_enable = 1'h1; // @[RegFile.scala 74:20:@48923.4]
  assign regs_515_clock = clock; // @[:@48932.4]
  assign regs_515_reset = io_reset; // @[:@48933.4 RegFile.scala 76:16:@48940.4]
  assign regs_515_io_in = 64'h0; // @[RegFile.scala 75:16:@48939.4]
  assign regs_515_io_reset = reset; // @[RegFile.scala 78:19:@48943.4]
  assign regs_515_io_enable = 1'h1; // @[RegFile.scala 74:20:@48937.4]
  assign regs_516_clock = clock; // @[:@48946.4]
  assign regs_516_reset = io_reset; // @[:@48947.4 RegFile.scala 76:16:@48954.4]
  assign regs_516_io_in = 64'h0; // @[RegFile.scala 75:16:@48953.4]
  assign regs_516_io_reset = reset; // @[RegFile.scala 78:19:@48957.4]
  assign regs_516_io_enable = 1'h1; // @[RegFile.scala 74:20:@48951.4]
  assign regs_517_clock = clock; // @[:@48960.4]
  assign regs_517_reset = io_reset; // @[:@48961.4 RegFile.scala 76:16:@48968.4]
  assign regs_517_io_in = 64'h0; // @[RegFile.scala 75:16:@48967.4]
  assign regs_517_io_reset = reset; // @[RegFile.scala 78:19:@48971.4]
  assign regs_517_io_enable = 1'h1; // @[RegFile.scala 74:20:@48965.4]
  assign regs_518_clock = clock; // @[:@48974.4]
  assign regs_518_reset = io_reset; // @[:@48975.4 RegFile.scala 76:16:@48982.4]
  assign regs_518_io_in = 64'h0; // @[RegFile.scala 75:16:@48981.4]
  assign regs_518_io_reset = reset; // @[RegFile.scala 78:19:@48985.4]
  assign regs_518_io_enable = 1'h1; // @[RegFile.scala 74:20:@48979.4]
  assign regs_519_clock = clock; // @[:@48988.4]
  assign regs_519_reset = io_reset; // @[:@48989.4 RegFile.scala 76:16:@48996.4]
  assign regs_519_io_in = 64'h0; // @[RegFile.scala 75:16:@48995.4]
  assign regs_519_io_reset = reset; // @[RegFile.scala 78:19:@48999.4]
  assign regs_519_io_enable = 1'h1; // @[RegFile.scala 74:20:@48993.4]
  assign regs_520_clock = clock; // @[:@49002.4]
  assign regs_520_reset = io_reset; // @[:@49003.4 RegFile.scala 76:16:@49010.4]
  assign regs_520_io_in = 64'h0; // @[RegFile.scala 75:16:@49009.4]
  assign regs_520_io_reset = reset; // @[RegFile.scala 78:19:@49013.4]
  assign regs_520_io_enable = 1'h1; // @[RegFile.scala 74:20:@49007.4]
  assign regs_521_clock = clock; // @[:@49016.4]
  assign regs_521_reset = io_reset; // @[:@49017.4 RegFile.scala 76:16:@49024.4]
  assign regs_521_io_in = 64'h0; // @[RegFile.scala 75:16:@49023.4]
  assign regs_521_io_reset = reset; // @[RegFile.scala 78:19:@49027.4]
  assign regs_521_io_enable = 1'h1; // @[RegFile.scala 74:20:@49021.4]
  assign regs_522_clock = clock; // @[:@49030.4]
  assign regs_522_reset = io_reset; // @[:@49031.4 RegFile.scala 76:16:@49038.4]
  assign regs_522_io_in = 64'h0; // @[RegFile.scala 75:16:@49037.4]
  assign regs_522_io_reset = reset; // @[RegFile.scala 78:19:@49041.4]
  assign regs_522_io_enable = 1'h1; // @[RegFile.scala 74:20:@49035.4]
  assign regs_523_clock = clock; // @[:@49044.4]
  assign regs_523_reset = io_reset; // @[:@49045.4 RegFile.scala 76:16:@49052.4]
  assign regs_523_io_in = 64'h0; // @[RegFile.scala 75:16:@49051.4]
  assign regs_523_io_reset = reset; // @[RegFile.scala 78:19:@49055.4]
  assign regs_523_io_enable = 1'h1; // @[RegFile.scala 74:20:@49049.4]
  assign regs_524_clock = clock; // @[:@49058.4]
  assign regs_524_reset = io_reset; // @[:@49059.4 RegFile.scala 76:16:@49066.4]
  assign regs_524_io_in = 64'h0; // @[RegFile.scala 75:16:@49065.4]
  assign regs_524_io_reset = reset; // @[RegFile.scala 78:19:@49069.4]
  assign regs_524_io_enable = 1'h1; // @[RegFile.scala 74:20:@49063.4]
  assign regs_525_clock = clock; // @[:@49072.4]
  assign regs_525_reset = io_reset; // @[:@49073.4 RegFile.scala 76:16:@49080.4]
  assign regs_525_io_in = 64'h0; // @[RegFile.scala 75:16:@49079.4]
  assign regs_525_io_reset = reset; // @[RegFile.scala 78:19:@49083.4]
  assign regs_525_io_enable = 1'h1; // @[RegFile.scala 74:20:@49077.4]
  assign regs_526_clock = clock; // @[:@49086.4]
  assign regs_526_reset = io_reset; // @[:@49087.4 RegFile.scala 76:16:@49094.4]
  assign regs_526_io_in = 64'h0; // @[RegFile.scala 75:16:@49093.4]
  assign regs_526_io_reset = reset; // @[RegFile.scala 78:19:@49097.4]
  assign regs_526_io_enable = 1'h1; // @[RegFile.scala 74:20:@49091.4]
  assign regs_527_clock = clock; // @[:@49100.4]
  assign regs_527_reset = io_reset; // @[:@49101.4 RegFile.scala 76:16:@49108.4]
  assign regs_527_io_in = 64'h0; // @[RegFile.scala 75:16:@49107.4]
  assign regs_527_io_reset = reset; // @[RegFile.scala 78:19:@49111.4]
  assign regs_527_io_enable = 1'h1; // @[RegFile.scala 74:20:@49105.4]
  assign regs_528_clock = clock; // @[:@49114.4]
  assign regs_528_reset = io_reset; // @[:@49115.4 RegFile.scala 76:16:@49122.4]
  assign regs_528_io_in = 64'h0; // @[RegFile.scala 75:16:@49121.4]
  assign regs_528_io_reset = reset; // @[RegFile.scala 78:19:@49125.4]
  assign regs_528_io_enable = 1'h1; // @[RegFile.scala 74:20:@49119.4]
  assign regs_529_clock = clock; // @[:@49128.4]
  assign regs_529_reset = io_reset; // @[:@49129.4 RegFile.scala 76:16:@49136.4]
  assign regs_529_io_in = 64'h0; // @[RegFile.scala 75:16:@49135.4]
  assign regs_529_io_reset = reset; // @[RegFile.scala 78:19:@49139.4]
  assign regs_529_io_enable = 1'h1; // @[RegFile.scala 74:20:@49133.4]
  assign regs_530_clock = clock; // @[:@49142.4]
  assign regs_530_reset = io_reset; // @[:@49143.4 RegFile.scala 76:16:@49150.4]
  assign regs_530_io_in = 64'h0; // @[RegFile.scala 75:16:@49149.4]
  assign regs_530_io_reset = reset; // @[RegFile.scala 78:19:@49153.4]
  assign regs_530_io_enable = 1'h1; // @[RegFile.scala 74:20:@49147.4]
  assign regs_531_clock = clock; // @[:@49156.4]
  assign regs_531_reset = io_reset; // @[:@49157.4 RegFile.scala 76:16:@49164.4]
  assign regs_531_io_in = 64'h0; // @[RegFile.scala 75:16:@49163.4]
  assign regs_531_io_reset = reset; // @[RegFile.scala 78:19:@49167.4]
  assign regs_531_io_enable = 1'h1; // @[RegFile.scala 74:20:@49161.4]
  assign regs_532_clock = clock; // @[:@49170.4]
  assign regs_532_reset = io_reset; // @[:@49171.4 RegFile.scala 76:16:@49178.4]
  assign regs_532_io_in = 64'h0; // @[RegFile.scala 75:16:@49177.4]
  assign regs_532_io_reset = reset; // @[RegFile.scala 78:19:@49181.4]
  assign regs_532_io_enable = 1'h1; // @[RegFile.scala 74:20:@49175.4]
  assign regs_533_clock = clock; // @[:@49184.4]
  assign regs_533_reset = io_reset; // @[:@49185.4 RegFile.scala 76:16:@49192.4]
  assign regs_533_io_in = 64'h0; // @[RegFile.scala 75:16:@49191.4]
  assign regs_533_io_reset = reset; // @[RegFile.scala 78:19:@49195.4]
  assign regs_533_io_enable = 1'h1; // @[RegFile.scala 74:20:@49189.4]
  assign rport_io_ins_0 = regs_0_io_out; // @[RegFile.scala 97:16:@49735.4]
  assign rport_io_ins_1 = regs_1_io_out; // @[RegFile.scala 97:16:@49736.4]
  assign rport_io_ins_2 = regs_2_io_out; // @[RegFile.scala 97:16:@49737.4]
  assign rport_io_ins_3 = regs_3_io_out; // @[RegFile.scala 97:16:@49738.4]
  assign rport_io_ins_4 = regs_4_io_out; // @[RegFile.scala 97:16:@49739.4]
  assign rport_io_ins_5 = regs_5_io_out; // @[RegFile.scala 97:16:@49740.4]
  assign rport_io_ins_6 = regs_6_io_out; // @[RegFile.scala 97:16:@49741.4]
  assign rport_io_ins_7 = regs_7_io_out; // @[RegFile.scala 97:16:@49742.4]
  assign rport_io_ins_8 = regs_8_io_out; // @[RegFile.scala 97:16:@49743.4]
  assign rport_io_ins_9 = regs_9_io_out; // @[RegFile.scala 97:16:@49744.4]
  assign rport_io_ins_10 = regs_10_io_out; // @[RegFile.scala 97:16:@49745.4]
  assign rport_io_ins_11 = regs_11_io_out; // @[RegFile.scala 97:16:@49746.4]
  assign rport_io_ins_12 = regs_12_io_out; // @[RegFile.scala 97:16:@49747.4]
  assign rport_io_ins_13 = regs_13_io_out; // @[RegFile.scala 97:16:@49748.4]
  assign rport_io_ins_14 = regs_14_io_out; // @[RegFile.scala 97:16:@49749.4]
  assign rport_io_ins_15 = regs_15_io_out; // @[RegFile.scala 97:16:@49750.4]
  assign rport_io_ins_16 = regs_16_io_out; // @[RegFile.scala 97:16:@49751.4]
  assign rport_io_ins_17 = regs_17_io_out; // @[RegFile.scala 97:16:@49752.4]
  assign rport_io_ins_18 = regs_18_io_out; // @[RegFile.scala 97:16:@49753.4]
  assign rport_io_ins_19 = regs_19_io_out; // @[RegFile.scala 97:16:@49754.4]
  assign rport_io_ins_20 = regs_20_io_out; // @[RegFile.scala 97:16:@49755.4]
  assign rport_io_ins_21 = regs_21_io_out; // @[RegFile.scala 97:16:@49756.4]
  assign rport_io_ins_22 = regs_22_io_out; // @[RegFile.scala 97:16:@49757.4]
  assign rport_io_ins_23 = regs_23_io_out; // @[RegFile.scala 97:16:@49758.4]
  assign rport_io_ins_24 = regs_24_io_out; // @[RegFile.scala 97:16:@49759.4]
  assign rport_io_ins_25 = regs_25_io_out; // @[RegFile.scala 97:16:@49760.4]
  assign rport_io_ins_26 = regs_26_io_out; // @[RegFile.scala 97:16:@49761.4]
  assign rport_io_ins_27 = regs_27_io_out; // @[RegFile.scala 97:16:@49762.4]
  assign rport_io_ins_28 = regs_28_io_out; // @[RegFile.scala 97:16:@49763.4]
  assign rport_io_ins_29 = regs_29_io_out; // @[RegFile.scala 97:16:@49764.4]
  assign rport_io_ins_30 = regs_30_io_out; // @[RegFile.scala 97:16:@49765.4]
  assign rport_io_ins_31 = regs_31_io_out; // @[RegFile.scala 97:16:@49766.4]
  assign rport_io_ins_32 = regs_32_io_out; // @[RegFile.scala 97:16:@49767.4]
  assign rport_io_ins_33 = regs_33_io_out; // @[RegFile.scala 97:16:@49768.4]
  assign rport_io_ins_34 = regs_34_io_out; // @[RegFile.scala 97:16:@49769.4]
  assign rport_io_ins_35 = regs_35_io_out; // @[RegFile.scala 97:16:@49770.4]
  assign rport_io_ins_36 = regs_36_io_out; // @[RegFile.scala 97:16:@49771.4]
  assign rport_io_ins_37 = regs_37_io_out; // @[RegFile.scala 97:16:@49772.4]
  assign rport_io_ins_38 = regs_38_io_out; // @[RegFile.scala 97:16:@49773.4]
  assign rport_io_ins_39 = regs_39_io_out; // @[RegFile.scala 97:16:@49774.4]
  assign rport_io_ins_40 = regs_40_io_out; // @[RegFile.scala 97:16:@49775.4]
  assign rport_io_ins_41 = regs_41_io_out; // @[RegFile.scala 97:16:@49776.4]
  assign rport_io_ins_42 = regs_42_io_out; // @[RegFile.scala 97:16:@49777.4]
  assign rport_io_ins_43 = regs_43_io_out; // @[RegFile.scala 97:16:@49778.4]
  assign rport_io_ins_44 = regs_44_io_out; // @[RegFile.scala 97:16:@49779.4]
  assign rport_io_ins_45 = regs_45_io_out; // @[RegFile.scala 97:16:@49780.4]
  assign rport_io_ins_46 = regs_46_io_out; // @[RegFile.scala 97:16:@49781.4]
  assign rport_io_ins_47 = regs_47_io_out; // @[RegFile.scala 97:16:@49782.4]
  assign rport_io_ins_48 = regs_48_io_out; // @[RegFile.scala 97:16:@49783.4]
  assign rport_io_ins_49 = regs_49_io_out; // @[RegFile.scala 97:16:@49784.4]
  assign rport_io_ins_50 = regs_50_io_out; // @[RegFile.scala 97:16:@49785.4]
  assign rport_io_ins_51 = regs_51_io_out; // @[RegFile.scala 97:16:@49786.4]
  assign rport_io_ins_52 = regs_52_io_out; // @[RegFile.scala 97:16:@49787.4]
  assign rport_io_ins_53 = regs_53_io_out; // @[RegFile.scala 97:16:@49788.4]
  assign rport_io_ins_54 = regs_54_io_out; // @[RegFile.scala 97:16:@49789.4]
  assign rport_io_ins_55 = regs_55_io_out; // @[RegFile.scala 97:16:@49790.4]
  assign rport_io_ins_56 = regs_56_io_out; // @[RegFile.scala 97:16:@49791.4]
  assign rport_io_ins_57 = regs_57_io_out; // @[RegFile.scala 97:16:@49792.4]
  assign rport_io_ins_58 = regs_58_io_out; // @[RegFile.scala 97:16:@49793.4]
  assign rport_io_ins_59 = regs_59_io_out; // @[RegFile.scala 97:16:@49794.4]
  assign rport_io_ins_60 = regs_60_io_out; // @[RegFile.scala 97:16:@49795.4]
  assign rport_io_ins_61 = regs_61_io_out; // @[RegFile.scala 97:16:@49796.4]
  assign rport_io_ins_62 = regs_62_io_out; // @[RegFile.scala 97:16:@49797.4]
  assign rport_io_ins_63 = regs_63_io_out; // @[RegFile.scala 97:16:@49798.4]
  assign rport_io_ins_64 = regs_64_io_out; // @[RegFile.scala 97:16:@49799.4]
  assign rport_io_ins_65 = regs_65_io_out; // @[RegFile.scala 97:16:@49800.4]
  assign rport_io_ins_66 = regs_66_io_out; // @[RegFile.scala 97:16:@49801.4]
  assign rport_io_ins_67 = regs_67_io_out; // @[RegFile.scala 97:16:@49802.4]
  assign rport_io_ins_68 = regs_68_io_out; // @[RegFile.scala 97:16:@49803.4]
  assign rport_io_ins_69 = regs_69_io_out; // @[RegFile.scala 97:16:@49804.4]
  assign rport_io_ins_70 = regs_70_io_out; // @[RegFile.scala 97:16:@49805.4]
  assign rport_io_ins_71 = regs_71_io_out; // @[RegFile.scala 97:16:@49806.4]
  assign rport_io_ins_72 = regs_72_io_out; // @[RegFile.scala 97:16:@49807.4]
  assign rport_io_ins_73 = regs_73_io_out; // @[RegFile.scala 97:16:@49808.4]
  assign rport_io_ins_74 = regs_74_io_out; // @[RegFile.scala 97:16:@49809.4]
  assign rport_io_ins_75 = regs_75_io_out; // @[RegFile.scala 97:16:@49810.4]
  assign rport_io_ins_76 = regs_76_io_out; // @[RegFile.scala 97:16:@49811.4]
  assign rport_io_ins_77 = regs_77_io_out; // @[RegFile.scala 97:16:@49812.4]
  assign rport_io_ins_78 = regs_78_io_out; // @[RegFile.scala 97:16:@49813.4]
  assign rport_io_ins_79 = regs_79_io_out; // @[RegFile.scala 97:16:@49814.4]
  assign rport_io_ins_80 = regs_80_io_out; // @[RegFile.scala 97:16:@49815.4]
  assign rport_io_ins_81 = regs_81_io_out; // @[RegFile.scala 97:16:@49816.4]
  assign rport_io_ins_82 = regs_82_io_out; // @[RegFile.scala 97:16:@49817.4]
  assign rport_io_ins_83 = regs_83_io_out; // @[RegFile.scala 97:16:@49818.4]
  assign rport_io_ins_84 = regs_84_io_out; // @[RegFile.scala 97:16:@49819.4]
  assign rport_io_ins_85 = regs_85_io_out; // @[RegFile.scala 97:16:@49820.4]
  assign rport_io_ins_86 = regs_86_io_out; // @[RegFile.scala 97:16:@49821.4]
  assign rport_io_ins_87 = regs_87_io_out; // @[RegFile.scala 97:16:@49822.4]
  assign rport_io_ins_88 = regs_88_io_out; // @[RegFile.scala 97:16:@49823.4]
  assign rport_io_ins_89 = regs_89_io_out; // @[RegFile.scala 97:16:@49824.4]
  assign rport_io_ins_90 = regs_90_io_out; // @[RegFile.scala 97:16:@49825.4]
  assign rport_io_ins_91 = regs_91_io_out; // @[RegFile.scala 97:16:@49826.4]
  assign rport_io_ins_92 = regs_92_io_out; // @[RegFile.scala 97:16:@49827.4]
  assign rport_io_ins_93 = regs_93_io_out; // @[RegFile.scala 97:16:@49828.4]
  assign rport_io_ins_94 = regs_94_io_out; // @[RegFile.scala 97:16:@49829.4]
  assign rport_io_ins_95 = regs_95_io_out; // @[RegFile.scala 97:16:@49830.4]
  assign rport_io_ins_96 = regs_96_io_out; // @[RegFile.scala 97:16:@49831.4]
  assign rport_io_ins_97 = regs_97_io_out; // @[RegFile.scala 97:16:@49832.4]
  assign rport_io_ins_98 = regs_98_io_out; // @[RegFile.scala 97:16:@49833.4]
  assign rport_io_ins_99 = regs_99_io_out; // @[RegFile.scala 97:16:@49834.4]
  assign rport_io_ins_100 = regs_100_io_out; // @[RegFile.scala 97:16:@49835.4]
  assign rport_io_ins_101 = regs_101_io_out; // @[RegFile.scala 97:16:@49836.4]
  assign rport_io_ins_102 = regs_102_io_out; // @[RegFile.scala 97:16:@49837.4]
  assign rport_io_ins_103 = regs_103_io_out; // @[RegFile.scala 97:16:@49838.4]
  assign rport_io_ins_104 = regs_104_io_out; // @[RegFile.scala 97:16:@49839.4]
  assign rport_io_ins_105 = regs_105_io_out; // @[RegFile.scala 97:16:@49840.4]
  assign rport_io_ins_106 = regs_106_io_out; // @[RegFile.scala 97:16:@49841.4]
  assign rport_io_ins_107 = regs_107_io_out; // @[RegFile.scala 97:16:@49842.4]
  assign rport_io_ins_108 = regs_108_io_out; // @[RegFile.scala 97:16:@49843.4]
  assign rport_io_ins_109 = regs_109_io_out; // @[RegFile.scala 97:16:@49844.4]
  assign rport_io_ins_110 = regs_110_io_out; // @[RegFile.scala 97:16:@49845.4]
  assign rport_io_ins_111 = regs_111_io_out; // @[RegFile.scala 97:16:@49846.4]
  assign rport_io_ins_112 = regs_112_io_out; // @[RegFile.scala 97:16:@49847.4]
  assign rport_io_ins_113 = regs_113_io_out; // @[RegFile.scala 97:16:@49848.4]
  assign rport_io_ins_114 = regs_114_io_out; // @[RegFile.scala 97:16:@49849.4]
  assign rport_io_ins_115 = regs_115_io_out; // @[RegFile.scala 97:16:@49850.4]
  assign rport_io_ins_116 = regs_116_io_out; // @[RegFile.scala 97:16:@49851.4]
  assign rport_io_ins_117 = regs_117_io_out; // @[RegFile.scala 97:16:@49852.4]
  assign rport_io_ins_118 = regs_118_io_out; // @[RegFile.scala 97:16:@49853.4]
  assign rport_io_ins_119 = regs_119_io_out; // @[RegFile.scala 97:16:@49854.4]
  assign rport_io_ins_120 = regs_120_io_out; // @[RegFile.scala 97:16:@49855.4]
  assign rport_io_ins_121 = regs_121_io_out; // @[RegFile.scala 97:16:@49856.4]
  assign rport_io_ins_122 = regs_122_io_out; // @[RegFile.scala 97:16:@49857.4]
  assign rport_io_ins_123 = regs_123_io_out; // @[RegFile.scala 97:16:@49858.4]
  assign rport_io_ins_124 = regs_124_io_out; // @[RegFile.scala 97:16:@49859.4]
  assign rport_io_ins_125 = regs_125_io_out; // @[RegFile.scala 97:16:@49860.4]
  assign rport_io_ins_126 = regs_126_io_out; // @[RegFile.scala 97:16:@49861.4]
  assign rport_io_ins_127 = regs_127_io_out; // @[RegFile.scala 97:16:@49862.4]
  assign rport_io_ins_128 = regs_128_io_out; // @[RegFile.scala 97:16:@49863.4]
  assign rport_io_ins_129 = regs_129_io_out; // @[RegFile.scala 97:16:@49864.4]
  assign rport_io_ins_130 = regs_130_io_out; // @[RegFile.scala 97:16:@49865.4]
  assign rport_io_ins_131 = regs_131_io_out; // @[RegFile.scala 97:16:@49866.4]
  assign rport_io_ins_132 = regs_132_io_out; // @[RegFile.scala 97:16:@49867.4]
  assign rport_io_ins_133 = regs_133_io_out; // @[RegFile.scala 97:16:@49868.4]
  assign rport_io_ins_134 = regs_134_io_out; // @[RegFile.scala 97:16:@49869.4]
  assign rport_io_ins_135 = regs_135_io_out; // @[RegFile.scala 97:16:@49870.4]
  assign rport_io_ins_136 = regs_136_io_out; // @[RegFile.scala 97:16:@49871.4]
  assign rport_io_ins_137 = regs_137_io_out; // @[RegFile.scala 97:16:@49872.4]
  assign rport_io_ins_138 = regs_138_io_out; // @[RegFile.scala 97:16:@49873.4]
  assign rport_io_ins_139 = regs_139_io_out; // @[RegFile.scala 97:16:@49874.4]
  assign rport_io_ins_140 = regs_140_io_out; // @[RegFile.scala 97:16:@49875.4]
  assign rport_io_ins_141 = regs_141_io_out; // @[RegFile.scala 97:16:@49876.4]
  assign rport_io_ins_142 = regs_142_io_out; // @[RegFile.scala 97:16:@49877.4]
  assign rport_io_ins_143 = regs_143_io_out; // @[RegFile.scala 97:16:@49878.4]
  assign rport_io_ins_144 = regs_144_io_out; // @[RegFile.scala 97:16:@49879.4]
  assign rport_io_ins_145 = regs_145_io_out; // @[RegFile.scala 97:16:@49880.4]
  assign rport_io_ins_146 = regs_146_io_out; // @[RegFile.scala 97:16:@49881.4]
  assign rport_io_ins_147 = regs_147_io_out; // @[RegFile.scala 97:16:@49882.4]
  assign rport_io_ins_148 = regs_148_io_out; // @[RegFile.scala 97:16:@49883.4]
  assign rport_io_ins_149 = regs_149_io_out; // @[RegFile.scala 97:16:@49884.4]
  assign rport_io_ins_150 = regs_150_io_out; // @[RegFile.scala 97:16:@49885.4]
  assign rport_io_ins_151 = regs_151_io_out; // @[RegFile.scala 97:16:@49886.4]
  assign rport_io_ins_152 = regs_152_io_out; // @[RegFile.scala 97:16:@49887.4]
  assign rport_io_ins_153 = regs_153_io_out; // @[RegFile.scala 97:16:@49888.4]
  assign rport_io_ins_154 = regs_154_io_out; // @[RegFile.scala 97:16:@49889.4]
  assign rport_io_ins_155 = regs_155_io_out; // @[RegFile.scala 97:16:@49890.4]
  assign rport_io_ins_156 = regs_156_io_out; // @[RegFile.scala 97:16:@49891.4]
  assign rport_io_ins_157 = regs_157_io_out; // @[RegFile.scala 97:16:@49892.4]
  assign rport_io_ins_158 = regs_158_io_out; // @[RegFile.scala 97:16:@49893.4]
  assign rport_io_ins_159 = regs_159_io_out; // @[RegFile.scala 97:16:@49894.4]
  assign rport_io_ins_160 = regs_160_io_out; // @[RegFile.scala 97:16:@49895.4]
  assign rport_io_ins_161 = regs_161_io_out; // @[RegFile.scala 97:16:@49896.4]
  assign rport_io_ins_162 = regs_162_io_out; // @[RegFile.scala 97:16:@49897.4]
  assign rport_io_ins_163 = regs_163_io_out; // @[RegFile.scala 97:16:@49898.4]
  assign rport_io_ins_164 = regs_164_io_out; // @[RegFile.scala 97:16:@49899.4]
  assign rport_io_ins_165 = regs_165_io_out; // @[RegFile.scala 97:16:@49900.4]
  assign rport_io_ins_166 = regs_166_io_out; // @[RegFile.scala 97:16:@49901.4]
  assign rport_io_ins_167 = regs_167_io_out; // @[RegFile.scala 97:16:@49902.4]
  assign rport_io_ins_168 = regs_168_io_out; // @[RegFile.scala 97:16:@49903.4]
  assign rport_io_ins_169 = regs_169_io_out; // @[RegFile.scala 97:16:@49904.4]
  assign rport_io_ins_170 = regs_170_io_out; // @[RegFile.scala 97:16:@49905.4]
  assign rport_io_ins_171 = regs_171_io_out; // @[RegFile.scala 97:16:@49906.4]
  assign rport_io_ins_172 = regs_172_io_out; // @[RegFile.scala 97:16:@49907.4]
  assign rport_io_ins_173 = regs_173_io_out; // @[RegFile.scala 97:16:@49908.4]
  assign rport_io_ins_174 = regs_174_io_out; // @[RegFile.scala 97:16:@49909.4]
  assign rport_io_ins_175 = regs_175_io_out; // @[RegFile.scala 97:16:@49910.4]
  assign rport_io_ins_176 = regs_176_io_out; // @[RegFile.scala 97:16:@49911.4]
  assign rport_io_ins_177 = regs_177_io_out; // @[RegFile.scala 97:16:@49912.4]
  assign rport_io_ins_178 = regs_178_io_out; // @[RegFile.scala 97:16:@49913.4]
  assign rport_io_ins_179 = regs_179_io_out; // @[RegFile.scala 97:16:@49914.4]
  assign rport_io_ins_180 = regs_180_io_out; // @[RegFile.scala 97:16:@49915.4]
  assign rport_io_ins_181 = regs_181_io_out; // @[RegFile.scala 97:16:@49916.4]
  assign rport_io_ins_182 = regs_182_io_out; // @[RegFile.scala 97:16:@49917.4]
  assign rport_io_ins_183 = regs_183_io_out; // @[RegFile.scala 97:16:@49918.4]
  assign rport_io_ins_184 = regs_184_io_out; // @[RegFile.scala 97:16:@49919.4]
  assign rport_io_ins_185 = regs_185_io_out; // @[RegFile.scala 97:16:@49920.4]
  assign rport_io_ins_186 = regs_186_io_out; // @[RegFile.scala 97:16:@49921.4]
  assign rport_io_ins_187 = regs_187_io_out; // @[RegFile.scala 97:16:@49922.4]
  assign rport_io_ins_188 = regs_188_io_out; // @[RegFile.scala 97:16:@49923.4]
  assign rport_io_ins_189 = regs_189_io_out; // @[RegFile.scala 97:16:@49924.4]
  assign rport_io_ins_190 = regs_190_io_out; // @[RegFile.scala 97:16:@49925.4]
  assign rport_io_ins_191 = regs_191_io_out; // @[RegFile.scala 97:16:@49926.4]
  assign rport_io_ins_192 = regs_192_io_out; // @[RegFile.scala 97:16:@49927.4]
  assign rport_io_ins_193 = regs_193_io_out; // @[RegFile.scala 97:16:@49928.4]
  assign rport_io_ins_194 = regs_194_io_out; // @[RegFile.scala 97:16:@49929.4]
  assign rport_io_ins_195 = regs_195_io_out; // @[RegFile.scala 97:16:@49930.4]
  assign rport_io_ins_196 = regs_196_io_out; // @[RegFile.scala 97:16:@49931.4]
  assign rport_io_ins_197 = regs_197_io_out; // @[RegFile.scala 97:16:@49932.4]
  assign rport_io_ins_198 = regs_198_io_out; // @[RegFile.scala 97:16:@49933.4]
  assign rport_io_ins_199 = regs_199_io_out; // @[RegFile.scala 97:16:@49934.4]
  assign rport_io_ins_200 = regs_200_io_out; // @[RegFile.scala 97:16:@49935.4]
  assign rport_io_ins_201 = regs_201_io_out; // @[RegFile.scala 97:16:@49936.4]
  assign rport_io_ins_202 = regs_202_io_out; // @[RegFile.scala 97:16:@49937.4]
  assign rport_io_ins_203 = regs_203_io_out; // @[RegFile.scala 97:16:@49938.4]
  assign rport_io_ins_204 = regs_204_io_out; // @[RegFile.scala 97:16:@49939.4]
  assign rport_io_ins_205 = regs_205_io_out; // @[RegFile.scala 97:16:@49940.4]
  assign rport_io_ins_206 = regs_206_io_out; // @[RegFile.scala 97:16:@49941.4]
  assign rport_io_ins_207 = regs_207_io_out; // @[RegFile.scala 97:16:@49942.4]
  assign rport_io_ins_208 = regs_208_io_out; // @[RegFile.scala 97:16:@49943.4]
  assign rport_io_ins_209 = regs_209_io_out; // @[RegFile.scala 97:16:@49944.4]
  assign rport_io_ins_210 = regs_210_io_out; // @[RegFile.scala 97:16:@49945.4]
  assign rport_io_ins_211 = regs_211_io_out; // @[RegFile.scala 97:16:@49946.4]
  assign rport_io_ins_212 = regs_212_io_out; // @[RegFile.scala 97:16:@49947.4]
  assign rport_io_ins_213 = regs_213_io_out; // @[RegFile.scala 97:16:@49948.4]
  assign rport_io_ins_214 = regs_214_io_out; // @[RegFile.scala 97:16:@49949.4]
  assign rport_io_ins_215 = regs_215_io_out; // @[RegFile.scala 97:16:@49950.4]
  assign rport_io_ins_216 = regs_216_io_out; // @[RegFile.scala 97:16:@49951.4]
  assign rport_io_ins_217 = regs_217_io_out; // @[RegFile.scala 97:16:@49952.4]
  assign rport_io_ins_218 = regs_218_io_out; // @[RegFile.scala 97:16:@49953.4]
  assign rport_io_ins_219 = regs_219_io_out; // @[RegFile.scala 97:16:@49954.4]
  assign rport_io_ins_220 = regs_220_io_out; // @[RegFile.scala 97:16:@49955.4]
  assign rport_io_ins_221 = regs_221_io_out; // @[RegFile.scala 97:16:@49956.4]
  assign rport_io_ins_222 = regs_222_io_out; // @[RegFile.scala 97:16:@49957.4]
  assign rport_io_ins_223 = regs_223_io_out; // @[RegFile.scala 97:16:@49958.4]
  assign rport_io_ins_224 = regs_224_io_out; // @[RegFile.scala 97:16:@49959.4]
  assign rport_io_ins_225 = regs_225_io_out; // @[RegFile.scala 97:16:@49960.4]
  assign rport_io_ins_226 = regs_226_io_out; // @[RegFile.scala 97:16:@49961.4]
  assign rport_io_ins_227 = regs_227_io_out; // @[RegFile.scala 97:16:@49962.4]
  assign rport_io_ins_228 = regs_228_io_out; // @[RegFile.scala 97:16:@49963.4]
  assign rport_io_ins_229 = regs_229_io_out; // @[RegFile.scala 97:16:@49964.4]
  assign rport_io_ins_230 = regs_230_io_out; // @[RegFile.scala 97:16:@49965.4]
  assign rport_io_ins_231 = regs_231_io_out; // @[RegFile.scala 97:16:@49966.4]
  assign rport_io_ins_232 = regs_232_io_out; // @[RegFile.scala 97:16:@49967.4]
  assign rport_io_ins_233 = regs_233_io_out; // @[RegFile.scala 97:16:@49968.4]
  assign rport_io_ins_234 = regs_234_io_out; // @[RegFile.scala 97:16:@49969.4]
  assign rport_io_ins_235 = regs_235_io_out; // @[RegFile.scala 97:16:@49970.4]
  assign rport_io_ins_236 = regs_236_io_out; // @[RegFile.scala 97:16:@49971.4]
  assign rport_io_ins_237 = regs_237_io_out; // @[RegFile.scala 97:16:@49972.4]
  assign rport_io_ins_238 = regs_238_io_out; // @[RegFile.scala 97:16:@49973.4]
  assign rport_io_ins_239 = regs_239_io_out; // @[RegFile.scala 97:16:@49974.4]
  assign rport_io_ins_240 = regs_240_io_out; // @[RegFile.scala 97:16:@49975.4]
  assign rport_io_ins_241 = regs_241_io_out; // @[RegFile.scala 97:16:@49976.4]
  assign rport_io_ins_242 = regs_242_io_out; // @[RegFile.scala 97:16:@49977.4]
  assign rport_io_ins_243 = regs_243_io_out; // @[RegFile.scala 97:16:@49978.4]
  assign rport_io_ins_244 = regs_244_io_out; // @[RegFile.scala 97:16:@49979.4]
  assign rport_io_ins_245 = regs_245_io_out; // @[RegFile.scala 97:16:@49980.4]
  assign rport_io_ins_246 = regs_246_io_out; // @[RegFile.scala 97:16:@49981.4]
  assign rport_io_ins_247 = regs_247_io_out; // @[RegFile.scala 97:16:@49982.4]
  assign rport_io_ins_248 = regs_248_io_out; // @[RegFile.scala 97:16:@49983.4]
  assign rport_io_ins_249 = regs_249_io_out; // @[RegFile.scala 97:16:@49984.4]
  assign rport_io_ins_250 = regs_250_io_out; // @[RegFile.scala 97:16:@49985.4]
  assign rport_io_ins_251 = regs_251_io_out; // @[RegFile.scala 97:16:@49986.4]
  assign rport_io_ins_252 = regs_252_io_out; // @[RegFile.scala 97:16:@49987.4]
  assign rport_io_ins_253 = regs_253_io_out; // @[RegFile.scala 97:16:@49988.4]
  assign rport_io_ins_254 = regs_254_io_out; // @[RegFile.scala 97:16:@49989.4]
  assign rport_io_ins_255 = regs_255_io_out; // @[RegFile.scala 97:16:@49990.4]
  assign rport_io_ins_256 = regs_256_io_out; // @[RegFile.scala 97:16:@49991.4]
  assign rport_io_ins_257 = regs_257_io_out; // @[RegFile.scala 97:16:@49992.4]
  assign rport_io_ins_258 = regs_258_io_out; // @[RegFile.scala 97:16:@49993.4]
  assign rport_io_ins_259 = regs_259_io_out; // @[RegFile.scala 97:16:@49994.4]
  assign rport_io_ins_260 = regs_260_io_out; // @[RegFile.scala 97:16:@49995.4]
  assign rport_io_ins_261 = regs_261_io_out; // @[RegFile.scala 97:16:@49996.4]
  assign rport_io_ins_262 = regs_262_io_out; // @[RegFile.scala 97:16:@49997.4]
  assign rport_io_ins_263 = regs_263_io_out; // @[RegFile.scala 97:16:@49998.4]
  assign rport_io_ins_264 = regs_264_io_out; // @[RegFile.scala 97:16:@49999.4]
  assign rport_io_ins_265 = regs_265_io_out; // @[RegFile.scala 97:16:@50000.4]
  assign rport_io_ins_266 = regs_266_io_out; // @[RegFile.scala 97:16:@50001.4]
  assign rport_io_ins_267 = regs_267_io_out; // @[RegFile.scala 97:16:@50002.4]
  assign rport_io_ins_268 = regs_268_io_out; // @[RegFile.scala 97:16:@50003.4]
  assign rport_io_ins_269 = regs_269_io_out; // @[RegFile.scala 97:16:@50004.4]
  assign rport_io_ins_270 = regs_270_io_out; // @[RegFile.scala 97:16:@50005.4]
  assign rport_io_ins_271 = regs_271_io_out; // @[RegFile.scala 97:16:@50006.4]
  assign rport_io_ins_272 = regs_272_io_out; // @[RegFile.scala 97:16:@50007.4]
  assign rport_io_ins_273 = regs_273_io_out; // @[RegFile.scala 97:16:@50008.4]
  assign rport_io_ins_274 = regs_274_io_out; // @[RegFile.scala 97:16:@50009.4]
  assign rport_io_ins_275 = regs_275_io_out; // @[RegFile.scala 97:16:@50010.4]
  assign rport_io_ins_276 = regs_276_io_out; // @[RegFile.scala 97:16:@50011.4]
  assign rport_io_ins_277 = regs_277_io_out; // @[RegFile.scala 97:16:@50012.4]
  assign rport_io_ins_278 = regs_278_io_out; // @[RegFile.scala 97:16:@50013.4]
  assign rport_io_ins_279 = regs_279_io_out; // @[RegFile.scala 97:16:@50014.4]
  assign rport_io_ins_280 = regs_280_io_out; // @[RegFile.scala 97:16:@50015.4]
  assign rport_io_ins_281 = regs_281_io_out; // @[RegFile.scala 97:16:@50016.4]
  assign rport_io_ins_282 = regs_282_io_out; // @[RegFile.scala 97:16:@50017.4]
  assign rport_io_ins_283 = regs_283_io_out; // @[RegFile.scala 97:16:@50018.4]
  assign rport_io_ins_284 = regs_284_io_out; // @[RegFile.scala 97:16:@50019.4]
  assign rport_io_ins_285 = regs_285_io_out; // @[RegFile.scala 97:16:@50020.4]
  assign rport_io_ins_286 = regs_286_io_out; // @[RegFile.scala 97:16:@50021.4]
  assign rport_io_ins_287 = regs_287_io_out; // @[RegFile.scala 97:16:@50022.4]
  assign rport_io_ins_288 = regs_288_io_out; // @[RegFile.scala 97:16:@50023.4]
  assign rport_io_ins_289 = regs_289_io_out; // @[RegFile.scala 97:16:@50024.4]
  assign rport_io_ins_290 = regs_290_io_out; // @[RegFile.scala 97:16:@50025.4]
  assign rport_io_ins_291 = regs_291_io_out; // @[RegFile.scala 97:16:@50026.4]
  assign rport_io_ins_292 = regs_292_io_out; // @[RegFile.scala 97:16:@50027.4]
  assign rport_io_ins_293 = regs_293_io_out; // @[RegFile.scala 97:16:@50028.4]
  assign rport_io_ins_294 = regs_294_io_out; // @[RegFile.scala 97:16:@50029.4]
  assign rport_io_ins_295 = regs_295_io_out; // @[RegFile.scala 97:16:@50030.4]
  assign rport_io_ins_296 = regs_296_io_out; // @[RegFile.scala 97:16:@50031.4]
  assign rport_io_ins_297 = regs_297_io_out; // @[RegFile.scala 97:16:@50032.4]
  assign rport_io_ins_298 = regs_298_io_out; // @[RegFile.scala 97:16:@50033.4]
  assign rport_io_ins_299 = regs_299_io_out; // @[RegFile.scala 97:16:@50034.4]
  assign rport_io_ins_300 = regs_300_io_out; // @[RegFile.scala 97:16:@50035.4]
  assign rport_io_ins_301 = regs_301_io_out; // @[RegFile.scala 97:16:@50036.4]
  assign rport_io_ins_302 = regs_302_io_out; // @[RegFile.scala 97:16:@50037.4]
  assign rport_io_ins_303 = regs_303_io_out; // @[RegFile.scala 97:16:@50038.4]
  assign rport_io_ins_304 = regs_304_io_out; // @[RegFile.scala 97:16:@50039.4]
  assign rport_io_ins_305 = regs_305_io_out; // @[RegFile.scala 97:16:@50040.4]
  assign rport_io_ins_306 = regs_306_io_out; // @[RegFile.scala 97:16:@50041.4]
  assign rport_io_ins_307 = regs_307_io_out; // @[RegFile.scala 97:16:@50042.4]
  assign rport_io_ins_308 = regs_308_io_out; // @[RegFile.scala 97:16:@50043.4]
  assign rport_io_ins_309 = regs_309_io_out; // @[RegFile.scala 97:16:@50044.4]
  assign rport_io_ins_310 = regs_310_io_out; // @[RegFile.scala 97:16:@50045.4]
  assign rport_io_ins_311 = regs_311_io_out; // @[RegFile.scala 97:16:@50046.4]
  assign rport_io_ins_312 = regs_312_io_out; // @[RegFile.scala 97:16:@50047.4]
  assign rport_io_ins_313 = regs_313_io_out; // @[RegFile.scala 97:16:@50048.4]
  assign rport_io_ins_314 = regs_314_io_out; // @[RegFile.scala 97:16:@50049.4]
  assign rport_io_ins_315 = regs_315_io_out; // @[RegFile.scala 97:16:@50050.4]
  assign rport_io_ins_316 = regs_316_io_out; // @[RegFile.scala 97:16:@50051.4]
  assign rport_io_ins_317 = regs_317_io_out; // @[RegFile.scala 97:16:@50052.4]
  assign rport_io_ins_318 = regs_318_io_out; // @[RegFile.scala 97:16:@50053.4]
  assign rport_io_ins_319 = regs_319_io_out; // @[RegFile.scala 97:16:@50054.4]
  assign rport_io_ins_320 = regs_320_io_out; // @[RegFile.scala 97:16:@50055.4]
  assign rport_io_ins_321 = regs_321_io_out; // @[RegFile.scala 97:16:@50056.4]
  assign rport_io_ins_322 = regs_322_io_out; // @[RegFile.scala 97:16:@50057.4]
  assign rport_io_ins_323 = regs_323_io_out; // @[RegFile.scala 97:16:@50058.4]
  assign rport_io_ins_324 = regs_324_io_out; // @[RegFile.scala 97:16:@50059.4]
  assign rport_io_ins_325 = regs_325_io_out; // @[RegFile.scala 97:16:@50060.4]
  assign rport_io_ins_326 = regs_326_io_out; // @[RegFile.scala 97:16:@50061.4]
  assign rport_io_ins_327 = regs_327_io_out; // @[RegFile.scala 97:16:@50062.4]
  assign rport_io_ins_328 = regs_328_io_out; // @[RegFile.scala 97:16:@50063.4]
  assign rport_io_ins_329 = regs_329_io_out; // @[RegFile.scala 97:16:@50064.4]
  assign rport_io_ins_330 = regs_330_io_out; // @[RegFile.scala 97:16:@50065.4]
  assign rport_io_ins_331 = regs_331_io_out; // @[RegFile.scala 97:16:@50066.4]
  assign rport_io_ins_332 = regs_332_io_out; // @[RegFile.scala 97:16:@50067.4]
  assign rport_io_ins_333 = regs_333_io_out; // @[RegFile.scala 97:16:@50068.4]
  assign rport_io_ins_334 = regs_334_io_out; // @[RegFile.scala 97:16:@50069.4]
  assign rport_io_ins_335 = regs_335_io_out; // @[RegFile.scala 97:16:@50070.4]
  assign rport_io_ins_336 = regs_336_io_out; // @[RegFile.scala 97:16:@50071.4]
  assign rport_io_ins_337 = regs_337_io_out; // @[RegFile.scala 97:16:@50072.4]
  assign rport_io_ins_338 = regs_338_io_out; // @[RegFile.scala 97:16:@50073.4]
  assign rport_io_ins_339 = regs_339_io_out; // @[RegFile.scala 97:16:@50074.4]
  assign rport_io_ins_340 = regs_340_io_out; // @[RegFile.scala 97:16:@50075.4]
  assign rport_io_ins_341 = regs_341_io_out; // @[RegFile.scala 97:16:@50076.4]
  assign rport_io_ins_342 = regs_342_io_out; // @[RegFile.scala 97:16:@50077.4]
  assign rport_io_ins_343 = regs_343_io_out; // @[RegFile.scala 97:16:@50078.4]
  assign rport_io_ins_344 = regs_344_io_out; // @[RegFile.scala 97:16:@50079.4]
  assign rport_io_ins_345 = regs_345_io_out; // @[RegFile.scala 97:16:@50080.4]
  assign rport_io_ins_346 = regs_346_io_out; // @[RegFile.scala 97:16:@50081.4]
  assign rport_io_ins_347 = regs_347_io_out; // @[RegFile.scala 97:16:@50082.4]
  assign rport_io_ins_348 = regs_348_io_out; // @[RegFile.scala 97:16:@50083.4]
  assign rport_io_ins_349 = regs_349_io_out; // @[RegFile.scala 97:16:@50084.4]
  assign rport_io_ins_350 = regs_350_io_out; // @[RegFile.scala 97:16:@50085.4]
  assign rport_io_ins_351 = regs_351_io_out; // @[RegFile.scala 97:16:@50086.4]
  assign rport_io_ins_352 = regs_352_io_out; // @[RegFile.scala 97:16:@50087.4]
  assign rport_io_ins_353 = regs_353_io_out; // @[RegFile.scala 97:16:@50088.4]
  assign rport_io_ins_354 = regs_354_io_out; // @[RegFile.scala 97:16:@50089.4]
  assign rport_io_ins_355 = regs_355_io_out; // @[RegFile.scala 97:16:@50090.4]
  assign rport_io_ins_356 = regs_356_io_out; // @[RegFile.scala 97:16:@50091.4]
  assign rport_io_ins_357 = regs_357_io_out; // @[RegFile.scala 97:16:@50092.4]
  assign rport_io_ins_358 = regs_358_io_out; // @[RegFile.scala 97:16:@50093.4]
  assign rport_io_ins_359 = regs_359_io_out; // @[RegFile.scala 97:16:@50094.4]
  assign rport_io_ins_360 = regs_360_io_out; // @[RegFile.scala 97:16:@50095.4]
  assign rport_io_ins_361 = regs_361_io_out; // @[RegFile.scala 97:16:@50096.4]
  assign rport_io_ins_362 = regs_362_io_out; // @[RegFile.scala 97:16:@50097.4]
  assign rport_io_ins_363 = regs_363_io_out; // @[RegFile.scala 97:16:@50098.4]
  assign rport_io_ins_364 = regs_364_io_out; // @[RegFile.scala 97:16:@50099.4]
  assign rport_io_ins_365 = regs_365_io_out; // @[RegFile.scala 97:16:@50100.4]
  assign rport_io_ins_366 = regs_366_io_out; // @[RegFile.scala 97:16:@50101.4]
  assign rport_io_ins_367 = regs_367_io_out; // @[RegFile.scala 97:16:@50102.4]
  assign rport_io_ins_368 = regs_368_io_out; // @[RegFile.scala 97:16:@50103.4]
  assign rport_io_ins_369 = regs_369_io_out; // @[RegFile.scala 97:16:@50104.4]
  assign rport_io_ins_370 = regs_370_io_out; // @[RegFile.scala 97:16:@50105.4]
  assign rport_io_ins_371 = regs_371_io_out; // @[RegFile.scala 97:16:@50106.4]
  assign rport_io_ins_372 = regs_372_io_out; // @[RegFile.scala 97:16:@50107.4]
  assign rport_io_ins_373 = regs_373_io_out; // @[RegFile.scala 97:16:@50108.4]
  assign rport_io_ins_374 = regs_374_io_out; // @[RegFile.scala 97:16:@50109.4]
  assign rport_io_ins_375 = regs_375_io_out; // @[RegFile.scala 97:16:@50110.4]
  assign rport_io_ins_376 = regs_376_io_out; // @[RegFile.scala 97:16:@50111.4]
  assign rport_io_ins_377 = regs_377_io_out; // @[RegFile.scala 97:16:@50112.4]
  assign rport_io_ins_378 = regs_378_io_out; // @[RegFile.scala 97:16:@50113.4]
  assign rport_io_ins_379 = regs_379_io_out; // @[RegFile.scala 97:16:@50114.4]
  assign rport_io_ins_380 = regs_380_io_out; // @[RegFile.scala 97:16:@50115.4]
  assign rport_io_ins_381 = regs_381_io_out; // @[RegFile.scala 97:16:@50116.4]
  assign rport_io_ins_382 = regs_382_io_out; // @[RegFile.scala 97:16:@50117.4]
  assign rport_io_ins_383 = regs_383_io_out; // @[RegFile.scala 97:16:@50118.4]
  assign rport_io_ins_384 = regs_384_io_out; // @[RegFile.scala 97:16:@50119.4]
  assign rport_io_ins_385 = regs_385_io_out; // @[RegFile.scala 97:16:@50120.4]
  assign rport_io_ins_386 = regs_386_io_out; // @[RegFile.scala 97:16:@50121.4]
  assign rport_io_ins_387 = regs_387_io_out; // @[RegFile.scala 97:16:@50122.4]
  assign rport_io_ins_388 = regs_388_io_out; // @[RegFile.scala 97:16:@50123.4]
  assign rport_io_ins_389 = regs_389_io_out; // @[RegFile.scala 97:16:@50124.4]
  assign rport_io_ins_390 = regs_390_io_out; // @[RegFile.scala 97:16:@50125.4]
  assign rport_io_ins_391 = regs_391_io_out; // @[RegFile.scala 97:16:@50126.4]
  assign rport_io_ins_392 = regs_392_io_out; // @[RegFile.scala 97:16:@50127.4]
  assign rport_io_ins_393 = regs_393_io_out; // @[RegFile.scala 97:16:@50128.4]
  assign rport_io_ins_394 = regs_394_io_out; // @[RegFile.scala 97:16:@50129.4]
  assign rport_io_ins_395 = regs_395_io_out; // @[RegFile.scala 97:16:@50130.4]
  assign rport_io_ins_396 = regs_396_io_out; // @[RegFile.scala 97:16:@50131.4]
  assign rport_io_ins_397 = regs_397_io_out; // @[RegFile.scala 97:16:@50132.4]
  assign rport_io_ins_398 = regs_398_io_out; // @[RegFile.scala 97:16:@50133.4]
  assign rport_io_ins_399 = regs_399_io_out; // @[RegFile.scala 97:16:@50134.4]
  assign rport_io_ins_400 = regs_400_io_out; // @[RegFile.scala 97:16:@50135.4]
  assign rport_io_ins_401 = regs_401_io_out; // @[RegFile.scala 97:16:@50136.4]
  assign rport_io_ins_402 = regs_402_io_out; // @[RegFile.scala 97:16:@50137.4]
  assign rport_io_ins_403 = regs_403_io_out; // @[RegFile.scala 97:16:@50138.4]
  assign rport_io_ins_404 = regs_404_io_out; // @[RegFile.scala 97:16:@50139.4]
  assign rport_io_ins_405 = regs_405_io_out; // @[RegFile.scala 97:16:@50140.4]
  assign rport_io_ins_406 = regs_406_io_out; // @[RegFile.scala 97:16:@50141.4]
  assign rport_io_ins_407 = regs_407_io_out; // @[RegFile.scala 97:16:@50142.4]
  assign rport_io_ins_408 = regs_408_io_out; // @[RegFile.scala 97:16:@50143.4]
  assign rport_io_ins_409 = regs_409_io_out; // @[RegFile.scala 97:16:@50144.4]
  assign rport_io_ins_410 = regs_410_io_out; // @[RegFile.scala 97:16:@50145.4]
  assign rport_io_ins_411 = regs_411_io_out; // @[RegFile.scala 97:16:@50146.4]
  assign rport_io_ins_412 = regs_412_io_out; // @[RegFile.scala 97:16:@50147.4]
  assign rport_io_ins_413 = regs_413_io_out; // @[RegFile.scala 97:16:@50148.4]
  assign rport_io_ins_414 = regs_414_io_out; // @[RegFile.scala 97:16:@50149.4]
  assign rport_io_ins_415 = regs_415_io_out; // @[RegFile.scala 97:16:@50150.4]
  assign rport_io_ins_416 = regs_416_io_out; // @[RegFile.scala 97:16:@50151.4]
  assign rport_io_ins_417 = regs_417_io_out; // @[RegFile.scala 97:16:@50152.4]
  assign rport_io_ins_418 = regs_418_io_out; // @[RegFile.scala 97:16:@50153.4]
  assign rport_io_ins_419 = regs_419_io_out; // @[RegFile.scala 97:16:@50154.4]
  assign rport_io_ins_420 = regs_420_io_out; // @[RegFile.scala 97:16:@50155.4]
  assign rport_io_ins_421 = regs_421_io_out; // @[RegFile.scala 97:16:@50156.4]
  assign rport_io_ins_422 = regs_422_io_out; // @[RegFile.scala 97:16:@50157.4]
  assign rport_io_ins_423 = regs_423_io_out; // @[RegFile.scala 97:16:@50158.4]
  assign rport_io_ins_424 = regs_424_io_out; // @[RegFile.scala 97:16:@50159.4]
  assign rport_io_ins_425 = regs_425_io_out; // @[RegFile.scala 97:16:@50160.4]
  assign rport_io_ins_426 = regs_426_io_out; // @[RegFile.scala 97:16:@50161.4]
  assign rport_io_ins_427 = regs_427_io_out; // @[RegFile.scala 97:16:@50162.4]
  assign rport_io_ins_428 = regs_428_io_out; // @[RegFile.scala 97:16:@50163.4]
  assign rport_io_ins_429 = regs_429_io_out; // @[RegFile.scala 97:16:@50164.4]
  assign rport_io_ins_430 = regs_430_io_out; // @[RegFile.scala 97:16:@50165.4]
  assign rport_io_ins_431 = regs_431_io_out; // @[RegFile.scala 97:16:@50166.4]
  assign rport_io_ins_432 = regs_432_io_out; // @[RegFile.scala 97:16:@50167.4]
  assign rport_io_ins_433 = regs_433_io_out; // @[RegFile.scala 97:16:@50168.4]
  assign rport_io_ins_434 = regs_434_io_out; // @[RegFile.scala 97:16:@50169.4]
  assign rport_io_ins_435 = regs_435_io_out; // @[RegFile.scala 97:16:@50170.4]
  assign rport_io_ins_436 = regs_436_io_out; // @[RegFile.scala 97:16:@50171.4]
  assign rport_io_ins_437 = regs_437_io_out; // @[RegFile.scala 97:16:@50172.4]
  assign rport_io_ins_438 = regs_438_io_out; // @[RegFile.scala 97:16:@50173.4]
  assign rport_io_ins_439 = regs_439_io_out; // @[RegFile.scala 97:16:@50174.4]
  assign rport_io_ins_440 = regs_440_io_out; // @[RegFile.scala 97:16:@50175.4]
  assign rport_io_ins_441 = regs_441_io_out; // @[RegFile.scala 97:16:@50176.4]
  assign rport_io_ins_442 = regs_442_io_out; // @[RegFile.scala 97:16:@50177.4]
  assign rport_io_ins_443 = regs_443_io_out; // @[RegFile.scala 97:16:@50178.4]
  assign rport_io_ins_444 = regs_444_io_out; // @[RegFile.scala 97:16:@50179.4]
  assign rport_io_ins_445 = regs_445_io_out; // @[RegFile.scala 97:16:@50180.4]
  assign rport_io_ins_446 = regs_446_io_out; // @[RegFile.scala 97:16:@50181.4]
  assign rport_io_ins_447 = regs_447_io_out; // @[RegFile.scala 97:16:@50182.4]
  assign rport_io_ins_448 = regs_448_io_out; // @[RegFile.scala 97:16:@50183.4]
  assign rport_io_ins_449 = regs_449_io_out; // @[RegFile.scala 97:16:@50184.4]
  assign rport_io_ins_450 = regs_450_io_out; // @[RegFile.scala 97:16:@50185.4]
  assign rport_io_ins_451 = regs_451_io_out; // @[RegFile.scala 97:16:@50186.4]
  assign rport_io_ins_452 = regs_452_io_out; // @[RegFile.scala 97:16:@50187.4]
  assign rport_io_ins_453 = regs_453_io_out; // @[RegFile.scala 97:16:@50188.4]
  assign rport_io_ins_454 = regs_454_io_out; // @[RegFile.scala 97:16:@50189.4]
  assign rport_io_ins_455 = regs_455_io_out; // @[RegFile.scala 97:16:@50190.4]
  assign rport_io_ins_456 = regs_456_io_out; // @[RegFile.scala 97:16:@50191.4]
  assign rport_io_ins_457 = regs_457_io_out; // @[RegFile.scala 97:16:@50192.4]
  assign rport_io_ins_458 = regs_458_io_out; // @[RegFile.scala 97:16:@50193.4]
  assign rport_io_ins_459 = regs_459_io_out; // @[RegFile.scala 97:16:@50194.4]
  assign rport_io_ins_460 = regs_460_io_out; // @[RegFile.scala 97:16:@50195.4]
  assign rport_io_ins_461 = regs_461_io_out; // @[RegFile.scala 97:16:@50196.4]
  assign rport_io_ins_462 = regs_462_io_out; // @[RegFile.scala 97:16:@50197.4]
  assign rport_io_ins_463 = regs_463_io_out; // @[RegFile.scala 97:16:@50198.4]
  assign rport_io_ins_464 = regs_464_io_out; // @[RegFile.scala 97:16:@50199.4]
  assign rport_io_ins_465 = regs_465_io_out; // @[RegFile.scala 97:16:@50200.4]
  assign rport_io_ins_466 = regs_466_io_out; // @[RegFile.scala 97:16:@50201.4]
  assign rport_io_ins_467 = regs_467_io_out; // @[RegFile.scala 97:16:@50202.4]
  assign rport_io_ins_468 = regs_468_io_out; // @[RegFile.scala 97:16:@50203.4]
  assign rport_io_ins_469 = regs_469_io_out; // @[RegFile.scala 97:16:@50204.4]
  assign rport_io_ins_470 = regs_470_io_out; // @[RegFile.scala 97:16:@50205.4]
  assign rport_io_ins_471 = regs_471_io_out; // @[RegFile.scala 97:16:@50206.4]
  assign rport_io_ins_472 = regs_472_io_out; // @[RegFile.scala 97:16:@50207.4]
  assign rport_io_ins_473 = regs_473_io_out; // @[RegFile.scala 97:16:@50208.4]
  assign rport_io_ins_474 = regs_474_io_out; // @[RegFile.scala 97:16:@50209.4]
  assign rport_io_ins_475 = regs_475_io_out; // @[RegFile.scala 97:16:@50210.4]
  assign rport_io_ins_476 = regs_476_io_out; // @[RegFile.scala 97:16:@50211.4]
  assign rport_io_ins_477 = regs_477_io_out; // @[RegFile.scala 97:16:@50212.4]
  assign rport_io_ins_478 = regs_478_io_out; // @[RegFile.scala 97:16:@50213.4]
  assign rport_io_ins_479 = regs_479_io_out; // @[RegFile.scala 97:16:@50214.4]
  assign rport_io_ins_480 = regs_480_io_out; // @[RegFile.scala 97:16:@50215.4]
  assign rport_io_ins_481 = regs_481_io_out; // @[RegFile.scala 97:16:@50216.4]
  assign rport_io_ins_482 = regs_482_io_out; // @[RegFile.scala 97:16:@50217.4]
  assign rport_io_ins_483 = regs_483_io_out; // @[RegFile.scala 97:16:@50218.4]
  assign rport_io_ins_484 = regs_484_io_out; // @[RegFile.scala 97:16:@50219.4]
  assign rport_io_ins_485 = regs_485_io_out; // @[RegFile.scala 97:16:@50220.4]
  assign rport_io_ins_486 = regs_486_io_out; // @[RegFile.scala 97:16:@50221.4]
  assign rport_io_ins_487 = regs_487_io_out; // @[RegFile.scala 97:16:@50222.4]
  assign rport_io_ins_488 = regs_488_io_out; // @[RegFile.scala 97:16:@50223.4]
  assign rport_io_ins_489 = regs_489_io_out; // @[RegFile.scala 97:16:@50224.4]
  assign rport_io_ins_490 = regs_490_io_out; // @[RegFile.scala 97:16:@50225.4]
  assign rport_io_ins_491 = regs_491_io_out; // @[RegFile.scala 97:16:@50226.4]
  assign rport_io_ins_492 = regs_492_io_out; // @[RegFile.scala 97:16:@50227.4]
  assign rport_io_ins_493 = regs_493_io_out; // @[RegFile.scala 97:16:@50228.4]
  assign rport_io_ins_494 = regs_494_io_out; // @[RegFile.scala 97:16:@50229.4]
  assign rport_io_ins_495 = regs_495_io_out; // @[RegFile.scala 97:16:@50230.4]
  assign rport_io_ins_496 = regs_496_io_out; // @[RegFile.scala 97:16:@50231.4]
  assign rport_io_ins_497 = regs_497_io_out; // @[RegFile.scala 97:16:@50232.4]
  assign rport_io_ins_498 = regs_498_io_out; // @[RegFile.scala 97:16:@50233.4]
  assign rport_io_ins_499 = regs_499_io_out; // @[RegFile.scala 97:16:@50234.4]
  assign rport_io_ins_500 = regs_500_io_out; // @[RegFile.scala 97:16:@50235.4]
  assign rport_io_ins_501 = regs_501_io_out; // @[RegFile.scala 97:16:@50236.4]
  assign rport_io_ins_502 = regs_502_io_out; // @[RegFile.scala 97:16:@50237.4]
  assign rport_io_ins_503 = regs_503_io_out; // @[RegFile.scala 97:16:@50238.4]
  assign rport_io_ins_504 = regs_504_io_out; // @[RegFile.scala 97:16:@50239.4]
  assign rport_io_ins_505 = regs_505_io_out; // @[RegFile.scala 97:16:@50240.4]
  assign rport_io_ins_506 = regs_506_io_out; // @[RegFile.scala 97:16:@50241.4]
  assign rport_io_ins_507 = regs_507_io_out; // @[RegFile.scala 97:16:@50242.4]
  assign rport_io_ins_508 = regs_508_io_out; // @[RegFile.scala 97:16:@50243.4]
  assign rport_io_ins_509 = regs_509_io_out; // @[RegFile.scala 97:16:@50244.4]
  assign rport_io_ins_510 = regs_510_io_out; // @[RegFile.scala 97:16:@50245.4]
  assign rport_io_ins_511 = regs_511_io_out; // @[RegFile.scala 97:16:@50246.4]
  assign rport_io_ins_512 = regs_512_io_out; // @[RegFile.scala 97:16:@50247.4]
  assign rport_io_ins_513 = regs_513_io_out; // @[RegFile.scala 97:16:@50248.4]
  assign rport_io_ins_514 = regs_514_io_out; // @[RegFile.scala 97:16:@50249.4]
  assign rport_io_ins_515 = regs_515_io_out; // @[RegFile.scala 97:16:@50250.4]
  assign rport_io_ins_516 = regs_516_io_out; // @[RegFile.scala 97:16:@50251.4]
  assign rport_io_ins_517 = regs_517_io_out; // @[RegFile.scala 97:16:@50252.4]
  assign rport_io_ins_518 = regs_518_io_out; // @[RegFile.scala 97:16:@50253.4]
  assign rport_io_ins_519 = regs_519_io_out; // @[RegFile.scala 97:16:@50254.4]
  assign rport_io_ins_520 = regs_520_io_out; // @[RegFile.scala 97:16:@50255.4]
  assign rport_io_ins_521 = regs_521_io_out; // @[RegFile.scala 97:16:@50256.4]
  assign rport_io_ins_522 = regs_522_io_out; // @[RegFile.scala 97:16:@50257.4]
  assign rport_io_ins_523 = regs_523_io_out; // @[RegFile.scala 97:16:@50258.4]
  assign rport_io_ins_524 = regs_524_io_out; // @[RegFile.scala 97:16:@50259.4]
  assign rport_io_ins_525 = regs_525_io_out; // @[RegFile.scala 97:16:@50260.4]
  assign rport_io_ins_526 = regs_526_io_out; // @[RegFile.scala 97:16:@50261.4]
  assign rport_io_ins_527 = regs_527_io_out; // @[RegFile.scala 97:16:@50262.4]
  assign rport_io_ins_528 = regs_528_io_out; // @[RegFile.scala 97:16:@50263.4]
  assign rport_io_ins_529 = regs_529_io_out; // @[RegFile.scala 97:16:@50264.4]
  assign rport_io_ins_530 = regs_530_io_out; // @[RegFile.scala 97:16:@50265.4]
  assign rport_io_ins_531 = regs_531_io_out; // @[RegFile.scala 97:16:@50266.4]
  assign rport_io_ins_532 = regs_532_io_out; // @[RegFile.scala 97:16:@50267.4]
  assign rport_io_ins_533 = regs_533_io_out; // @[RegFile.scala 97:16:@50268.4]
  assign rport_io_sel = io_raddr[9:0]; // @[RegFile.scala 106:18:@50269.4]
endmodule
module RetimeWrapper_614( // @[:@50291.2]
  input         clock, // @[:@50292.4]
  input         reset, // @[:@50293.4]
  input  [39:0] io_in, // @[:@50294.4]
  output [39:0] io_out // @[:@50294.4]
);
  wire [39:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@50296.4]
  wire [39:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@50296.4]
  wire [39:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@50296.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@50296.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@50296.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@50296.4]
  RetimeShiftRegister #(.WIDTH(40), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@50296.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@50309.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@50308.4]
  assign sr_init = 40'h0; // @[RetimeShiftRegister.scala 19:16:@50307.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@50306.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@50305.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@50303.4]
endmodule
module FringeFF_534( // @[:@50311.2]
  input         clock, // @[:@50312.4]
  input         reset, // @[:@50313.4]
  input  [39:0] io_in, // @[:@50314.4]
  output [39:0] io_out, // @[:@50314.4]
  input         io_enable // @[:@50314.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@50317.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@50317.4]
  wire [39:0] RetimeWrapper_io_in; // @[package.scala 93:22:@50317.4]
  wire [39:0] RetimeWrapper_io_out; // @[package.scala 93:22:@50317.4]
  wire [39:0] _T_18; // @[package.scala 96:25:@50322.4 package.scala 96:25:@50323.4]
  RetimeWrapper_614 RetimeWrapper ( // @[package.scala 93:22:@50317.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@50322.4 package.scala 96:25:@50323.4]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@50334.4]
  assign RetimeWrapper_clock = clock; // @[:@50318.4]
  assign RetimeWrapper_reset = reset; // @[:@50319.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _T_18; // @[package.scala 94:16:@50320.4]
endmodule
module FringeCounter( // @[:@50336.2]
  input   clock, // @[:@50337.4]
  input   reset, // @[:@50338.4]
  input   io_enable, // @[:@50339.4]
  output  io_done // @[:@50339.4]
);
  wire  reg$_clock; // @[FringeCounter.scala 24:19:@50341.4]
  wire  reg$_reset; // @[FringeCounter.scala 24:19:@50341.4]
  wire [39:0] reg$_io_in; // @[FringeCounter.scala 24:19:@50341.4]
  wire [39:0] reg$_io_out; // @[FringeCounter.scala 24:19:@50341.4]
  wire  reg$_io_enable; // @[FringeCounter.scala 24:19:@50341.4]
  wire [40:0] count; // @[Cat.scala 30:58:@50348.4]
  wire [41:0] _T_25; // @[FringeCounter.scala 31:22:@50349.4]
  wire [40:0] newval; // @[FringeCounter.scala 31:22:@50350.4]
  wire  isMax; // @[FringeCounter.scala 32:22:@50351.4]
  wire [40:0] next; // @[FringeCounter.scala 33:17:@50353.4]
  FringeFF_534 reg$ ( // @[FringeCounter.scala 24:19:@50341.4]
    .clock(reg$_clock),
    .reset(reg$_reset),
    .io_in(reg$_io_in),
    .io_out(reg$_io_out),
    .io_enable(reg$_io_enable)
  );
  assign count = {1'h0,reg$_io_out}; // @[Cat.scala 30:58:@50348.4]
  assign _T_25 = count + 41'h1; // @[FringeCounter.scala 31:22:@50349.4]
  assign newval = count + 41'h1; // @[FringeCounter.scala 31:22:@50350.4]
  assign isMax = newval >= 41'h2cb417800; // @[FringeCounter.scala 32:22:@50351.4]
  assign next = isMax ? count : newval; // @[FringeCounter.scala 33:17:@50353.4]
  assign io_done = io_enable & isMax; // @[FringeCounter.scala 43:11:@50364.4]
  assign reg$_clock = clock; // @[:@50342.4]
  assign reg$_reset = reset; // @[:@50343.4]
  assign reg$_io_in = next[39:0]; // @[FringeCounter.scala 35:15:@50355.6 FringeCounter.scala 37:15:@50358.6]
  assign reg$_io_enable = io_enable; // @[FringeCounter.scala 27:17:@50346.4]
endmodule
module FringeFF_535( // @[:@50398.2]
  input   clock, // @[:@50399.4]
  input   reset, // @[:@50400.4]
  input   io_in, // @[:@50401.4]
  input   io_reset, // @[:@50401.4]
  output  io_out, // @[:@50401.4]
  input   io_enable // @[:@50401.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@50404.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@50404.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@50404.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@50404.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@50404.4]
  wire  _T_18; // @[package.scala 96:25:@50409.4 package.scala 96:25:@50410.4]
  wire  _GEN_0; // @[FringeFF.scala 21:27:@50415.6]
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@50404.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@50409.4 package.scala 96:25:@50410.4]
  assign _GEN_0 = io_reset ? 1'h0 : _T_18; // @[FringeFF.scala 21:27:@50415.6]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@50421.4]
  assign RetimeWrapper_clock = clock; // @[:@50405.4]
  assign RetimeWrapper_reset = reset; // @[:@50406.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@50408.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _GEN_0; // @[package.scala 94:16:@50407.4]
endmodule
module Depulser( // @[:@50423.2]
  input   clock, // @[:@50424.4]
  input   reset, // @[:@50425.4]
  input   io_in, // @[:@50426.4]
  input   io_rst, // @[:@50426.4]
  output  io_out // @[:@50426.4]
);
  wire  r_clock; // @[Depulser.scala 14:17:@50428.4]
  wire  r_reset; // @[Depulser.scala 14:17:@50428.4]
  wire  r_io_in; // @[Depulser.scala 14:17:@50428.4]
  wire  r_io_reset; // @[Depulser.scala 14:17:@50428.4]
  wire  r_io_out; // @[Depulser.scala 14:17:@50428.4]
  wire  r_io_enable; // @[Depulser.scala 14:17:@50428.4]
  FringeFF_535 r ( // @[Depulser.scala 14:17:@50428.4]
    .clock(r_clock),
    .reset(r_reset),
    .io_in(r_io_in),
    .io_reset(r_io_reset),
    .io_out(r_io_out),
    .io_enable(r_io_enable)
  );
  assign io_out = r_io_out; // @[Depulser.scala 19:10:@50437.4]
  assign r_clock = clock; // @[:@50429.4]
  assign r_reset = reset; // @[:@50430.4]
  assign r_io_in = io_rst ? 1'h0 : io_in; // @[Depulser.scala 15:11:@50432.4]
  assign r_io_reset = io_rst; // @[Depulser.scala 18:14:@50436.4]
  assign r_io_enable = io_in | io_rst; // @[Depulser.scala 17:15:@50435.4]
endmodule
module Fringe( // @[:@50439.2]
  input         clock, // @[:@50440.4]
  input         reset, // @[:@50441.4]
  input  [31:0] io_raddr, // @[:@50442.4]
  input         io_wen, // @[:@50442.4]
  input  [31:0] io_waddr, // @[:@50442.4]
  input  [63:0] io_wdata, // @[:@50442.4]
  output [63:0] io_rdata, // @[:@50442.4]
  output        io_enable, // @[:@50442.4]
  input         io_done, // @[:@50442.4]
  output        io_reset, // @[:@50442.4]
  output [63:0] io_argIns_0, // @[:@50442.4]
  input         io_argOuts_0_valid, // @[:@50442.4]
  input  [63:0] io_argOuts_0_bits, // @[:@50442.4]
  input         io_argOuts_1_valid, // @[:@50442.4]
  input  [63:0] io_argOuts_1_bits, // @[:@50442.4]
  input         io_argOuts_2_valid, // @[:@50442.4]
  input  [63:0] io_argOuts_2_bits, // @[:@50442.4]
  input         io_argOuts_3_valid, // @[:@50442.4]
  input  [63:0] io_argOuts_3_bits, // @[:@50442.4]
  input         io_argOuts_4_valid, // @[:@50442.4]
  input  [63:0] io_argOuts_4_bits, // @[:@50442.4]
  input         io_argOuts_5_valid, // @[:@50442.4]
  input  [63:0] io_argOuts_5_bits, // @[:@50442.4]
  input         io_argOuts_6_valid, // @[:@50442.4]
  input  [63:0] io_argOuts_6_bits, // @[:@50442.4]
  input         io_argOuts_7_valid, // @[:@50442.4]
  input  [63:0] io_argOuts_7_bits, // @[:@50442.4]
  input         io_argOuts_8_valid, // @[:@50442.4]
  input  [63:0] io_argOuts_8_bits, // @[:@50442.4]
  input         io_argOuts_9_valid, // @[:@50442.4]
  input  [63:0] io_argOuts_9_bits, // @[:@50442.4]
  input         io_argOuts_10_valid, // @[:@50442.4]
  input  [63:0] io_argOuts_10_bits, // @[:@50442.4]
  input         io_argOuts_11_valid, // @[:@50442.4]
  input  [63:0] io_argOuts_11_bits, // @[:@50442.4]
  input         io_argOuts_12_valid, // @[:@50442.4]
  input  [63:0] io_argOuts_12_bits, // @[:@50442.4]
  input         io_argOuts_13_valid, // @[:@50442.4]
  input  [63:0] io_argOuts_13_bits, // @[:@50442.4]
  input         io_argOuts_14_valid, // @[:@50442.4]
  input  [63:0] io_argOuts_14_bits, // @[:@50442.4]
  input         io_argOuts_15_valid, // @[:@50442.4]
  input  [63:0] io_argOuts_15_bits, // @[:@50442.4]
  input         io_argOuts_16_valid, // @[:@50442.4]
  input  [63:0] io_argOuts_16_bits, // @[:@50442.4]
  input         io_argOuts_17_valid, // @[:@50442.4]
  input  [63:0] io_argOuts_17_bits, // @[:@50442.4]
  input         io_argOuts_18_valid, // @[:@50442.4]
  input  [63:0] io_argOuts_18_bits, // @[:@50442.4]
  input         io_argOuts_19_valid, // @[:@50442.4]
  input  [63:0] io_argOuts_19_bits, // @[:@50442.4]
  input         io_argOuts_20_valid, // @[:@50442.4]
  input  [63:0] io_argOuts_20_bits, // @[:@50442.4]
  input         io_argOuts_21_valid, // @[:@50442.4]
  input  [63:0] io_argOuts_21_bits, // @[:@50442.4]
  input         io_argOuts_22_valid, // @[:@50442.4]
  input  [63:0] io_argOuts_22_bits, // @[:@50442.4]
  input         io_argOuts_23_valid, // @[:@50442.4]
  input  [63:0] io_argOuts_23_bits, // @[:@50442.4]
  input         io_argOuts_24_valid, // @[:@50442.4]
  input  [63:0] io_argOuts_24_bits, // @[:@50442.4]
  input         io_argOuts_25_valid, // @[:@50442.4]
  input  [63:0] io_argOuts_25_bits, // @[:@50442.4]
  input         io_argOuts_26_valid, // @[:@50442.4]
  input  [63:0] io_argOuts_26_bits, // @[:@50442.4]
  input         io_argOuts_27_valid, // @[:@50442.4]
  input  [63:0] io_argOuts_27_bits, // @[:@50442.4]
  input         io_argOuts_28_valid, // @[:@50442.4]
  input  [63:0] io_argOuts_28_bits, // @[:@50442.4]
  input         io_argOuts_29_valid, // @[:@50442.4]
  input  [63:0] io_argOuts_29_bits, // @[:@50442.4]
  input         io_argOuts_30_valid, // @[:@50442.4]
  input  [63:0] io_argOuts_30_bits, // @[:@50442.4]
  input         io_argOuts_31_valid, // @[:@50442.4]
  input  [63:0] io_argOuts_31_bits, // @[:@50442.4]
  input         io_heap_0_req_valid, // @[:@50442.4]
  input         io_heap_0_req_bits_allocDealloc, // @[:@50442.4]
  input  [63:0] io_heap_0_req_bits_sizeAddr, // @[:@50442.4]
  output        io_heap_0_resp_valid, // @[:@50442.4]
  output        io_heap_0_resp_bits_allocDealloc, // @[:@50442.4]
  output [63:0] io_heap_0_resp_bits_sizeAddr // @[:@50442.4]
);
  wire  heap_io_accel_0_req_valid; // @[Fringe.scala 107:20:@51595.4]
  wire  heap_io_accel_0_req_bits_allocDealloc; // @[Fringe.scala 107:20:@51595.4]
  wire [63:0] heap_io_accel_0_req_bits_sizeAddr; // @[Fringe.scala 107:20:@51595.4]
  wire  heap_io_accel_0_resp_valid; // @[Fringe.scala 107:20:@51595.4]
  wire  heap_io_accel_0_resp_bits_allocDealloc; // @[Fringe.scala 107:20:@51595.4]
  wire [63:0] heap_io_accel_0_resp_bits_sizeAddr; // @[Fringe.scala 107:20:@51595.4]
  wire  heap_io_host_0_req_valid; // @[Fringe.scala 107:20:@51595.4]
  wire  heap_io_host_0_req_bits_allocDealloc; // @[Fringe.scala 107:20:@51595.4]
  wire [63:0] heap_io_host_0_req_bits_sizeAddr; // @[Fringe.scala 107:20:@51595.4]
  wire  heap_io_host_0_resp_valid; // @[Fringe.scala 107:20:@51595.4]
  wire  heap_io_host_0_resp_bits_allocDealloc; // @[Fringe.scala 107:20:@51595.4]
  wire [63:0] heap_io_host_0_resp_bits_sizeAddr; // @[Fringe.scala 107:20:@51595.4]
  wire  regs_clock; // @[Fringe.scala 116:20:@51604.4]
  wire  regs_reset; // @[Fringe.scala 116:20:@51604.4]
  wire [31:0] regs_io_raddr; // @[Fringe.scala 116:20:@51604.4]
  wire  regs_io_wen; // @[Fringe.scala 116:20:@51604.4]
  wire [31:0] regs_io_waddr; // @[Fringe.scala 116:20:@51604.4]
  wire [63:0] regs_io_wdata; // @[Fringe.scala 116:20:@51604.4]
  wire [63:0] regs_io_rdata; // @[Fringe.scala 116:20:@51604.4]
  wire  regs_io_reset; // @[Fringe.scala 116:20:@51604.4]
  wire [63:0] regs_io_argIns_0; // @[Fringe.scala 116:20:@51604.4]
  wire [63:0] regs_io_argIns_1; // @[Fringe.scala 116:20:@51604.4]
  wire [63:0] regs_io_argIns_2; // @[Fringe.scala 116:20:@51604.4]
  wire  regs_io_argOuts_0_valid; // @[Fringe.scala 116:20:@51604.4]
  wire [63:0] regs_io_argOuts_0_bits; // @[Fringe.scala 116:20:@51604.4]
  wire  regs_io_argOuts_1_valid; // @[Fringe.scala 116:20:@51604.4]
  wire [63:0] regs_io_argOuts_1_bits; // @[Fringe.scala 116:20:@51604.4]
  wire  regs_io_argOuts_2_valid; // @[Fringe.scala 116:20:@51604.4]
  wire [63:0] regs_io_argOuts_2_bits; // @[Fringe.scala 116:20:@51604.4]
  wire  regs_io_argOuts_3_valid; // @[Fringe.scala 116:20:@51604.4]
  wire [63:0] regs_io_argOuts_3_bits; // @[Fringe.scala 116:20:@51604.4]
  wire  regs_io_argOuts_4_valid; // @[Fringe.scala 116:20:@51604.4]
  wire [63:0] regs_io_argOuts_4_bits; // @[Fringe.scala 116:20:@51604.4]
  wire  regs_io_argOuts_5_valid; // @[Fringe.scala 116:20:@51604.4]
  wire [63:0] regs_io_argOuts_5_bits; // @[Fringe.scala 116:20:@51604.4]
  wire  regs_io_argOuts_6_valid; // @[Fringe.scala 116:20:@51604.4]
  wire [63:0] regs_io_argOuts_6_bits; // @[Fringe.scala 116:20:@51604.4]
  wire  regs_io_argOuts_7_valid; // @[Fringe.scala 116:20:@51604.4]
  wire [63:0] regs_io_argOuts_7_bits; // @[Fringe.scala 116:20:@51604.4]
  wire  regs_io_argOuts_8_valid; // @[Fringe.scala 116:20:@51604.4]
  wire [63:0] regs_io_argOuts_8_bits; // @[Fringe.scala 116:20:@51604.4]
  wire  regs_io_argOuts_9_valid; // @[Fringe.scala 116:20:@51604.4]
  wire [63:0] regs_io_argOuts_9_bits; // @[Fringe.scala 116:20:@51604.4]
  wire  regs_io_argOuts_10_valid; // @[Fringe.scala 116:20:@51604.4]
  wire [63:0] regs_io_argOuts_10_bits; // @[Fringe.scala 116:20:@51604.4]
  wire  regs_io_argOuts_11_valid; // @[Fringe.scala 116:20:@51604.4]
  wire [63:0] regs_io_argOuts_11_bits; // @[Fringe.scala 116:20:@51604.4]
  wire  regs_io_argOuts_12_valid; // @[Fringe.scala 116:20:@51604.4]
  wire [63:0] regs_io_argOuts_12_bits; // @[Fringe.scala 116:20:@51604.4]
  wire  regs_io_argOuts_13_valid; // @[Fringe.scala 116:20:@51604.4]
  wire [63:0] regs_io_argOuts_13_bits; // @[Fringe.scala 116:20:@51604.4]
  wire  regs_io_argOuts_14_valid; // @[Fringe.scala 116:20:@51604.4]
  wire [63:0] regs_io_argOuts_14_bits; // @[Fringe.scala 116:20:@51604.4]
  wire  regs_io_argOuts_15_valid; // @[Fringe.scala 116:20:@51604.4]
  wire [63:0] regs_io_argOuts_15_bits; // @[Fringe.scala 116:20:@51604.4]
  wire  regs_io_argOuts_16_valid; // @[Fringe.scala 116:20:@51604.4]
  wire [63:0] regs_io_argOuts_16_bits; // @[Fringe.scala 116:20:@51604.4]
  wire  regs_io_argOuts_17_valid; // @[Fringe.scala 116:20:@51604.4]
  wire [63:0] regs_io_argOuts_17_bits; // @[Fringe.scala 116:20:@51604.4]
  wire  regs_io_argOuts_18_valid; // @[Fringe.scala 116:20:@51604.4]
  wire [63:0] regs_io_argOuts_18_bits; // @[Fringe.scala 116:20:@51604.4]
  wire  regs_io_argOuts_19_valid; // @[Fringe.scala 116:20:@51604.4]
  wire [63:0] regs_io_argOuts_19_bits; // @[Fringe.scala 116:20:@51604.4]
  wire  regs_io_argOuts_20_valid; // @[Fringe.scala 116:20:@51604.4]
  wire [63:0] regs_io_argOuts_20_bits; // @[Fringe.scala 116:20:@51604.4]
  wire  regs_io_argOuts_21_valid; // @[Fringe.scala 116:20:@51604.4]
  wire [63:0] regs_io_argOuts_21_bits; // @[Fringe.scala 116:20:@51604.4]
  wire  regs_io_argOuts_22_valid; // @[Fringe.scala 116:20:@51604.4]
  wire [63:0] regs_io_argOuts_22_bits; // @[Fringe.scala 116:20:@51604.4]
  wire  regs_io_argOuts_23_valid; // @[Fringe.scala 116:20:@51604.4]
  wire [63:0] regs_io_argOuts_23_bits; // @[Fringe.scala 116:20:@51604.4]
  wire  regs_io_argOuts_24_valid; // @[Fringe.scala 116:20:@51604.4]
  wire [63:0] regs_io_argOuts_24_bits; // @[Fringe.scala 116:20:@51604.4]
  wire  regs_io_argOuts_25_valid; // @[Fringe.scala 116:20:@51604.4]
  wire [63:0] regs_io_argOuts_25_bits; // @[Fringe.scala 116:20:@51604.4]
  wire  regs_io_argOuts_26_valid; // @[Fringe.scala 116:20:@51604.4]
  wire [63:0] regs_io_argOuts_26_bits; // @[Fringe.scala 116:20:@51604.4]
  wire  regs_io_argOuts_27_valid; // @[Fringe.scala 116:20:@51604.4]
  wire [63:0] regs_io_argOuts_27_bits; // @[Fringe.scala 116:20:@51604.4]
  wire  regs_io_argOuts_28_valid; // @[Fringe.scala 116:20:@51604.4]
  wire [63:0] regs_io_argOuts_28_bits; // @[Fringe.scala 116:20:@51604.4]
  wire  regs_io_argOuts_29_valid; // @[Fringe.scala 116:20:@51604.4]
  wire [63:0] regs_io_argOuts_29_bits; // @[Fringe.scala 116:20:@51604.4]
  wire  regs_io_argOuts_30_valid; // @[Fringe.scala 116:20:@51604.4]
  wire [63:0] regs_io_argOuts_30_bits; // @[Fringe.scala 116:20:@51604.4]
  wire  regs_io_argOuts_31_valid; // @[Fringe.scala 116:20:@51604.4]
  wire [63:0] regs_io_argOuts_31_bits; // @[Fringe.scala 116:20:@51604.4]
  wire  regs_io_argOuts_32_valid; // @[Fringe.scala 116:20:@51604.4]
  wire [63:0] regs_io_argOuts_32_bits; // @[Fringe.scala 116:20:@51604.4]
  wire  timeoutCtr_clock; // @[Fringe.scala 143:26:@53777.4]
  wire  timeoutCtr_reset; // @[Fringe.scala 143:26:@53777.4]
  wire  timeoutCtr_io_enable; // @[Fringe.scala 143:26:@53777.4]
  wire  timeoutCtr_io_done; // @[Fringe.scala 143:26:@53777.4]
  wire  depulser_clock; // @[Fringe.scala 153:24:@53795.4]
  wire  depulser_reset; // @[Fringe.scala 153:24:@53795.4]
  wire  depulser_io_in; // @[Fringe.scala 153:24:@53795.4]
  wire  depulser_io_rst; // @[Fringe.scala 153:24:@53795.4]
  wire  depulser_io_out; // @[Fringe.scala 153:24:@53795.4]
  wire [63:0] _T_1012; // @[:@53754.4 :@53755.4]
  wire  curStatus_done; // @[Fringe.scala 133:45:@53756.4]
  wire  curStatus_timeout; // @[Fringe.scala 133:45:@53758.4]
  wire [2:0] curStatus_allocDealloc; // @[Fringe.scala 133:45:@53760.4]
  wire [58:0] curStatus_sizeAddr; // @[Fringe.scala 133:45:@53762.4]
  wire  _T_1017; // @[Fringe.scala 134:28:@53764.4]
  wire  _T_1021; // @[Fringe.scala 134:42:@53766.4]
  wire  _T_1022; // @[Fringe.scala 135:27:@53768.4]
  wire [63:0] _T_1032; // @[Fringe.scala 156:22:@53803.4]
  reg  _T_1039; // @[package.scala 152:20:@53806.4]
  reg [31:0] _RAND_0;
  wire  _T_1040; // @[package.scala 153:13:@53808.4]
  wire  _T_1041; // @[package.scala 153:8:@53809.4]
  wire  _T_1044; // @[Fringe.scala 160:55:@53813.4]
  wire  status_bits_done; // @[Fringe.scala 160:26:@53814.4]
  wire  _T_1047; // @[Fringe.scala 161:58:@53817.4]
  wire  status_bits_timeout; // @[Fringe.scala 161:29:@53818.4]
  wire [1:0] _T_1051; // @[Fringe.scala 162:57:@53820.4]
  wire [1:0] _T_1053; // @[Fringe.scala 162:34:@53821.4]
  wire [63:0] _T_1055; // @[Fringe.scala 163:30:@53823.4]
  wire [1:0] _T_1056; // @[Fringe.scala 171:37:@53826.4]
  wire [58:0] status_bits_sizeAddr; // @[Fringe.scala 158:20:@53805.4 Fringe.scala 163:24:@53824.4]
  wire [2:0] status_bits_allocDealloc; // @[Fringe.scala 158:20:@53805.4 Fringe.scala 162:28:@53822.4]
  wire [61:0] _T_1057; // @[Fringe.scala 171:37:@53827.4]
  wire  alloc; // @[Fringe.scala 202:38:@55205.4]
  wire  dealloc; // @[Fringe.scala 203:40:@55206.4]
  wire  _T_1561; // @[Fringe.scala 204:37:@55207.4]
  reg  _T_1564; // @[package.scala 152:20:@55208.4]
  reg [31:0] _RAND_1;
  wire  _T_1565; // @[package.scala 153:13:@55210.4]
  DRAMHeap heap ( // @[Fringe.scala 107:20:@51595.4]
    .io_accel_0_req_valid(heap_io_accel_0_req_valid),
    .io_accel_0_req_bits_allocDealloc(heap_io_accel_0_req_bits_allocDealloc),
    .io_accel_0_req_bits_sizeAddr(heap_io_accel_0_req_bits_sizeAddr),
    .io_accel_0_resp_valid(heap_io_accel_0_resp_valid),
    .io_accel_0_resp_bits_allocDealloc(heap_io_accel_0_resp_bits_allocDealloc),
    .io_accel_0_resp_bits_sizeAddr(heap_io_accel_0_resp_bits_sizeAddr),
    .io_host_0_req_valid(heap_io_host_0_req_valid),
    .io_host_0_req_bits_allocDealloc(heap_io_host_0_req_bits_allocDealloc),
    .io_host_0_req_bits_sizeAddr(heap_io_host_0_req_bits_sizeAddr),
    .io_host_0_resp_valid(heap_io_host_0_resp_valid),
    .io_host_0_resp_bits_allocDealloc(heap_io_host_0_resp_bits_allocDealloc),
    .io_host_0_resp_bits_sizeAddr(heap_io_host_0_resp_bits_sizeAddr)
  );
  RegFile regs ( // @[Fringe.scala 116:20:@51604.4]
    .clock(regs_clock),
    .reset(regs_reset),
    .io_raddr(regs_io_raddr),
    .io_wen(regs_io_wen),
    .io_waddr(regs_io_waddr),
    .io_wdata(regs_io_wdata),
    .io_rdata(regs_io_rdata),
    .io_reset(regs_io_reset),
    .io_argIns_0(regs_io_argIns_0),
    .io_argIns_1(regs_io_argIns_1),
    .io_argIns_2(regs_io_argIns_2),
    .io_argOuts_0_valid(regs_io_argOuts_0_valid),
    .io_argOuts_0_bits(regs_io_argOuts_0_bits),
    .io_argOuts_1_valid(regs_io_argOuts_1_valid),
    .io_argOuts_1_bits(regs_io_argOuts_1_bits),
    .io_argOuts_2_valid(regs_io_argOuts_2_valid),
    .io_argOuts_2_bits(regs_io_argOuts_2_bits),
    .io_argOuts_3_valid(regs_io_argOuts_3_valid),
    .io_argOuts_3_bits(regs_io_argOuts_3_bits),
    .io_argOuts_4_valid(regs_io_argOuts_4_valid),
    .io_argOuts_4_bits(regs_io_argOuts_4_bits),
    .io_argOuts_5_valid(regs_io_argOuts_5_valid),
    .io_argOuts_5_bits(regs_io_argOuts_5_bits),
    .io_argOuts_6_valid(regs_io_argOuts_6_valid),
    .io_argOuts_6_bits(regs_io_argOuts_6_bits),
    .io_argOuts_7_valid(regs_io_argOuts_7_valid),
    .io_argOuts_7_bits(regs_io_argOuts_7_bits),
    .io_argOuts_8_valid(regs_io_argOuts_8_valid),
    .io_argOuts_8_bits(regs_io_argOuts_8_bits),
    .io_argOuts_9_valid(regs_io_argOuts_9_valid),
    .io_argOuts_9_bits(regs_io_argOuts_9_bits),
    .io_argOuts_10_valid(regs_io_argOuts_10_valid),
    .io_argOuts_10_bits(regs_io_argOuts_10_bits),
    .io_argOuts_11_valid(regs_io_argOuts_11_valid),
    .io_argOuts_11_bits(regs_io_argOuts_11_bits),
    .io_argOuts_12_valid(regs_io_argOuts_12_valid),
    .io_argOuts_12_bits(regs_io_argOuts_12_bits),
    .io_argOuts_13_valid(regs_io_argOuts_13_valid),
    .io_argOuts_13_bits(regs_io_argOuts_13_bits),
    .io_argOuts_14_valid(regs_io_argOuts_14_valid),
    .io_argOuts_14_bits(regs_io_argOuts_14_bits),
    .io_argOuts_15_valid(regs_io_argOuts_15_valid),
    .io_argOuts_15_bits(regs_io_argOuts_15_bits),
    .io_argOuts_16_valid(regs_io_argOuts_16_valid),
    .io_argOuts_16_bits(regs_io_argOuts_16_bits),
    .io_argOuts_17_valid(regs_io_argOuts_17_valid),
    .io_argOuts_17_bits(regs_io_argOuts_17_bits),
    .io_argOuts_18_valid(regs_io_argOuts_18_valid),
    .io_argOuts_18_bits(regs_io_argOuts_18_bits),
    .io_argOuts_19_valid(regs_io_argOuts_19_valid),
    .io_argOuts_19_bits(regs_io_argOuts_19_bits),
    .io_argOuts_20_valid(regs_io_argOuts_20_valid),
    .io_argOuts_20_bits(regs_io_argOuts_20_bits),
    .io_argOuts_21_valid(regs_io_argOuts_21_valid),
    .io_argOuts_21_bits(regs_io_argOuts_21_bits),
    .io_argOuts_22_valid(regs_io_argOuts_22_valid),
    .io_argOuts_22_bits(regs_io_argOuts_22_bits),
    .io_argOuts_23_valid(regs_io_argOuts_23_valid),
    .io_argOuts_23_bits(regs_io_argOuts_23_bits),
    .io_argOuts_24_valid(regs_io_argOuts_24_valid),
    .io_argOuts_24_bits(regs_io_argOuts_24_bits),
    .io_argOuts_25_valid(regs_io_argOuts_25_valid),
    .io_argOuts_25_bits(regs_io_argOuts_25_bits),
    .io_argOuts_26_valid(regs_io_argOuts_26_valid),
    .io_argOuts_26_bits(regs_io_argOuts_26_bits),
    .io_argOuts_27_valid(regs_io_argOuts_27_valid),
    .io_argOuts_27_bits(regs_io_argOuts_27_bits),
    .io_argOuts_28_valid(regs_io_argOuts_28_valid),
    .io_argOuts_28_bits(regs_io_argOuts_28_bits),
    .io_argOuts_29_valid(regs_io_argOuts_29_valid),
    .io_argOuts_29_bits(regs_io_argOuts_29_bits),
    .io_argOuts_30_valid(regs_io_argOuts_30_valid),
    .io_argOuts_30_bits(regs_io_argOuts_30_bits),
    .io_argOuts_31_valid(regs_io_argOuts_31_valid),
    .io_argOuts_31_bits(regs_io_argOuts_31_bits),
    .io_argOuts_32_valid(regs_io_argOuts_32_valid),
    .io_argOuts_32_bits(regs_io_argOuts_32_bits)
  );
  FringeCounter timeoutCtr ( // @[Fringe.scala 143:26:@53777.4]
    .clock(timeoutCtr_clock),
    .reset(timeoutCtr_reset),
    .io_enable(timeoutCtr_io_enable),
    .io_done(timeoutCtr_io_done)
  );
  Depulser depulser ( // @[Fringe.scala 153:24:@53795.4]
    .clock(depulser_clock),
    .reset(depulser_reset),
    .io_in(depulser_io_in),
    .io_rst(depulser_io_rst),
    .io_out(depulser_io_out)
  );
  assign _T_1012 = regs_io_argIns_1; // @[:@53754.4 :@53755.4]
  assign curStatus_done = _T_1012[0]; // @[Fringe.scala 133:45:@53756.4]
  assign curStatus_timeout = _T_1012[1]; // @[Fringe.scala 133:45:@53758.4]
  assign curStatus_allocDealloc = _T_1012[4:2]; // @[Fringe.scala 133:45:@53760.4]
  assign curStatus_sizeAddr = _T_1012[63:5]; // @[Fringe.scala 133:45:@53762.4]
  assign _T_1017 = regs_io_argIns_0[0]; // @[Fringe.scala 134:28:@53764.4]
  assign _T_1021 = curStatus_done == 1'h0; // @[Fringe.scala 134:42:@53766.4]
  assign _T_1022 = regs_io_argIns_0[1]; // @[Fringe.scala 135:27:@53768.4]
  assign _T_1032 = ~ regs_io_argIns_0; // @[Fringe.scala 156:22:@53803.4]
  assign _T_1040 = _T_1039 ^ heap_io_host_0_req_valid; // @[package.scala 153:13:@53808.4]
  assign _T_1041 = heap_io_host_0_req_valid & _T_1040; // @[package.scala 153:8:@53809.4]
  assign _T_1044 = _T_1017 & depulser_io_out; // @[Fringe.scala 160:55:@53813.4]
  assign status_bits_done = depulser_io_out ? _T_1044 : curStatus_done; // @[Fringe.scala 160:26:@53814.4]
  assign _T_1047 = _T_1017 & timeoutCtr_io_done; // @[Fringe.scala 161:58:@53817.4]
  assign status_bits_timeout = depulser_io_out ? _T_1047 : curStatus_timeout; // @[Fringe.scala 161:29:@53818.4]
  assign _T_1051 = heap_io_host_0_req_bits_allocDealloc ? 2'h1 : 2'h2; // @[Fringe.scala 162:57:@53820.4]
  assign _T_1053 = heap_io_host_0_req_valid ? _T_1051 : 2'h0; // @[Fringe.scala 162:34:@53821.4]
  assign _T_1055 = heap_io_host_0_req_valid ? heap_io_host_0_req_bits_sizeAddr : 64'h0; // @[Fringe.scala 163:30:@53823.4]
  assign _T_1056 = {status_bits_timeout,status_bits_done}; // @[Fringe.scala 171:37:@53826.4]
  assign status_bits_sizeAddr = _T_1055[58:0]; // @[Fringe.scala 158:20:@53805.4 Fringe.scala 163:24:@53824.4]
  assign status_bits_allocDealloc = {{1'd0}, _T_1053}; // @[Fringe.scala 158:20:@53805.4 Fringe.scala 162:28:@53822.4]
  assign _T_1057 = {status_bits_sizeAddr,status_bits_allocDealloc}; // @[Fringe.scala 171:37:@53827.4]
  assign alloc = curStatus_allocDealloc == 3'h3; // @[Fringe.scala 202:38:@55205.4]
  assign dealloc = curStatus_allocDealloc == 3'h4; // @[Fringe.scala 203:40:@55206.4]
  assign _T_1561 = alloc | dealloc; // @[Fringe.scala 204:37:@55207.4]
  assign _T_1565 = _T_1564 ^ _T_1561; // @[package.scala 153:13:@55210.4]
  assign io_rdata = regs_io_rdata; // @[Fringe.scala 125:14:@53752.4]
  assign io_enable = _T_1017 & _T_1021; // @[Fringe.scala 136:13:@53772.4]
  assign io_reset = _T_1022 | reset; // @[Fringe.scala 137:12:@53773.4]
  assign io_argIns_0 = regs_io_argIns_2; // @[Fringe.scala 151:51:@53794.4]
  assign io_heap_0_resp_valid = heap_io_accel_0_resp_valid; // @[Fringe.scala 108:17:@51600.4]
  assign io_heap_0_resp_bits_allocDealloc = heap_io_accel_0_resp_bits_allocDealloc; // @[Fringe.scala 108:17:@51599.4]
  assign io_heap_0_resp_bits_sizeAddr = heap_io_accel_0_resp_bits_sizeAddr; // @[Fringe.scala 108:17:@51598.4]
  assign heap_io_accel_0_req_valid = io_heap_0_req_valid; // @[Fringe.scala 108:17:@51603.4]
  assign heap_io_accel_0_req_bits_allocDealloc = io_heap_0_req_bits_allocDealloc; // @[Fringe.scala 108:17:@51602.4]
  assign heap_io_accel_0_req_bits_sizeAddr = io_heap_0_req_bits_sizeAddr; // @[Fringe.scala 108:17:@51601.4]
  assign heap_io_host_0_resp_valid = _T_1561 & _T_1565; // @[Fringe.scala 204:22:@55212.4]
  assign heap_io_host_0_resp_bits_allocDealloc = curStatus_allocDealloc == 3'h3; // @[Fringe.scala 205:34:@55213.4]
  assign heap_io_host_0_resp_bits_sizeAddr = {{5'd0}, curStatus_sizeAddr}; // @[Fringe.scala 206:30:@55214.4]
  assign regs_clock = clock; // @[:@51605.4]
  assign regs_reset = reset; // @[:@51606.4 Fringe.scala 139:14:@53776.4]
  assign regs_io_raddr = io_raddr; // @[Fringe.scala 118:17:@53748.4]
  assign regs_io_wen = io_wen; // @[Fringe.scala 120:15:@53750.4]
  assign regs_io_waddr = io_waddr; // @[Fringe.scala 119:17:@53749.4]
  assign regs_io_wdata = io_wdata; // @[Fringe.scala 121:17:@53751.4]
  assign regs_io_reset = _T_1022 | reset; // @[Fringe.scala 138:17:@53774.4]
  assign regs_io_argOuts_0_valid = depulser_io_out | _T_1041; // @[Fringe.scala 170:23:@53825.4]
  assign regs_io_argOuts_0_bits = {_T_1057,_T_1056}; // @[Fringe.scala 171:22:@53829.4]
  assign regs_io_argOuts_1_valid = io_argOuts_0_valid; // @[Fringe.scala 176:23:@53832.4]
  assign regs_io_argOuts_1_bits = io_argOuts_0_bits; // @[Fringe.scala 175:22:@53831.4]
  assign regs_io_argOuts_2_valid = io_argOuts_1_valid; // @[Fringe.scala 176:23:@53835.4]
  assign regs_io_argOuts_2_bits = io_argOuts_1_bits; // @[Fringe.scala 175:22:@53834.4]
  assign regs_io_argOuts_3_valid = io_argOuts_2_valid; // @[Fringe.scala 176:23:@53838.4]
  assign regs_io_argOuts_3_bits = io_argOuts_2_bits; // @[Fringe.scala 175:22:@53837.4]
  assign regs_io_argOuts_4_valid = io_argOuts_3_valid; // @[Fringe.scala 176:23:@53841.4]
  assign regs_io_argOuts_4_bits = io_argOuts_3_bits; // @[Fringe.scala 175:22:@53840.4]
  assign regs_io_argOuts_5_valid = io_argOuts_4_valid; // @[Fringe.scala 176:23:@53844.4]
  assign regs_io_argOuts_5_bits = io_argOuts_4_bits; // @[Fringe.scala 175:22:@53843.4]
  assign regs_io_argOuts_6_valid = io_argOuts_5_valid; // @[Fringe.scala 176:23:@53847.4]
  assign regs_io_argOuts_6_bits = io_argOuts_5_bits; // @[Fringe.scala 175:22:@53846.4]
  assign regs_io_argOuts_7_valid = io_argOuts_6_valid; // @[Fringe.scala 176:23:@53850.4]
  assign regs_io_argOuts_7_bits = io_argOuts_6_bits; // @[Fringe.scala 175:22:@53849.4]
  assign regs_io_argOuts_8_valid = io_argOuts_7_valid; // @[Fringe.scala 176:23:@53853.4]
  assign regs_io_argOuts_8_bits = io_argOuts_7_bits; // @[Fringe.scala 175:22:@53852.4]
  assign regs_io_argOuts_9_valid = io_argOuts_8_valid; // @[Fringe.scala 176:23:@53856.4]
  assign regs_io_argOuts_9_bits = io_argOuts_8_bits; // @[Fringe.scala 175:22:@53855.4]
  assign regs_io_argOuts_10_valid = io_argOuts_9_valid; // @[Fringe.scala 176:23:@53859.4]
  assign regs_io_argOuts_10_bits = io_argOuts_9_bits; // @[Fringe.scala 175:22:@53858.4]
  assign regs_io_argOuts_11_valid = io_argOuts_10_valid; // @[Fringe.scala 176:23:@53862.4]
  assign regs_io_argOuts_11_bits = io_argOuts_10_bits; // @[Fringe.scala 175:22:@53861.4]
  assign regs_io_argOuts_12_valid = io_argOuts_11_valid; // @[Fringe.scala 176:23:@53865.4]
  assign regs_io_argOuts_12_bits = io_argOuts_11_bits; // @[Fringe.scala 175:22:@53864.4]
  assign regs_io_argOuts_13_valid = io_argOuts_12_valid; // @[Fringe.scala 176:23:@53868.4]
  assign regs_io_argOuts_13_bits = io_argOuts_12_bits; // @[Fringe.scala 175:22:@53867.4]
  assign regs_io_argOuts_14_valid = io_argOuts_13_valid; // @[Fringe.scala 176:23:@53871.4]
  assign regs_io_argOuts_14_bits = io_argOuts_13_bits; // @[Fringe.scala 175:22:@53870.4]
  assign regs_io_argOuts_15_valid = io_argOuts_14_valid; // @[Fringe.scala 176:23:@53874.4]
  assign regs_io_argOuts_15_bits = io_argOuts_14_bits; // @[Fringe.scala 175:22:@53873.4]
  assign regs_io_argOuts_16_valid = io_argOuts_15_valid; // @[Fringe.scala 176:23:@53877.4]
  assign regs_io_argOuts_16_bits = io_argOuts_15_bits; // @[Fringe.scala 175:22:@53876.4]
  assign regs_io_argOuts_17_valid = io_argOuts_16_valid; // @[Fringe.scala 176:23:@53880.4]
  assign regs_io_argOuts_17_bits = io_argOuts_16_bits; // @[Fringe.scala 175:22:@53879.4]
  assign regs_io_argOuts_18_valid = io_argOuts_17_valid; // @[Fringe.scala 176:23:@53883.4]
  assign regs_io_argOuts_18_bits = io_argOuts_17_bits; // @[Fringe.scala 175:22:@53882.4]
  assign regs_io_argOuts_19_valid = io_argOuts_18_valid; // @[Fringe.scala 176:23:@53886.4]
  assign regs_io_argOuts_19_bits = io_argOuts_18_bits; // @[Fringe.scala 175:22:@53885.4]
  assign regs_io_argOuts_20_valid = io_argOuts_19_valid; // @[Fringe.scala 176:23:@53889.4]
  assign regs_io_argOuts_20_bits = io_argOuts_19_bits; // @[Fringe.scala 175:22:@53888.4]
  assign regs_io_argOuts_21_valid = io_argOuts_20_valid; // @[Fringe.scala 176:23:@53892.4]
  assign regs_io_argOuts_21_bits = io_argOuts_20_bits; // @[Fringe.scala 175:22:@53891.4]
  assign regs_io_argOuts_22_valid = io_argOuts_21_valid; // @[Fringe.scala 176:23:@53895.4]
  assign regs_io_argOuts_22_bits = io_argOuts_21_bits; // @[Fringe.scala 175:22:@53894.4]
  assign regs_io_argOuts_23_valid = io_argOuts_22_valid; // @[Fringe.scala 176:23:@53898.4]
  assign regs_io_argOuts_23_bits = io_argOuts_22_bits; // @[Fringe.scala 175:22:@53897.4]
  assign regs_io_argOuts_24_valid = io_argOuts_23_valid; // @[Fringe.scala 176:23:@53901.4]
  assign regs_io_argOuts_24_bits = io_argOuts_23_bits; // @[Fringe.scala 175:22:@53900.4]
  assign regs_io_argOuts_25_valid = io_argOuts_24_valid; // @[Fringe.scala 176:23:@53904.4]
  assign regs_io_argOuts_25_bits = io_argOuts_24_bits; // @[Fringe.scala 175:22:@53903.4]
  assign regs_io_argOuts_26_valid = io_argOuts_25_valid; // @[Fringe.scala 176:23:@53907.4]
  assign regs_io_argOuts_26_bits = io_argOuts_25_bits; // @[Fringe.scala 175:22:@53906.4]
  assign regs_io_argOuts_27_valid = io_argOuts_26_valid; // @[Fringe.scala 176:23:@53910.4]
  assign regs_io_argOuts_27_bits = io_argOuts_26_bits; // @[Fringe.scala 175:22:@53909.4]
  assign regs_io_argOuts_28_valid = io_argOuts_27_valid; // @[Fringe.scala 176:23:@53913.4]
  assign regs_io_argOuts_28_bits = io_argOuts_27_bits; // @[Fringe.scala 175:22:@53912.4]
  assign regs_io_argOuts_29_valid = io_argOuts_28_valid; // @[Fringe.scala 176:23:@53916.4]
  assign regs_io_argOuts_29_bits = io_argOuts_28_bits; // @[Fringe.scala 175:22:@53915.4]
  assign regs_io_argOuts_30_valid = io_argOuts_29_valid; // @[Fringe.scala 176:23:@53919.4]
  assign regs_io_argOuts_30_bits = io_argOuts_29_bits; // @[Fringe.scala 175:22:@53918.4]
  assign regs_io_argOuts_31_valid = io_argOuts_30_valid; // @[Fringe.scala 176:23:@53922.4]
  assign regs_io_argOuts_31_bits = io_argOuts_30_bits; // @[Fringe.scala 175:22:@53921.4]
  assign regs_io_argOuts_32_valid = io_argOuts_31_valid; // @[Fringe.scala 176:23:@53925.4]
  assign regs_io_argOuts_32_bits = io_argOuts_31_bits; // @[Fringe.scala 175:22:@53924.4]
  assign timeoutCtr_clock = clock; // @[:@53778.4]
  assign timeoutCtr_reset = reset; // @[:@53779.4]
  assign timeoutCtr_io_enable = _T_1017 & _T_1021; // @[Fringe.scala 149:24:@53793.4]
  assign depulser_clock = clock; // @[:@53796.4]
  assign depulser_reset = reset; // @[:@53797.4]
  assign depulser_io_in = io_done | timeoutCtr_io_done; // @[Fringe.scala 155:18:@53802.4]
  assign depulser_io_rst = _T_1032[0]; // @[Fringe.scala 156:19:@53804.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1039 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1564 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_1039 <= 1'h0;
    end else begin
      _T_1039 <= heap_io_host_0_req_valid;
    end
    if (reset) begin
      _T_1564 <= 1'h0;
    end else begin
      _T_1564 <= _T_1561;
    end
  end
endmodule
module AXI4LiteToRFBridgeKCU1500( // @[:@55229.2]
  input         clock, // @[:@55230.4]
  input         reset, // @[:@55231.4]
  input  [31:0] io_S_AXI_AWADDR, // @[:@55232.4]
  input  [2:0]  io_S_AXI_AWPROT, // @[:@55232.4]
  input         io_S_AXI_AWVALID, // @[:@55232.4]
  output        io_S_AXI_AWREADY, // @[:@55232.4]
  input  [31:0] io_S_AXI_ARADDR, // @[:@55232.4]
  input  [2:0]  io_S_AXI_ARPROT, // @[:@55232.4]
  input         io_S_AXI_ARVALID, // @[:@55232.4]
  output        io_S_AXI_ARREADY, // @[:@55232.4]
  input  [31:0] io_S_AXI_WDATA, // @[:@55232.4]
  input  [3:0]  io_S_AXI_WSTRB, // @[:@55232.4]
  input         io_S_AXI_WVALID, // @[:@55232.4]
  output        io_S_AXI_WREADY, // @[:@55232.4]
  output [31:0] io_S_AXI_RDATA, // @[:@55232.4]
  output [1:0]  io_S_AXI_RRESP, // @[:@55232.4]
  output        io_S_AXI_RVALID, // @[:@55232.4]
  input         io_S_AXI_RREADY, // @[:@55232.4]
  output [1:0]  io_S_AXI_BRESP, // @[:@55232.4]
  output        io_S_AXI_BVALID, // @[:@55232.4]
  input         io_S_AXI_BREADY, // @[:@55232.4]
  output [31:0] io_raddr, // @[:@55232.4]
  output        io_wen, // @[:@55232.4]
  output [31:0] io_waddr, // @[:@55232.4]
  output [31:0] io_wdata, // @[:@55232.4]
  input  [31:0] io_rdata // @[:@55232.4]
);
  wire [31:0] d_rf_rdata; // @[AXI4LiteToRFBridge.scala 109:17:@55234.4]
  wire [31:0] d_rf_wdata; // @[AXI4LiteToRFBridge.scala 109:17:@55234.4]
  wire [31:0] d_rf_waddr; // @[AXI4LiteToRFBridge.scala 109:17:@55234.4]
  wire  d_rf_wen; // @[AXI4LiteToRFBridge.scala 109:17:@55234.4]
  wire [31:0] d_rf_raddr; // @[AXI4LiteToRFBridge.scala 109:17:@55234.4]
  wire  d_S_AXI_ARESETN; // @[AXI4LiteToRFBridge.scala 109:17:@55234.4]
  wire  d_S_AXI_ACLK; // @[AXI4LiteToRFBridge.scala 109:17:@55234.4]
  wire [31:0] d_S_AXI_AWADDR; // @[AXI4LiteToRFBridge.scala 109:17:@55234.4]
  wire [2:0] d_S_AXI_AWPROT; // @[AXI4LiteToRFBridge.scala 109:17:@55234.4]
  wire  d_S_AXI_AWVALID; // @[AXI4LiteToRFBridge.scala 109:17:@55234.4]
  wire  d_S_AXI_AWREADY; // @[AXI4LiteToRFBridge.scala 109:17:@55234.4]
  wire [31:0] d_S_AXI_ARADDR; // @[AXI4LiteToRFBridge.scala 109:17:@55234.4]
  wire [2:0] d_S_AXI_ARPROT; // @[AXI4LiteToRFBridge.scala 109:17:@55234.4]
  wire  d_S_AXI_ARVALID; // @[AXI4LiteToRFBridge.scala 109:17:@55234.4]
  wire  d_S_AXI_ARREADY; // @[AXI4LiteToRFBridge.scala 109:17:@55234.4]
  wire [31:0] d_S_AXI_WDATA; // @[AXI4LiteToRFBridge.scala 109:17:@55234.4]
  wire [3:0] d_S_AXI_WSTRB; // @[AXI4LiteToRFBridge.scala 109:17:@55234.4]
  wire  d_S_AXI_WVALID; // @[AXI4LiteToRFBridge.scala 109:17:@55234.4]
  wire  d_S_AXI_WREADY; // @[AXI4LiteToRFBridge.scala 109:17:@55234.4]
  wire [31:0] d_S_AXI_RDATA; // @[AXI4LiteToRFBridge.scala 109:17:@55234.4]
  wire [1:0] d_S_AXI_RRESP; // @[AXI4LiteToRFBridge.scala 109:17:@55234.4]
  wire  d_S_AXI_RVALID; // @[AXI4LiteToRFBridge.scala 109:17:@55234.4]
  wire  d_S_AXI_RREADY; // @[AXI4LiteToRFBridge.scala 109:17:@55234.4]
  wire [1:0] d_S_AXI_BRESP; // @[AXI4LiteToRFBridge.scala 109:17:@55234.4]
  wire  d_S_AXI_BVALID; // @[AXI4LiteToRFBridge.scala 109:17:@55234.4]
  wire  d_S_AXI_BREADY; // @[AXI4LiteToRFBridge.scala 109:17:@55234.4]
  AXI4LiteToRFBridgeVerilog d ( // @[AXI4LiteToRFBridge.scala 109:17:@55234.4]
    .rf_rdata(d_rf_rdata),
    .rf_wdata(d_rf_wdata),
    .rf_waddr(d_rf_waddr),
    .rf_wen(d_rf_wen),
    .rf_raddr(d_rf_raddr),
    .S_AXI_ARESETN(d_S_AXI_ARESETN),
    .S_AXI_ACLK(d_S_AXI_ACLK),
    .S_AXI_AWADDR(d_S_AXI_AWADDR),
    .S_AXI_AWPROT(d_S_AXI_AWPROT),
    .S_AXI_AWVALID(d_S_AXI_AWVALID),
    .S_AXI_AWREADY(d_S_AXI_AWREADY),
    .S_AXI_ARADDR(d_S_AXI_ARADDR),
    .S_AXI_ARPROT(d_S_AXI_ARPROT),
    .S_AXI_ARVALID(d_S_AXI_ARVALID),
    .S_AXI_ARREADY(d_S_AXI_ARREADY),
    .S_AXI_WDATA(d_S_AXI_WDATA),
    .S_AXI_WSTRB(d_S_AXI_WSTRB),
    .S_AXI_WVALID(d_S_AXI_WVALID),
    .S_AXI_WREADY(d_S_AXI_WREADY),
    .S_AXI_RDATA(d_S_AXI_RDATA),
    .S_AXI_RRESP(d_S_AXI_RRESP),
    .S_AXI_RVALID(d_S_AXI_RVALID),
    .S_AXI_RREADY(d_S_AXI_RREADY),
    .S_AXI_BRESP(d_S_AXI_BRESP),
    .S_AXI_BVALID(d_S_AXI_BVALID),
    .S_AXI_BREADY(d_S_AXI_BREADY)
  );
  assign io_S_AXI_AWREADY = d_S_AXI_AWREADY; // @[AXI4LiteToRFBridge.scala 111:14:@55258.4]
  assign io_S_AXI_ARREADY = d_S_AXI_ARREADY; // @[AXI4LiteToRFBridge.scala 111:14:@55254.4]
  assign io_S_AXI_WREADY = d_S_AXI_WREADY; // @[AXI4LiteToRFBridge.scala 111:14:@55250.4]
  assign io_S_AXI_RDATA = d_S_AXI_RDATA; // @[AXI4LiteToRFBridge.scala 111:14:@55249.4]
  assign io_S_AXI_RRESP = d_S_AXI_RRESP; // @[AXI4LiteToRFBridge.scala 111:14:@55248.4]
  assign io_S_AXI_RVALID = d_S_AXI_RVALID; // @[AXI4LiteToRFBridge.scala 111:14:@55247.4]
  assign io_S_AXI_BRESP = d_S_AXI_BRESP; // @[AXI4LiteToRFBridge.scala 111:14:@55245.4]
  assign io_S_AXI_BVALID = d_S_AXI_BVALID; // @[AXI4LiteToRFBridge.scala 111:14:@55244.4]
  assign io_raddr = d_rf_raddr; // @[AXI4LiteToRFBridge.scala 115:12:@55266.4]
  assign io_wen = d_rf_wen; // @[AXI4LiteToRFBridge.scala 118:12:@55269.4]
  assign io_waddr = d_rf_waddr; // @[AXI4LiteToRFBridge.scala 116:12:@55267.4]
  assign io_wdata = d_rf_wdata; // @[AXI4LiteToRFBridge.scala 117:12:@55268.4]
  assign d_rf_rdata = io_rdata; // @[AXI4LiteToRFBridge.scala 119:17:@55270.4]
  assign d_S_AXI_ARESETN = ~ reset; // @[AXI4LiteToRFBridge.scala 113:22:@55265.4]
  assign d_S_AXI_ACLK = clock; // @[AXI4LiteToRFBridge.scala 112:19:@55262.4]
  assign d_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[AXI4LiteToRFBridge.scala 111:14:@55261.4]
  assign d_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[AXI4LiteToRFBridge.scala 111:14:@55260.4]
  assign d_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[AXI4LiteToRFBridge.scala 111:14:@55259.4]
  assign d_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[AXI4LiteToRFBridge.scala 111:14:@55257.4]
  assign d_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[AXI4LiteToRFBridge.scala 111:14:@55256.4]
  assign d_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[AXI4LiteToRFBridge.scala 111:14:@55255.4]
  assign d_S_AXI_WDATA = io_S_AXI_WDATA; // @[AXI4LiteToRFBridge.scala 111:14:@55253.4]
  assign d_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[AXI4LiteToRFBridge.scala 111:14:@55252.4]
  assign d_S_AXI_WVALID = io_S_AXI_WVALID; // @[AXI4LiteToRFBridge.scala 111:14:@55251.4]
  assign d_S_AXI_RREADY = io_S_AXI_RREADY; // @[AXI4LiteToRFBridge.scala 111:14:@55246.4]
  assign d_S_AXI_BREADY = io_S_AXI_BREADY; // @[AXI4LiteToRFBridge.scala 111:14:@55243.4]
endmodule
module MAGToAXI4Bridge( // @[:@55272.2]
  output [7:0] io_M_AXI_AWLEN, // @[:@55275.4]
  output [7:0] io_M_AXI_ARLEN // @[:@55275.4]
);
  wire [32:0] _T_218; // @[MAGToAXI4Bridge.scala 27:29:@55432.4]
  wire [32:0] _T_219; // @[MAGToAXI4Bridge.scala 27:29:@55433.4]
  wire [31:0] _T_220; // @[MAGToAXI4Bridge.scala 27:29:@55434.4]
  assign _T_218 = 32'h0 - 32'h1; // @[MAGToAXI4Bridge.scala 27:29:@55432.4]
  assign _T_219 = $unsigned(_T_218); // @[MAGToAXI4Bridge.scala 27:29:@55433.4]
  assign _T_220 = _T_219[31:0]; // @[MAGToAXI4Bridge.scala 27:29:@55434.4]
  assign io_M_AXI_AWLEN = _T_220[7:0]; // @[MAGToAXI4Bridge.scala 41:21:@55452.4]
  assign io_M_AXI_ARLEN = _T_220[7:0]; // @[MAGToAXI4Bridge.scala 27:21:@55435.4]
endmodule
module FringeZynq( // @[:@55600.2]
  input         clock, // @[:@55601.4]
  input         reset, // @[:@55602.4]
  input  [31:0] io_S_AXI_AWADDR, // @[:@55603.4]
  input  [2:0]  io_S_AXI_AWPROT, // @[:@55603.4]
  input         io_S_AXI_AWVALID, // @[:@55603.4]
  output        io_S_AXI_AWREADY, // @[:@55603.4]
  input  [31:0] io_S_AXI_ARADDR, // @[:@55603.4]
  input  [2:0]  io_S_AXI_ARPROT, // @[:@55603.4]
  input         io_S_AXI_ARVALID, // @[:@55603.4]
  output        io_S_AXI_ARREADY, // @[:@55603.4]
  input  [31:0] io_S_AXI_WDATA, // @[:@55603.4]
  input  [3:0]  io_S_AXI_WSTRB, // @[:@55603.4]
  input         io_S_AXI_WVALID, // @[:@55603.4]
  output        io_S_AXI_WREADY, // @[:@55603.4]
  output [31:0] io_S_AXI_RDATA, // @[:@55603.4]
  output [1:0]  io_S_AXI_RRESP, // @[:@55603.4]
  output        io_S_AXI_RVALID, // @[:@55603.4]
  input         io_S_AXI_RREADY, // @[:@55603.4]
  output [1:0]  io_S_AXI_BRESP, // @[:@55603.4]
  output        io_S_AXI_BVALID, // @[:@55603.4]
  input         io_S_AXI_BREADY, // @[:@55603.4]
  output [7:0]  io_M_AXI_0_AWLEN, // @[:@55603.4]
  output [7:0]  io_M_AXI_0_ARLEN, // @[:@55603.4]
  output        io_enable, // @[:@55603.4]
  input         io_done, // @[:@55603.4]
  output        io_reset, // @[:@55603.4]
  output [63:0] io_argIns_0, // @[:@55603.4]
  input         io_argOuts_0_valid, // @[:@55603.4]
  input  [63:0] io_argOuts_0_bits, // @[:@55603.4]
  input         io_argOuts_1_valid, // @[:@55603.4]
  input  [63:0] io_argOuts_1_bits, // @[:@55603.4]
  input         io_argOuts_2_valid, // @[:@55603.4]
  input  [63:0] io_argOuts_2_bits, // @[:@55603.4]
  input         io_argOuts_3_valid, // @[:@55603.4]
  input  [63:0] io_argOuts_3_bits, // @[:@55603.4]
  input         io_argOuts_4_valid, // @[:@55603.4]
  input  [63:0] io_argOuts_4_bits, // @[:@55603.4]
  input         io_argOuts_5_valid, // @[:@55603.4]
  input  [63:0] io_argOuts_5_bits, // @[:@55603.4]
  input         io_argOuts_6_valid, // @[:@55603.4]
  input  [63:0] io_argOuts_6_bits, // @[:@55603.4]
  input         io_argOuts_7_valid, // @[:@55603.4]
  input  [63:0] io_argOuts_7_bits, // @[:@55603.4]
  input         io_argOuts_8_valid, // @[:@55603.4]
  input  [63:0] io_argOuts_8_bits, // @[:@55603.4]
  input         io_argOuts_9_valid, // @[:@55603.4]
  input  [63:0] io_argOuts_9_bits, // @[:@55603.4]
  input         io_argOuts_10_valid, // @[:@55603.4]
  input  [63:0] io_argOuts_10_bits, // @[:@55603.4]
  input         io_argOuts_11_valid, // @[:@55603.4]
  input  [63:0] io_argOuts_11_bits, // @[:@55603.4]
  input         io_argOuts_12_valid, // @[:@55603.4]
  input  [63:0] io_argOuts_12_bits, // @[:@55603.4]
  input         io_argOuts_13_valid, // @[:@55603.4]
  input  [63:0] io_argOuts_13_bits, // @[:@55603.4]
  input         io_argOuts_14_valid, // @[:@55603.4]
  input  [63:0] io_argOuts_14_bits, // @[:@55603.4]
  input         io_argOuts_15_valid, // @[:@55603.4]
  input  [63:0] io_argOuts_15_bits, // @[:@55603.4]
  input         io_argOuts_16_valid, // @[:@55603.4]
  input  [63:0] io_argOuts_16_bits, // @[:@55603.4]
  input         io_argOuts_17_valid, // @[:@55603.4]
  input  [63:0] io_argOuts_17_bits, // @[:@55603.4]
  input         io_argOuts_18_valid, // @[:@55603.4]
  input  [63:0] io_argOuts_18_bits, // @[:@55603.4]
  input         io_argOuts_19_valid, // @[:@55603.4]
  input  [63:0] io_argOuts_19_bits, // @[:@55603.4]
  input         io_argOuts_20_valid, // @[:@55603.4]
  input  [63:0] io_argOuts_20_bits, // @[:@55603.4]
  input         io_argOuts_21_valid, // @[:@55603.4]
  input  [63:0] io_argOuts_21_bits, // @[:@55603.4]
  input         io_argOuts_22_valid, // @[:@55603.4]
  input  [63:0] io_argOuts_22_bits, // @[:@55603.4]
  input         io_argOuts_23_valid, // @[:@55603.4]
  input  [63:0] io_argOuts_23_bits, // @[:@55603.4]
  input         io_argOuts_24_valid, // @[:@55603.4]
  input  [63:0] io_argOuts_24_bits, // @[:@55603.4]
  input         io_argOuts_25_valid, // @[:@55603.4]
  input  [63:0] io_argOuts_25_bits, // @[:@55603.4]
  input         io_argOuts_26_valid, // @[:@55603.4]
  input  [63:0] io_argOuts_26_bits, // @[:@55603.4]
  input         io_argOuts_27_valid, // @[:@55603.4]
  input  [63:0] io_argOuts_27_bits, // @[:@55603.4]
  input         io_argOuts_28_valid, // @[:@55603.4]
  input  [63:0] io_argOuts_28_bits, // @[:@55603.4]
  input         io_argOuts_29_valid, // @[:@55603.4]
  input  [63:0] io_argOuts_29_bits, // @[:@55603.4]
  input         io_argOuts_30_valid, // @[:@55603.4]
  input  [63:0] io_argOuts_30_bits, // @[:@55603.4]
  input         io_argOuts_31_valid, // @[:@55603.4]
  input  [63:0] io_argOuts_31_bits, // @[:@55603.4]
  input         io_heap_0_req_valid, // @[:@55603.4]
  input         io_heap_0_req_bits_allocDealloc, // @[:@55603.4]
  input  [63:0] io_heap_0_req_bits_sizeAddr, // @[:@55603.4]
  output        io_heap_0_resp_valid, // @[:@55603.4]
  output        io_heap_0_resp_bits_allocDealloc, // @[:@55603.4]
  output [63:0] io_heap_0_resp_bits_sizeAddr // @[:@55603.4]
);
  wire  fringeCommon_clock; // @[FringeZynq.scala 68:28:@56089.4]
  wire  fringeCommon_reset; // @[FringeZynq.scala 68:28:@56089.4]
  wire [31:0] fringeCommon_io_raddr; // @[FringeZynq.scala 68:28:@56089.4]
  wire  fringeCommon_io_wen; // @[FringeZynq.scala 68:28:@56089.4]
  wire [31:0] fringeCommon_io_waddr; // @[FringeZynq.scala 68:28:@56089.4]
  wire [63:0] fringeCommon_io_wdata; // @[FringeZynq.scala 68:28:@56089.4]
  wire [63:0] fringeCommon_io_rdata; // @[FringeZynq.scala 68:28:@56089.4]
  wire  fringeCommon_io_enable; // @[FringeZynq.scala 68:28:@56089.4]
  wire  fringeCommon_io_done; // @[FringeZynq.scala 68:28:@56089.4]
  wire  fringeCommon_io_reset; // @[FringeZynq.scala 68:28:@56089.4]
  wire [63:0] fringeCommon_io_argIns_0; // @[FringeZynq.scala 68:28:@56089.4]
  wire  fringeCommon_io_argOuts_0_valid; // @[FringeZynq.scala 68:28:@56089.4]
  wire [63:0] fringeCommon_io_argOuts_0_bits; // @[FringeZynq.scala 68:28:@56089.4]
  wire  fringeCommon_io_argOuts_1_valid; // @[FringeZynq.scala 68:28:@56089.4]
  wire [63:0] fringeCommon_io_argOuts_1_bits; // @[FringeZynq.scala 68:28:@56089.4]
  wire  fringeCommon_io_argOuts_2_valid; // @[FringeZynq.scala 68:28:@56089.4]
  wire [63:0] fringeCommon_io_argOuts_2_bits; // @[FringeZynq.scala 68:28:@56089.4]
  wire  fringeCommon_io_argOuts_3_valid; // @[FringeZynq.scala 68:28:@56089.4]
  wire [63:0] fringeCommon_io_argOuts_3_bits; // @[FringeZynq.scala 68:28:@56089.4]
  wire  fringeCommon_io_argOuts_4_valid; // @[FringeZynq.scala 68:28:@56089.4]
  wire [63:0] fringeCommon_io_argOuts_4_bits; // @[FringeZynq.scala 68:28:@56089.4]
  wire  fringeCommon_io_argOuts_5_valid; // @[FringeZynq.scala 68:28:@56089.4]
  wire [63:0] fringeCommon_io_argOuts_5_bits; // @[FringeZynq.scala 68:28:@56089.4]
  wire  fringeCommon_io_argOuts_6_valid; // @[FringeZynq.scala 68:28:@56089.4]
  wire [63:0] fringeCommon_io_argOuts_6_bits; // @[FringeZynq.scala 68:28:@56089.4]
  wire  fringeCommon_io_argOuts_7_valid; // @[FringeZynq.scala 68:28:@56089.4]
  wire [63:0] fringeCommon_io_argOuts_7_bits; // @[FringeZynq.scala 68:28:@56089.4]
  wire  fringeCommon_io_argOuts_8_valid; // @[FringeZynq.scala 68:28:@56089.4]
  wire [63:0] fringeCommon_io_argOuts_8_bits; // @[FringeZynq.scala 68:28:@56089.4]
  wire  fringeCommon_io_argOuts_9_valid; // @[FringeZynq.scala 68:28:@56089.4]
  wire [63:0] fringeCommon_io_argOuts_9_bits; // @[FringeZynq.scala 68:28:@56089.4]
  wire  fringeCommon_io_argOuts_10_valid; // @[FringeZynq.scala 68:28:@56089.4]
  wire [63:0] fringeCommon_io_argOuts_10_bits; // @[FringeZynq.scala 68:28:@56089.4]
  wire  fringeCommon_io_argOuts_11_valid; // @[FringeZynq.scala 68:28:@56089.4]
  wire [63:0] fringeCommon_io_argOuts_11_bits; // @[FringeZynq.scala 68:28:@56089.4]
  wire  fringeCommon_io_argOuts_12_valid; // @[FringeZynq.scala 68:28:@56089.4]
  wire [63:0] fringeCommon_io_argOuts_12_bits; // @[FringeZynq.scala 68:28:@56089.4]
  wire  fringeCommon_io_argOuts_13_valid; // @[FringeZynq.scala 68:28:@56089.4]
  wire [63:0] fringeCommon_io_argOuts_13_bits; // @[FringeZynq.scala 68:28:@56089.4]
  wire  fringeCommon_io_argOuts_14_valid; // @[FringeZynq.scala 68:28:@56089.4]
  wire [63:0] fringeCommon_io_argOuts_14_bits; // @[FringeZynq.scala 68:28:@56089.4]
  wire  fringeCommon_io_argOuts_15_valid; // @[FringeZynq.scala 68:28:@56089.4]
  wire [63:0] fringeCommon_io_argOuts_15_bits; // @[FringeZynq.scala 68:28:@56089.4]
  wire  fringeCommon_io_argOuts_16_valid; // @[FringeZynq.scala 68:28:@56089.4]
  wire [63:0] fringeCommon_io_argOuts_16_bits; // @[FringeZynq.scala 68:28:@56089.4]
  wire  fringeCommon_io_argOuts_17_valid; // @[FringeZynq.scala 68:28:@56089.4]
  wire [63:0] fringeCommon_io_argOuts_17_bits; // @[FringeZynq.scala 68:28:@56089.4]
  wire  fringeCommon_io_argOuts_18_valid; // @[FringeZynq.scala 68:28:@56089.4]
  wire [63:0] fringeCommon_io_argOuts_18_bits; // @[FringeZynq.scala 68:28:@56089.4]
  wire  fringeCommon_io_argOuts_19_valid; // @[FringeZynq.scala 68:28:@56089.4]
  wire [63:0] fringeCommon_io_argOuts_19_bits; // @[FringeZynq.scala 68:28:@56089.4]
  wire  fringeCommon_io_argOuts_20_valid; // @[FringeZynq.scala 68:28:@56089.4]
  wire [63:0] fringeCommon_io_argOuts_20_bits; // @[FringeZynq.scala 68:28:@56089.4]
  wire  fringeCommon_io_argOuts_21_valid; // @[FringeZynq.scala 68:28:@56089.4]
  wire [63:0] fringeCommon_io_argOuts_21_bits; // @[FringeZynq.scala 68:28:@56089.4]
  wire  fringeCommon_io_argOuts_22_valid; // @[FringeZynq.scala 68:28:@56089.4]
  wire [63:0] fringeCommon_io_argOuts_22_bits; // @[FringeZynq.scala 68:28:@56089.4]
  wire  fringeCommon_io_argOuts_23_valid; // @[FringeZynq.scala 68:28:@56089.4]
  wire [63:0] fringeCommon_io_argOuts_23_bits; // @[FringeZynq.scala 68:28:@56089.4]
  wire  fringeCommon_io_argOuts_24_valid; // @[FringeZynq.scala 68:28:@56089.4]
  wire [63:0] fringeCommon_io_argOuts_24_bits; // @[FringeZynq.scala 68:28:@56089.4]
  wire  fringeCommon_io_argOuts_25_valid; // @[FringeZynq.scala 68:28:@56089.4]
  wire [63:0] fringeCommon_io_argOuts_25_bits; // @[FringeZynq.scala 68:28:@56089.4]
  wire  fringeCommon_io_argOuts_26_valid; // @[FringeZynq.scala 68:28:@56089.4]
  wire [63:0] fringeCommon_io_argOuts_26_bits; // @[FringeZynq.scala 68:28:@56089.4]
  wire  fringeCommon_io_argOuts_27_valid; // @[FringeZynq.scala 68:28:@56089.4]
  wire [63:0] fringeCommon_io_argOuts_27_bits; // @[FringeZynq.scala 68:28:@56089.4]
  wire  fringeCommon_io_argOuts_28_valid; // @[FringeZynq.scala 68:28:@56089.4]
  wire [63:0] fringeCommon_io_argOuts_28_bits; // @[FringeZynq.scala 68:28:@56089.4]
  wire  fringeCommon_io_argOuts_29_valid; // @[FringeZynq.scala 68:28:@56089.4]
  wire [63:0] fringeCommon_io_argOuts_29_bits; // @[FringeZynq.scala 68:28:@56089.4]
  wire  fringeCommon_io_argOuts_30_valid; // @[FringeZynq.scala 68:28:@56089.4]
  wire [63:0] fringeCommon_io_argOuts_30_bits; // @[FringeZynq.scala 68:28:@56089.4]
  wire  fringeCommon_io_argOuts_31_valid; // @[FringeZynq.scala 68:28:@56089.4]
  wire [63:0] fringeCommon_io_argOuts_31_bits; // @[FringeZynq.scala 68:28:@56089.4]
  wire  fringeCommon_io_heap_0_req_valid; // @[FringeZynq.scala 68:28:@56089.4]
  wire  fringeCommon_io_heap_0_req_bits_allocDealloc; // @[FringeZynq.scala 68:28:@56089.4]
  wire [63:0] fringeCommon_io_heap_0_req_bits_sizeAddr; // @[FringeZynq.scala 68:28:@56089.4]
  wire  fringeCommon_io_heap_0_resp_valid; // @[FringeZynq.scala 68:28:@56089.4]
  wire  fringeCommon_io_heap_0_resp_bits_allocDealloc; // @[FringeZynq.scala 68:28:@56089.4]
  wire [63:0] fringeCommon_io_heap_0_resp_bits_sizeAddr; // @[FringeZynq.scala 68:28:@56089.4]
  wire  AXI4LiteToRFBridgeKCU1500_clock; // @[FringeZynq.scala 78:31:@56797.4]
  wire  AXI4LiteToRFBridgeKCU1500_reset; // @[FringeZynq.scala 78:31:@56797.4]
  wire [31:0] AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWADDR; // @[FringeZynq.scala 78:31:@56797.4]
  wire [2:0] AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWPROT; // @[FringeZynq.scala 78:31:@56797.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWVALID; // @[FringeZynq.scala 78:31:@56797.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWREADY; // @[FringeZynq.scala 78:31:@56797.4]
  wire [31:0] AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARADDR; // @[FringeZynq.scala 78:31:@56797.4]
  wire [2:0] AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARPROT; // @[FringeZynq.scala 78:31:@56797.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARVALID; // @[FringeZynq.scala 78:31:@56797.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARREADY; // @[FringeZynq.scala 78:31:@56797.4]
  wire [31:0] AXI4LiteToRFBridgeKCU1500_io_S_AXI_WDATA; // @[FringeZynq.scala 78:31:@56797.4]
  wire [3:0] AXI4LiteToRFBridgeKCU1500_io_S_AXI_WSTRB; // @[FringeZynq.scala 78:31:@56797.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_WVALID; // @[FringeZynq.scala 78:31:@56797.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_WREADY; // @[FringeZynq.scala 78:31:@56797.4]
  wire [31:0] AXI4LiteToRFBridgeKCU1500_io_S_AXI_RDATA; // @[FringeZynq.scala 78:31:@56797.4]
  wire [1:0] AXI4LiteToRFBridgeKCU1500_io_S_AXI_RRESP; // @[FringeZynq.scala 78:31:@56797.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_RVALID; // @[FringeZynq.scala 78:31:@56797.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_RREADY; // @[FringeZynq.scala 78:31:@56797.4]
  wire [1:0] AXI4LiteToRFBridgeKCU1500_io_S_AXI_BRESP; // @[FringeZynq.scala 78:31:@56797.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_BVALID; // @[FringeZynq.scala 78:31:@56797.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_BREADY; // @[FringeZynq.scala 78:31:@56797.4]
  wire [31:0] AXI4LiteToRFBridgeKCU1500_io_raddr; // @[FringeZynq.scala 78:31:@56797.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_wen; // @[FringeZynq.scala 78:31:@56797.4]
  wire [31:0] AXI4LiteToRFBridgeKCU1500_io_waddr; // @[FringeZynq.scala 78:31:@56797.4]
  wire [31:0] AXI4LiteToRFBridgeKCU1500_io_wdata; // @[FringeZynq.scala 78:31:@56797.4]
  wire [31:0] AXI4LiteToRFBridgeKCU1500_io_rdata; // @[FringeZynq.scala 78:31:@56797.4]
  wire [7:0] MAGToAXI4Bridge_io_M_AXI_AWLEN; // @[FringeZynq.scala 130:27:@57056.4]
  wire [7:0] MAGToAXI4Bridge_io_M_AXI_ARLEN; // @[FringeZynq.scala 130:27:@57056.4]
  Fringe fringeCommon ( // @[FringeZynq.scala 68:28:@56089.4]
    .clock(fringeCommon_clock),
    .reset(fringeCommon_reset),
    .io_raddr(fringeCommon_io_raddr),
    .io_wen(fringeCommon_io_wen),
    .io_waddr(fringeCommon_io_waddr),
    .io_wdata(fringeCommon_io_wdata),
    .io_rdata(fringeCommon_io_rdata),
    .io_enable(fringeCommon_io_enable),
    .io_done(fringeCommon_io_done),
    .io_reset(fringeCommon_io_reset),
    .io_argIns_0(fringeCommon_io_argIns_0),
    .io_argOuts_0_valid(fringeCommon_io_argOuts_0_valid),
    .io_argOuts_0_bits(fringeCommon_io_argOuts_0_bits),
    .io_argOuts_1_valid(fringeCommon_io_argOuts_1_valid),
    .io_argOuts_1_bits(fringeCommon_io_argOuts_1_bits),
    .io_argOuts_2_valid(fringeCommon_io_argOuts_2_valid),
    .io_argOuts_2_bits(fringeCommon_io_argOuts_2_bits),
    .io_argOuts_3_valid(fringeCommon_io_argOuts_3_valid),
    .io_argOuts_3_bits(fringeCommon_io_argOuts_3_bits),
    .io_argOuts_4_valid(fringeCommon_io_argOuts_4_valid),
    .io_argOuts_4_bits(fringeCommon_io_argOuts_4_bits),
    .io_argOuts_5_valid(fringeCommon_io_argOuts_5_valid),
    .io_argOuts_5_bits(fringeCommon_io_argOuts_5_bits),
    .io_argOuts_6_valid(fringeCommon_io_argOuts_6_valid),
    .io_argOuts_6_bits(fringeCommon_io_argOuts_6_bits),
    .io_argOuts_7_valid(fringeCommon_io_argOuts_7_valid),
    .io_argOuts_7_bits(fringeCommon_io_argOuts_7_bits),
    .io_argOuts_8_valid(fringeCommon_io_argOuts_8_valid),
    .io_argOuts_8_bits(fringeCommon_io_argOuts_8_bits),
    .io_argOuts_9_valid(fringeCommon_io_argOuts_9_valid),
    .io_argOuts_9_bits(fringeCommon_io_argOuts_9_bits),
    .io_argOuts_10_valid(fringeCommon_io_argOuts_10_valid),
    .io_argOuts_10_bits(fringeCommon_io_argOuts_10_bits),
    .io_argOuts_11_valid(fringeCommon_io_argOuts_11_valid),
    .io_argOuts_11_bits(fringeCommon_io_argOuts_11_bits),
    .io_argOuts_12_valid(fringeCommon_io_argOuts_12_valid),
    .io_argOuts_12_bits(fringeCommon_io_argOuts_12_bits),
    .io_argOuts_13_valid(fringeCommon_io_argOuts_13_valid),
    .io_argOuts_13_bits(fringeCommon_io_argOuts_13_bits),
    .io_argOuts_14_valid(fringeCommon_io_argOuts_14_valid),
    .io_argOuts_14_bits(fringeCommon_io_argOuts_14_bits),
    .io_argOuts_15_valid(fringeCommon_io_argOuts_15_valid),
    .io_argOuts_15_bits(fringeCommon_io_argOuts_15_bits),
    .io_argOuts_16_valid(fringeCommon_io_argOuts_16_valid),
    .io_argOuts_16_bits(fringeCommon_io_argOuts_16_bits),
    .io_argOuts_17_valid(fringeCommon_io_argOuts_17_valid),
    .io_argOuts_17_bits(fringeCommon_io_argOuts_17_bits),
    .io_argOuts_18_valid(fringeCommon_io_argOuts_18_valid),
    .io_argOuts_18_bits(fringeCommon_io_argOuts_18_bits),
    .io_argOuts_19_valid(fringeCommon_io_argOuts_19_valid),
    .io_argOuts_19_bits(fringeCommon_io_argOuts_19_bits),
    .io_argOuts_20_valid(fringeCommon_io_argOuts_20_valid),
    .io_argOuts_20_bits(fringeCommon_io_argOuts_20_bits),
    .io_argOuts_21_valid(fringeCommon_io_argOuts_21_valid),
    .io_argOuts_21_bits(fringeCommon_io_argOuts_21_bits),
    .io_argOuts_22_valid(fringeCommon_io_argOuts_22_valid),
    .io_argOuts_22_bits(fringeCommon_io_argOuts_22_bits),
    .io_argOuts_23_valid(fringeCommon_io_argOuts_23_valid),
    .io_argOuts_23_bits(fringeCommon_io_argOuts_23_bits),
    .io_argOuts_24_valid(fringeCommon_io_argOuts_24_valid),
    .io_argOuts_24_bits(fringeCommon_io_argOuts_24_bits),
    .io_argOuts_25_valid(fringeCommon_io_argOuts_25_valid),
    .io_argOuts_25_bits(fringeCommon_io_argOuts_25_bits),
    .io_argOuts_26_valid(fringeCommon_io_argOuts_26_valid),
    .io_argOuts_26_bits(fringeCommon_io_argOuts_26_bits),
    .io_argOuts_27_valid(fringeCommon_io_argOuts_27_valid),
    .io_argOuts_27_bits(fringeCommon_io_argOuts_27_bits),
    .io_argOuts_28_valid(fringeCommon_io_argOuts_28_valid),
    .io_argOuts_28_bits(fringeCommon_io_argOuts_28_bits),
    .io_argOuts_29_valid(fringeCommon_io_argOuts_29_valid),
    .io_argOuts_29_bits(fringeCommon_io_argOuts_29_bits),
    .io_argOuts_30_valid(fringeCommon_io_argOuts_30_valid),
    .io_argOuts_30_bits(fringeCommon_io_argOuts_30_bits),
    .io_argOuts_31_valid(fringeCommon_io_argOuts_31_valid),
    .io_argOuts_31_bits(fringeCommon_io_argOuts_31_bits),
    .io_heap_0_req_valid(fringeCommon_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(fringeCommon_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(fringeCommon_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(fringeCommon_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(fringeCommon_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(fringeCommon_io_heap_0_resp_bits_sizeAddr)
  );
  AXI4LiteToRFBridgeKCU1500 AXI4LiteToRFBridgeKCU1500 ( // @[FringeZynq.scala 78:31:@56797.4]
    .clock(AXI4LiteToRFBridgeKCU1500_clock),
    .reset(AXI4LiteToRFBridgeKCU1500_reset),
    .io_S_AXI_AWADDR(AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWADDR),
    .io_S_AXI_AWPROT(AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWPROT),
    .io_S_AXI_AWVALID(AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWVALID),
    .io_S_AXI_AWREADY(AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWREADY),
    .io_S_AXI_ARADDR(AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARADDR),
    .io_S_AXI_ARPROT(AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARPROT),
    .io_S_AXI_ARVALID(AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARVALID),
    .io_S_AXI_ARREADY(AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARREADY),
    .io_S_AXI_WDATA(AXI4LiteToRFBridgeKCU1500_io_S_AXI_WDATA),
    .io_S_AXI_WSTRB(AXI4LiteToRFBridgeKCU1500_io_S_AXI_WSTRB),
    .io_S_AXI_WVALID(AXI4LiteToRFBridgeKCU1500_io_S_AXI_WVALID),
    .io_S_AXI_WREADY(AXI4LiteToRFBridgeKCU1500_io_S_AXI_WREADY),
    .io_S_AXI_RDATA(AXI4LiteToRFBridgeKCU1500_io_S_AXI_RDATA),
    .io_S_AXI_RRESP(AXI4LiteToRFBridgeKCU1500_io_S_AXI_RRESP),
    .io_S_AXI_RVALID(AXI4LiteToRFBridgeKCU1500_io_S_AXI_RVALID),
    .io_S_AXI_RREADY(AXI4LiteToRFBridgeKCU1500_io_S_AXI_RREADY),
    .io_S_AXI_BRESP(AXI4LiteToRFBridgeKCU1500_io_S_AXI_BRESP),
    .io_S_AXI_BVALID(AXI4LiteToRFBridgeKCU1500_io_S_AXI_BVALID),
    .io_S_AXI_BREADY(AXI4LiteToRFBridgeKCU1500_io_S_AXI_BREADY),
    .io_raddr(AXI4LiteToRFBridgeKCU1500_io_raddr),
    .io_wen(AXI4LiteToRFBridgeKCU1500_io_wen),
    .io_waddr(AXI4LiteToRFBridgeKCU1500_io_waddr),
    .io_wdata(AXI4LiteToRFBridgeKCU1500_io_wdata),
    .io_rdata(AXI4LiteToRFBridgeKCU1500_io_rdata)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge ( // @[FringeZynq.scala 130:27:@57056.4]
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_io_M_AXI_AWLEN),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_io_M_AXI_ARLEN)
  );
  assign io_S_AXI_AWREADY = AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWREADY; // @[FringeZynq.scala 79:28:@56815.4]
  assign io_S_AXI_ARREADY = AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARREADY; // @[FringeZynq.scala 79:28:@56811.4]
  assign io_S_AXI_WREADY = AXI4LiteToRFBridgeKCU1500_io_S_AXI_WREADY; // @[FringeZynq.scala 79:28:@56807.4]
  assign io_S_AXI_RDATA = AXI4LiteToRFBridgeKCU1500_io_S_AXI_RDATA; // @[FringeZynq.scala 79:28:@56806.4]
  assign io_S_AXI_RRESP = AXI4LiteToRFBridgeKCU1500_io_S_AXI_RRESP; // @[FringeZynq.scala 79:28:@56805.4]
  assign io_S_AXI_RVALID = AXI4LiteToRFBridgeKCU1500_io_S_AXI_RVALID; // @[FringeZynq.scala 79:28:@56804.4]
  assign io_S_AXI_BRESP = AXI4LiteToRFBridgeKCU1500_io_S_AXI_BRESP; // @[FringeZynq.scala 79:28:@56802.4]
  assign io_S_AXI_BVALID = AXI4LiteToRFBridgeKCU1500_io_S_AXI_BVALID; // @[FringeZynq.scala 79:28:@56801.4]
  assign io_M_AXI_0_AWLEN = MAGToAXI4Bridge_io_M_AXI_AWLEN; // @[FringeZynq.scala 132:10:@57208.4]
  assign io_M_AXI_0_ARLEN = MAGToAXI4Bridge_io_M_AXI_ARLEN; // @[FringeZynq.scala 132:10:@57196.4]
  assign io_enable = fringeCommon_io_enable; // @[FringeZynq.scala 114:13:@56827.4]
  assign io_reset = fringeCommon_io_reset; // @[FringeZynq.scala 118:12:@56831.4]
  assign io_argIns_0 = fringeCommon_io_argIns_0; // @[FringeZynq.scala 120:13:@56832.4]
  assign io_heap_0_resp_valid = fringeCommon_io_heap_0_resp_valid; // @[FringeZynq.scala 126:11:@57052.4]
  assign io_heap_0_resp_bits_allocDealloc = fringeCommon_io_heap_0_resp_bits_allocDealloc; // @[FringeZynq.scala 126:11:@57051.4]
  assign io_heap_0_resp_bits_sizeAddr = fringeCommon_io_heap_0_resp_bits_sizeAddr; // @[FringeZynq.scala 126:11:@57050.4]
  assign fringeCommon_clock = clock; // @[:@56090.4]
  assign fringeCommon_reset = reset; // @[:@56091.4 FringeZynq.scala 81:24:@56820.4 FringeZynq.scala 116:22:@56830.4]
  assign fringeCommon_io_raddr = AXI4LiteToRFBridgeKCU1500_io_raddr; // @[FringeZynq.scala 82:27:@56821.4]
  assign fringeCommon_io_wen = AXI4LiteToRFBridgeKCU1500_io_wen; // @[FringeZynq.scala 83:27:@56822.4]
  assign fringeCommon_io_waddr = AXI4LiteToRFBridgeKCU1500_io_waddr; // @[FringeZynq.scala 84:27:@56823.4]
  assign fringeCommon_io_wdata = {{32'd0}, AXI4LiteToRFBridgeKCU1500_io_wdata}; // @[FringeZynq.scala 85:27:@56824.4]
  assign fringeCommon_io_done = io_done; // @[FringeZynq.scala 115:24:@56828.4]
  assign fringeCommon_io_argOuts_0_valid = io_argOuts_0_valid; // @[FringeZynq.scala 121:27:@56834.4]
  assign fringeCommon_io_argOuts_0_bits = io_argOuts_0_bits; // @[FringeZynq.scala 121:27:@56833.4]
  assign fringeCommon_io_argOuts_1_valid = io_argOuts_1_valid; // @[FringeZynq.scala 121:27:@56837.4]
  assign fringeCommon_io_argOuts_1_bits = io_argOuts_1_bits; // @[FringeZynq.scala 121:27:@56836.4]
  assign fringeCommon_io_argOuts_2_valid = io_argOuts_2_valid; // @[FringeZynq.scala 121:27:@56840.4]
  assign fringeCommon_io_argOuts_2_bits = io_argOuts_2_bits; // @[FringeZynq.scala 121:27:@56839.4]
  assign fringeCommon_io_argOuts_3_valid = io_argOuts_3_valid; // @[FringeZynq.scala 121:27:@56843.4]
  assign fringeCommon_io_argOuts_3_bits = io_argOuts_3_bits; // @[FringeZynq.scala 121:27:@56842.4]
  assign fringeCommon_io_argOuts_4_valid = io_argOuts_4_valid; // @[FringeZynq.scala 121:27:@56846.4]
  assign fringeCommon_io_argOuts_4_bits = io_argOuts_4_bits; // @[FringeZynq.scala 121:27:@56845.4]
  assign fringeCommon_io_argOuts_5_valid = io_argOuts_5_valid; // @[FringeZynq.scala 121:27:@56849.4]
  assign fringeCommon_io_argOuts_5_bits = io_argOuts_5_bits; // @[FringeZynq.scala 121:27:@56848.4]
  assign fringeCommon_io_argOuts_6_valid = io_argOuts_6_valid; // @[FringeZynq.scala 121:27:@56852.4]
  assign fringeCommon_io_argOuts_6_bits = io_argOuts_6_bits; // @[FringeZynq.scala 121:27:@56851.4]
  assign fringeCommon_io_argOuts_7_valid = io_argOuts_7_valid; // @[FringeZynq.scala 121:27:@56855.4]
  assign fringeCommon_io_argOuts_7_bits = io_argOuts_7_bits; // @[FringeZynq.scala 121:27:@56854.4]
  assign fringeCommon_io_argOuts_8_valid = io_argOuts_8_valid; // @[FringeZynq.scala 121:27:@56858.4]
  assign fringeCommon_io_argOuts_8_bits = io_argOuts_8_bits; // @[FringeZynq.scala 121:27:@56857.4]
  assign fringeCommon_io_argOuts_9_valid = io_argOuts_9_valid; // @[FringeZynq.scala 121:27:@56861.4]
  assign fringeCommon_io_argOuts_9_bits = io_argOuts_9_bits; // @[FringeZynq.scala 121:27:@56860.4]
  assign fringeCommon_io_argOuts_10_valid = io_argOuts_10_valid; // @[FringeZynq.scala 121:27:@56864.4]
  assign fringeCommon_io_argOuts_10_bits = io_argOuts_10_bits; // @[FringeZynq.scala 121:27:@56863.4]
  assign fringeCommon_io_argOuts_11_valid = io_argOuts_11_valid; // @[FringeZynq.scala 121:27:@56867.4]
  assign fringeCommon_io_argOuts_11_bits = io_argOuts_11_bits; // @[FringeZynq.scala 121:27:@56866.4]
  assign fringeCommon_io_argOuts_12_valid = io_argOuts_12_valid; // @[FringeZynq.scala 121:27:@56870.4]
  assign fringeCommon_io_argOuts_12_bits = io_argOuts_12_bits; // @[FringeZynq.scala 121:27:@56869.4]
  assign fringeCommon_io_argOuts_13_valid = io_argOuts_13_valid; // @[FringeZynq.scala 121:27:@56873.4]
  assign fringeCommon_io_argOuts_13_bits = io_argOuts_13_bits; // @[FringeZynq.scala 121:27:@56872.4]
  assign fringeCommon_io_argOuts_14_valid = io_argOuts_14_valid; // @[FringeZynq.scala 121:27:@56876.4]
  assign fringeCommon_io_argOuts_14_bits = io_argOuts_14_bits; // @[FringeZynq.scala 121:27:@56875.4]
  assign fringeCommon_io_argOuts_15_valid = io_argOuts_15_valid; // @[FringeZynq.scala 121:27:@56879.4]
  assign fringeCommon_io_argOuts_15_bits = io_argOuts_15_bits; // @[FringeZynq.scala 121:27:@56878.4]
  assign fringeCommon_io_argOuts_16_valid = io_argOuts_16_valid; // @[FringeZynq.scala 121:27:@56882.4]
  assign fringeCommon_io_argOuts_16_bits = io_argOuts_16_bits; // @[FringeZynq.scala 121:27:@56881.4]
  assign fringeCommon_io_argOuts_17_valid = io_argOuts_17_valid; // @[FringeZynq.scala 121:27:@56885.4]
  assign fringeCommon_io_argOuts_17_bits = io_argOuts_17_bits; // @[FringeZynq.scala 121:27:@56884.4]
  assign fringeCommon_io_argOuts_18_valid = io_argOuts_18_valid; // @[FringeZynq.scala 121:27:@56888.4]
  assign fringeCommon_io_argOuts_18_bits = io_argOuts_18_bits; // @[FringeZynq.scala 121:27:@56887.4]
  assign fringeCommon_io_argOuts_19_valid = io_argOuts_19_valid; // @[FringeZynq.scala 121:27:@56891.4]
  assign fringeCommon_io_argOuts_19_bits = io_argOuts_19_bits; // @[FringeZynq.scala 121:27:@56890.4]
  assign fringeCommon_io_argOuts_20_valid = io_argOuts_20_valid; // @[FringeZynq.scala 121:27:@56894.4]
  assign fringeCommon_io_argOuts_20_bits = io_argOuts_20_bits; // @[FringeZynq.scala 121:27:@56893.4]
  assign fringeCommon_io_argOuts_21_valid = io_argOuts_21_valid; // @[FringeZynq.scala 121:27:@56897.4]
  assign fringeCommon_io_argOuts_21_bits = io_argOuts_21_bits; // @[FringeZynq.scala 121:27:@56896.4]
  assign fringeCommon_io_argOuts_22_valid = io_argOuts_22_valid; // @[FringeZynq.scala 121:27:@56900.4]
  assign fringeCommon_io_argOuts_22_bits = io_argOuts_22_bits; // @[FringeZynq.scala 121:27:@56899.4]
  assign fringeCommon_io_argOuts_23_valid = io_argOuts_23_valid; // @[FringeZynq.scala 121:27:@56903.4]
  assign fringeCommon_io_argOuts_23_bits = io_argOuts_23_bits; // @[FringeZynq.scala 121:27:@56902.4]
  assign fringeCommon_io_argOuts_24_valid = io_argOuts_24_valid; // @[FringeZynq.scala 121:27:@56906.4]
  assign fringeCommon_io_argOuts_24_bits = io_argOuts_24_bits; // @[FringeZynq.scala 121:27:@56905.4]
  assign fringeCommon_io_argOuts_25_valid = io_argOuts_25_valid; // @[FringeZynq.scala 121:27:@56909.4]
  assign fringeCommon_io_argOuts_25_bits = io_argOuts_25_bits; // @[FringeZynq.scala 121:27:@56908.4]
  assign fringeCommon_io_argOuts_26_valid = io_argOuts_26_valid; // @[FringeZynq.scala 121:27:@56912.4]
  assign fringeCommon_io_argOuts_26_bits = io_argOuts_26_bits; // @[FringeZynq.scala 121:27:@56911.4]
  assign fringeCommon_io_argOuts_27_valid = io_argOuts_27_valid; // @[FringeZynq.scala 121:27:@56915.4]
  assign fringeCommon_io_argOuts_27_bits = io_argOuts_27_bits; // @[FringeZynq.scala 121:27:@56914.4]
  assign fringeCommon_io_argOuts_28_valid = io_argOuts_28_valid; // @[FringeZynq.scala 121:27:@56918.4]
  assign fringeCommon_io_argOuts_28_bits = io_argOuts_28_bits; // @[FringeZynq.scala 121:27:@56917.4]
  assign fringeCommon_io_argOuts_29_valid = io_argOuts_29_valid; // @[FringeZynq.scala 121:27:@56921.4]
  assign fringeCommon_io_argOuts_29_bits = io_argOuts_29_bits; // @[FringeZynq.scala 121:27:@56920.4]
  assign fringeCommon_io_argOuts_30_valid = io_argOuts_30_valid; // @[FringeZynq.scala 121:27:@56924.4]
  assign fringeCommon_io_argOuts_30_bits = io_argOuts_30_bits; // @[FringeZynq.scala 121:27:@56923.4]
  assign fringeCommon_io_argOuts_31_valid = io_argOuts_31_valid; // @[FringeZynq.scala 121:27:@56927.4]
  assign fringeCommon_io_argOuts_31_bits = io_argOuts_31_bits; // @[FringeZynq.scala 121:27:@56926.4]
  assign fringeCommon_io_heap_0_req_valid = io_heap_0_req_valid; // @[FringeZynq.scala 126:11:@57055.4]
  assign fringeCommon_io_heap_0_req_bits_allocDealloc = io_heap_0_req_bits_allocDealloc; // @[FringeZynq.scala 126:11:@57054.4]
  assign fringeCommon_io_heap_0_req_bits_sizeAddr = io_heap_0_req_bits_sizeAddr; // @[FringeZynq.scala 126:11:@57053.4]
  assign AXI4LiteToRFBridgeKCU1500_clock = clock; // @[:@56798.4]
  assign AXI4LiteToRFBridgeKCU1500_reset = reset; // @[:@56799.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[FringeZynq.scala 79:28:@56818.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[FringeZynq.scala 79:28:@56817.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[FringeZynq.scala 79:28:@56816.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[FringeZynq.scala 79:28:@56814.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[FringeZynq.scala 79:28:@56813.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[FringeZynq.scala 79:28:@56812.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_WDATA = io_S_AXI_WDATA; // @[FringeZynq.scala 79:28:@56810.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[FringeZynq.scala 79:28:@56809.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_WVALID = io_S_AXI_WVALID; // @[FringeZynq.scala 79:28:@56808.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_RREADY = io_S_AXI_RREADY; // @[FringeZynq.scala 79:28:@56803.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_BREADY = io_S_AXI_BREADY; // @[FringeZynq.scala 79:28:@56800.4]
  assign AXI4LiteToRFBridgeKCU1500_io_rdata = fringeCommon_io_rdata[31:0]; // @[FringeZynq.scala 86:28:@56825.4]
endmodule
module SpatialIP( // @[:@57213.2]
  input          clock, // @[:@57214.4]
  input          reset, // @[:@57215.4]
  input          io_raddr, // @[:@57216.4]
  input          io_wen, // @[:@57216.4]
  input          io_waddr, // @[:@57216.4]
  input          io_wdata, // @[:@57216.4]
  output         io_rdata, // @[:@57216.4]
  input  [31:0]  io_S_AXI_AWADDR, // @[:@57216.4]
  input  [2:0]   io_S_AXI_AWPROT, // @[:@57216.4]
  input          io_S_AXI_AWVALID, // @[:@57216.4]
  output         io_S_AXI_AWREADY, // @[:@57216.4]
  input  [31:0]  io_S_AXI_ARADDR, // @[:@57216.4]
  input  [2:0]   io_S_AXI_ARPROT, // @[:@57216.4]
  input          io_S_AXI_ARVALID, // @[:@57216.4]
  output         io_S_AXI_ARREADY, // @[:@57216.4]
  input  [31:0]  io_S_AXI_WDATA, // @[:@57216.4]
  input  [3:0]   io_S_AXI_WSTRB, // @[:@57216.4]
  input          io_S_AXI_WVALID, // @[:@57216.4]
  output         io_S_AXI_WREADY, // @[:@57216.4]
  output [31:0]  io_S_AXI_RDATA, // @[:@57216.4]
  output [1:0]   io_S_AXI_RRESP, // @[:@57216.4]
  output         io_S_AXI_RVALID, // @[:@57216.4]
  input          io_S_AXI_RREADY, // @[:@57216.4]
  output [1:0]   io_S_AXI_BRESP, // @[:@57216.4]
  output         io_S_AXI_BVALID, // @[:@57216.4]
  input          io_S_AXI_BREADY, // @[:@57216.4]
  output [3:0]   io_M_AXI_0_AWID, // @[:@57216.4]
  output [3:0]   io_M_AXI_0_AWUSER, // @[:@57216.4]
  output [31:0]  io_M_AXI_0_AWADDR, // @[:@57216.4]
  output [7:0]   io_M_AXI_0_AWLEN, // @[:@57216.4]
  output [2:0]   io_M_AXI_0_AWSIZE, // @[:@57216.4]
  output [1:0]   io_M_AXI_0_AWBURST, // @[:@57216.4]
  output         io_M_AXI_0_AWLOCK, // @[:@57216.4]
  output [3:0]   io_M_AXI_0_AWCACHE, // @[:@57216.4]
  output [2:0]   io_M_AXI_0_AWPROT, // @[:@57216.4]
  output [3:0]   io_M_AXI_0_AWQOS, // @[:@57216.4]
  output         io_M_AXI_0_AWVALID, // @[:@57216.4]
  input          io_M_AXI_0_AWREADY, // @[:@57216.4]
  output [3:0]   io_M_AXI_0_ARID, // @[:@57216.4]
  output [3:0]   io_M_AXI_0_ARUSER, // @[:@57216.4]
  output [31:0]  io_M_AXI_0_ARADDR, // @[:@57216.4]
  output [7:0]   io_M_AXI_0_ARLEN, // @[:@57216.4]
  output [2:0]   io_M_AXI_0_ARSIZE, // @[:@57216.4]
  output [1:0]   io_M_AXI_0_ARBURST, // @[:@57216.4]
  output         io_M_AXI_0_ARLOCK, // @[:@57216.4]
  output [3:0]   io_M_AXI_0_ARCACHE, // @[:@57216.4]
  output [2:0]   io_M_AXI_0_ARPROT, // @[:@57216.4]
  output [3:0]   io_M_AXI_0_ARQOS, // @[:@57216.4]
  output         io_M_AXI_0_ARVALID, // @[:@57216.4]
  input          io_M_AXI_0_ARREADY, // @[:@57216.4]
  output [511:0] io_M_AXI_0_WDATA, // @[:@57216.4]
  output [63:0]  io_M_AXI_0_WSTRB, // @[:@57216.4]
  output         io_M_AXI_0_WLAST, // @[:@57216.4]
  output         io_M_AXI_0_WVALID, // @[:@57216.4]
  input          io_M_AXI_0_WREADY, // @[:@57216.4]
  input  [3:0]   io_M_AXI_0_RID, // @[:@57216.4]
  input  [31:0]  io_M_AXI_0_RUSER, // @[:@57216.4]
  input  [511:0] io_M_AXI_0_RDATA, // @[:@57216.4]
  input  [1:0]   io_M_AXI_0_RRESP, // @[:@57216.4]
  input          io_M_AXI_0_RLAST, // @[:@57216.4]
  input          io_M_AXI_0_RVALID, // @[:@57216.4]
  output         io_M_AXI_0_RREADY, // @[:@57216.4]
  input  [3:0]   io_M_AXI_0_BID, // @[:@57216.4]
  input  [3:0]   io_M_AXI_0_BUSER, // @[:@57216.4]
  input  [1:0]   io_M_AXI_0_BRESP, // @[:@57216.4]
  input          io_M_AXI_0_BVALID, // @[:@57216.4]
  output         io_M_AXI_0_BREADY, // @[:@57216.4]
  input          io_AXIS_IN_TVALID, // @[:@57216.4]
  output         io_AXIS_IN_TREADY, // @[:@57216.4]
  input  [255:0] io_AXIS_IN_TDATA, // @[:@57216.4]
  input  [31:0]  io_AXIS_IN_TSTRB, // @[:@57216.4]
  input  [31:0]  io_AXIS_IN_TKEEP, // @[:@57216.4]
  input          io_AXIS_IN_TLAST, // @[:@57216.4]
  input  [3:0]   io_AXIS_IN_TID, // @[:@57216.4]
  input  [3:0]   io_AXIS_IN_TDEST, // @[:@57216.4]
  output         io_AXIS_OUT_TVALID, // @[:@57216.4]
  input          io_AXIS_OUT_TREADY, // @[:@57216.4]
  output [255:0] io_AXIS_OUT_TDATA, // @[:@57216.4]
  output [31:0]  io_AXIS_OUT_TSTRB, // @[:@57216.4]
  output [31:0]  io_AXIS_OUT_TKEEP, // @[:@57216.4]
  output         io_AXIS_OUT_TLAST, // @[:@57216.4]
  output [3:0]   io_AXIS_OUT_TID, // @[:@57216.4]
  output [3:0]   io_AXIS_OUT_TDEST // @[:@57216.4]
);
  wire  accel_clock; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_reset; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_enable; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_done; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_reset; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_memStreams_loads_0_cmd_ready; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_memStreams_loads_0_cmd_valid; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_memStreams_loads_0_cmd_bits_addr; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_loads_0_cmd_bits_size; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_memStreams_loads_0_data_ready; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_memStreams_loads_0_data_valid; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_0; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_1; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_2; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_3; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_4; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_5; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_6; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_7; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_8; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_9; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_10; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_11; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_12; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_13; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_14; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_15; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_memStreams_stores_0_cmd_ready; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_memStreams_stores_0_cmd_valid; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_memStreams_stores_0_cmd_bits_addr; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_stores_0_cmd_bits_size; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_memStreams_stores_0_data_ready; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_memStreams_stores_0_data_valid; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_0; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_1; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_2; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_3; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_4; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_5; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_6; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_7; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_8; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_9; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_10; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_11; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_12; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_13; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_14; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_15; // @[Instantiator.scala 85:44:@57218.4]
  wire [15:0] accel_io_memStreams_stores_0_data_bits_wstrb; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_memStreams_stores_0_wresp_ready; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_memStreams_stores_0_wresp_valid; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_memStreams_stores_0_wresp_bits; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_memStreams_gathers_0_cmd_ready; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_memStreams_gathers_0_cmd_valid; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_0; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_1; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_2; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_3; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_4; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_5; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_6; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_7; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_8; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_9; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_10; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_11; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_12; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_13; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_14; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_15; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_memStreams_gathers_0_data_ready; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_memStreams_gathers_0_data_valid; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_0; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_1; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_2; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_3; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_4; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_5; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_6; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_7; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_8; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_9; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_10; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_11; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_12; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_13; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_14; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_15; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_memStreams_scatters_0_cmd_ready; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_memStreams_scatters_0_cmd_valid; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_0; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_1; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_2; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_3; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_4; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_5; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_6; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_7; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_8; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_9; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_10; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_11; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_12; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_13; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_14; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_15; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_memStreams_scatters_0_wresp_ready; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_memStreams_scatters_0_wresp_valid; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_memStreams_scatters_0_wresp_bits; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_axiStreamsIn_0_TVALID; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_axiStreamsIn_0_TREADY; // @[Instantiator.scala 85:44:@57218.4]
  wire [255:0] accel_io_axiStreamsIn_0_TDATA; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_axiStreamsIn_0_TSTRB; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_axiStreamsIn_0_TKEEP; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_axiStreamsIn_0_TLAST; // @[Instantiator.scala 85:44:@57218.4]
  wire [7:0] accel_io_axiStreamsIn_0_TID; // @[Instantiator.scala 85:44:@57218.4]
  wire [7:0] accel_io_axiStreamsIn_0_TDEST; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_axiStreamsOut_0_TVALID; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_axiStreamsOut_0_TREADY; // @[Instantiator.scala 85:44:@57218.4]
  wire [255:0] accel_io_axiStreamsOut_0_TDATA; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_axiStreamsOut_0_TSTRB; // @[Instantiator.scala 85:44:@57218.4]
  wire [31:0] accel_io_axiStreamsOut_0_TKEEP; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_axiStreamsOut_0_TLAST; // @[Instantiator.scala 85:44:@57218.4]
  wire [7:0] accel_io_axiStreamsOut_0_TID; // @[Instantiator.scala 85:44:@57218.4]
  wire [7:0] accel_io_axiStreamsOut_0_TDEST; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_heap_0_req_valid; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_heap_0_req_bits_allocDealloc; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_heap_0_req_bits_sizeAddr; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_heap_0_resp_valid; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_heap_0_resp_bits_allocDealloc; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_heap_0_resp_bits_sizeAddr; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argIns_0; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_0_port_ready; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_0_port_valid; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_0_port_bits; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_0_echo; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_1_port_ready; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_1_port_valid; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_1_port_bits; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_1_echo; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_2_port_ready; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_2_port_valid; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_2_port_bits; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_2_echo; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_3_port_ready; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_3_port_valid; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_3_port_bits; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_3_echo; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_4_port_ready; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_4_port_valid; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_4_port_bits; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_4_echo; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_5_port_ready; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_5_port_valid; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_5_port_bits; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_5_echo; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_6_port_ready; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_6_port_valid; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_6_port_bits; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_6_echo; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_7_port_ready; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_7_port_valid; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_7_port_bits; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_7_echo; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_8_port_ready; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_8_port_valid; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_8_port_bits; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_8_echo; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_9_port_ready; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_9_port_valid; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_9_port_bits; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_9_echo; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_10_port_ready; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_10_port_valid; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_10_port_bits; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_10_echo; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_11_port_ready; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_11_port_valid; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_11_port_bits; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_11_echo; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_12_port_ready; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_12_port_valid; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_12_port_bits; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_12_echo; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_13_port_ready; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_13_port_valid; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_13_port_bits; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_13_echo; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_14_port_ready; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_14_port_valid; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_14_port_bits; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_14_echo; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_15_port_ready; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_15_port_valid; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_15_port_bits; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_15_echo; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_16_port_ready; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_16_port_valid; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_16_port_bits; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_16_echo; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_17_port_ready; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_17_port_valid; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_17_port_bits; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_17_echo; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_18_port_ready; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_18_port_valid; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_18_port_bits; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_18_echo; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_19_port_ready; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_19_port_valid; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_19_port_bits; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_19_echo; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_20_port_ready; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_20_port_valid; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_20_port_bits; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_20_echo; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_21_port_ready; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_21_port_valid; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_21_port_bits; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_21_echo; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_22_port_ready; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_22_port_valid; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_22_port_bits; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_22_echo; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_23_port_ready; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_23_port_valid; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_23_port_bits; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_23_echo; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_24_port_ready; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_24_port_valid; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_24_port_bits; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_24_echo; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_25_port_ready; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_25_port_valid; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_25_port_bits; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_25_echo; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_26_port_ready; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_26_port_valid; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_26_port_bits; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_26_echo; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_27_port_ready; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_27_port_valid; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_27_port_bits; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_27_echo; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_28_port_ready; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_28_port_valid; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_28_port_bits; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_28_echo; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_29_port_ready; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_29_port_valid; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_29_port_bits; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_29_echo; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_30_port_ready; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_30_port_valid; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_30_port_bits; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_30_echo; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_31_port_ready; // @[Instantiator.scala 85:44:@57218.4]
  wire  accel_io_argOuts_31_port_valid; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_31_port_bits; // @[Instantiator.scala 85:44:@57218.4]
  wire [63:0] accel_io_argOuts_31_echo; // @[Instantiator.scala 85:44:@57218.4]
  wire  FringeZynq_clock; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_reset; // @[KCU1500.scala 21:24:@57496.4]
  wire [31:0] FringeZynq_io_S_AXI_AWADDR; // @[KCU1500.scala 21:24:@57496.4]
  wire [2:0] FringeZynq_io_S_AXI_AWPROT; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_S_AXI_AWVALID; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_S_AXI_AWREADY; // @[KCU1500.scala 21:24:@57496.4]
  wire [31:0] FringeZynq_io_S_AXI_ARADDR; // @[KCU1500.scala 21:24:@57496.4]
  wire [2:0] FringeZynq_io_S_AXI_ARPROT; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_S_AXI_ARVALID; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_S_AXI_ARREADY; // @[KCU1500.scala 21:24:@57496.4]
  wire [31:0] FringeZynq_io_S_AXI_WDATA; // @[KCU1500.scala 21:24:@57496.4]
  wire [3:0] FringeZynq_io_S_AXI_WSTRB; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_S_AXI_WVALID; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_S_AXI_WREADY; // @[KCU1500.scala 21:24:@57496.4]
  wire [31:0] FringeZynq_io_S_AXI_RDATA; // @[KCU1500.scala 21:24:@57496.4]
  wire [1:0] FringeZynq_io_S_AXI_RRESP; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_S_AXI_RVALID; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_S_AXI_RREADY; // @[KCU1500.scala 21:24:@57496.4]
  wire [1:0] FringeZynq_io_S_AXI_BRESP; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_S_AXI_BVALID; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_S_AXI_BREADY; // @[KCU1500.scala 21:24:@57496.4]
  wire [7:0] FringeZynq_io_M_AXI_0_AWLEN; // @[KCU1500.scala 21:24:@57496.4]
  wire [7:0] FringeZynq_io_M_AXI_0_ARLEN; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_enable; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_done; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_reset; // @[KCU1500.scala 21:24:@57496.4]
  wire [63:0] FringeZynq_io_argIns_0; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_argOuts_0_valid; // @[KCU1500.scala 21:24:@57496.4]
  wire [63:0] FringeZynq_io_argOuts_0_bits; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_argOuts_1_valid; // @[KCU1500.scala 21:24:@57496.4]
  wire [63:0] FringeZynq_io_argOuts_1_bits; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_argOuts_2_valid; // @[KCU1500.scala 21:24:@57496.4]
  wire [63:0] FringeZynq_io_argOuts_2_bits; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_argOuts_3_valid; // @[KCU1500.scala 21:24:@57496.4]
  wire [63:0] FringeZynq_io_argOuts_3_bits; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_argOuts_4_valid; // @[KCU1500.scala 21:24:@57496.4]
  wire [63:0] FringeZynq_io_argOuts_4_bits; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_argOuts_5_valid; // @[KCU1500.scala 21:24:@57496.4]
  wire [63:0] FringeZynq_io_argOuts_5_bits; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_argOuts_6_valid; // @[KCU1500.scala 21:24:@57496.4]
  wire [63:0] FringeZynq_io_argOuts_6_bits; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_argOuts_7_valid; // @[KCU1500.scala 21:24:@57496.4]
  wire [63:0] FringeZynq_io_argOuts_7_bits; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_argOuts_8_valid; // @[KCU1500.scala 21:24:@57496.4]
  wire [63:0] FringeZynq_io_argOuts_8_bits; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_argOuts_9_valid; // @[KCU1500.scala 21:24:@57496.4]
  wire [63:0] FringeZynq_io_argOuts_9_bits; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_argOuts_10_valid; // @[KCU1500.scala 21:24:@57496.4]
  wire [63:0] FringeZynq_io_argOuts_10_bits; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_argOuts_11_valid; // @[KCU1500.scala 21:24:@57496.4]
  wire [63:0] FringeZynq_io_argOuts_11_bits; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_argOuts_12_valid; // @[KCU1500.scala 21:24:@57496.4]
  wire [63:0] FringeZynq_io_argOuts_12_bits; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_argOuts_13_valid; // @[KCU1500.scala 21:24:@57496.4]
  wire [63:0] FringeZynq_io_argOuts_13_bits; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_argOuts_14_valid; // @[KCU1500.scala 21:24:@57496.4]
  wire [63:0] FringeZynq_io_argOuts_14_bits; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_argOuts_15_valid; // @[KCU1500.scala 21:24:@57496.4]
  wire [63:0] FringeZynq_io_argOuts_15_bits; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_argOuts_16_valid; // @[KCU1500.scala 21:24:@57496.4]
  wire [63:0] FringeZynq_io_argOuts_16_bits; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_argOuts_17_valid; // @[KCU1500.scala 21:24:@57496.4]
  wire [63:0] FringeZynq_io_argOuts_17_bits; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_argOuts_18_valid; // @[KCU1500.scala 21:24:@57496.4]
  wire [63:0] FringeZynq_io_argOuts_18_bits; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_argOuts_19_valid; // @[KCU1500.scala 21:24:@57496.4]
  wire [63:0] FringeZynq_io_argOuts_19_bits; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_argOuts_20_valid; // @[KCU1500.scala 21:24:@57496.4]
  wire [63:0] FringeZynq_io_argOuts_20_bits; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_argOuts_21_valid; // @[KCU1500.scala 21:24:@57496.4]
  wire [63:0] FringeZynq_io_argOuts_21_bits; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_argOuts_22_valid; // @[KCU1500.scala 21:24:@57496.4]
  wire [63:0] FringeZynq_io_argOuts_22_bits; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_argOuts_23_valid; // @[KCU1500.scala 21:24:@57496.4]
  wire [63:0] FringeZynq_io_argOuts_23_bits; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_argOuts_24_valid; // @[KCU1500.scala 21:24:@57496.4]
  wire [63:0] FringeZynq_io_argOuts_24_bits; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_argOuts_25_valid; // @[KCU1500.scala 21:24:@57496.4]
  wire [63:0] FringeZynq_io_argOuts_25_bits; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_argOuts_26_valid; // @[KCU1500.scala 21:24:@57496.4]
  wire [63:0] FringeZynq_io_argOuts_26_bits; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_argOuts_27_valid; // @[KCU1500.scala 21:24:@57496.4]
  wire [63:0] FringeZynq_io_argOuts_27_bits; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_argOuts_28_valid; // @[KCU1500.scala 21:24:@57496.4]
  wire [63:0] FringeZynq_io_argOuts_28_bits; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_argOuts_29_valid; // @[KCU1500.scala 21:24:@57496.4]
  wire [63:0] FringeZynq_io_argOuts_29_bits; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_argOuts_30_valid; // @[KCU1500.scala 21:24:@57496.4]
  wire [63:0] FringeZynq_io_argOuts_30_bits; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_argOuts_31_valid; // @[KCU1500.scala 21:24:@57496.4]
  wire [63:0] FringeZynq_io_argOuts_31_bits; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_heap_0_req_valid; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_heap_0_req_bits_allocDealloc; // @[KCU1500.scala 21:24:@57496.4]
  wire [63:0] FringeZynq_io_heap_0_req_bits_sizeAddr; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_heap_0_resp_valid; // @[KCU1500.scala 21:24:@57496.4]
  wire  FringeZynq_io_heap_0_resp_bits_allocDealloc; // @[KCU1500.scala 21:24:@57496.4]
  wire [63:0] FringeZynq_io_heap_0_resp_bits_sizeAddr; // @[KCU1500.scala 21:24:@57496.4]
  AccelUnit accel ( // @[Instantiator.scala 85:44:@57218.4]
    .clock(accel_clock),
    .reset(accel_reset),
    .io_enable(accel_io_enable),
    .io_done(accel_io_done),
    .io_reset(accel_io_reset),
    .io_memStreams_loads_0_cmd_ready(accel_io_memStreams_loads_0_cmd_ready),
    .io_memStreams_loads_0_cmd_valid(accel_io_memStreams_loads_0_cmd_valid),
    .io_memStreams_loads_0_cmd_bits_addr(accel_io_memStreams_loads_0_cmd_bits_addr),
    .io_memStreams_loads_0_cmd_bits_size(accel_io_memStreams_loads_0_cmd_bits_size),
    .io_memStreams_loads_0_data_ready(accel_io_memStreams_loads_0_data_ready),
    .io_memStreams_loads_0_data_valid(accel_io_memStreams_loads_0_data_valid),
    .io_memStreams_loads_0_data_bits_rdata_0(accel_io_memStreams_loads_0_data_bits_rdata_0),
    .io_memStreams_loads_0_data_bits_rdata_1(accel_io_memStreams_loads_0_data_bits_rdata_1),
    .io_memStreams_loads_0_data_bits_rdata_2(accel_io_memStreams_loads_0_data_bits_rdata_2),
    .io_memStreams_loads_0_data_bits_rdata_3(accel_io_memStreams_loads_0_data_bits_rdata_3),
    .io_memStreams_loads_0_data_bits_rdata_4(accel_io_memStreams_loads_0_data_bits_rdata_4),
    .io_memStreams_loads_0_data_bits_rdata_5(accel_io_memStreams_loads_0_data_bits_rdata_5),
    .io_memStreams_loads_0_data_bits_rdata_6(accel_io_memStreams_loads_0_data_bits_rdata_6),
    .io_memStreams_loads_0_data_bits_rdata_7(accel_io_memStreams_loads_0_data_bits_rdata_7),
    .io_memStreams_loads_0_data_bits_rdata_8(accel_io_memStreams_loads_0_data_bits_rdata_8),
    .io_memStreams_loads_0_data_bits_rdata_9(accel_io_memStreams_loads_0_data_bits_rdata_9),
    .io_memStreams_loads_0_data_bits_rdata_10(accel_io_memStreams_loads_0_data_bits_rdata_10),
    .io_memStreams_loads_0_data_bits_rdata_11(accel_io_memStreams_loads_0_data_bits_rdata_11),
    .io_memStreams_loads_0_data_bits_rdata_12(accel_io_memStreams_loads_0_data_bits_rdata_12),
    .io_memStreams_loads_0_data_bits_rdata_13(accel_io_memStreams_loads_0_data_bits_rdata_13),
    .io_memStreams_loads_0_data_bits_rdata_14(accel_io_memStreams_loads_0_data_bits_rdata_14),
    .io_memStreams_loads_0_data_bits_rdata_15(accel_io_memStreams_loads_0_data_bits_rdata_15),
    .io_memStreams_stores_0_cmd_ready(accel_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(accel_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(accel_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(accel_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(accel_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(accel_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(accel_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wdata_1(accel_io_memStreams_stores_0_data_bits_wdata_1),
    .io_memStreams_stores_0_data_bits_wdata_2(accel_io_memStreams_stores_0_data_bits_wdata_2),
    .io_memStreams_stores_0_data_bits_wdata_3(accel_io_memStreams_stores_0_data_bits_wdata_3),
    .io_memStreams_stores_0_data_bits_wdata_4(accel_io_memStreams_stores_0_data_bits_wdata_4),
    .io_memStreams_stores_0_data_bits_wdata_5(accel_io_memStreams_stores_0_data_bits_wdata_5),
    .io_memStreams_stores_0_data_bits_wdata_6(accel_io_memStreams_stores_0_data_bits_wdata_6),
    .io_memStreams_stores_0_data_bits_wdata_7(accel_io_memStreams_stores_0_data_bits_wdata_7),
    .io_memStreams_stores_0_data_bits_wdata_8(accel_io_memStreams_stores_0_data_bits_wdata_8),
    .io_memStreams_stores_0_data_bits_wdata_9(accel_io_memStreams_stores_0_data_bits_wdata_9),
    .io_memStreams_stores_0_data_bits_wdata_10(accel_io_memStreams_stores_0_data_bits_wdata_10),
    .io_memStreams_stores_0_data_bits_wdata_11(accel_io_memStreams_stores_0_data_bits_wdata_11),
    .io_memStreams_stores_0_data_bits_wdata_12(accel_io_memStreams_stores_0_data_bits_wdata_12),
    .io_memStreams_stores_0_data_bits_wdata_13(accel_io_memStreams_stores_0_data_bits_wdata_13),
    .io_memStreams_stores_0_data_bits_wdata_14(accel_io_memStreams_stores_0_data_bits_wdata_14),
    .io_memStreams_stores_0_data_bits_wdata_15(accel_io_memStreams_stores_0_data_bits_wdata_15),
    .io_memStreams_stores_0_data_bits_wstrb(accel_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(accel_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(accel_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(accel_io_memStreams_stores_0_wresp_bits),
    .io_memStreams_gathers_0_cmd_ready(accel_io_memStreams_gathers_0_cmd_ready),
    .io_memStreams_gathers_0_cmd_valid(accel_io_memStreams_gathers_0_cmd_valid),
    .io_memStreams_gathers_0_cmd_bits_addr_0(accel_io_memStreams_gathers_0_cmd_bits_addr_0),
    .io_memStreams_gathers_0_cmd_bits_addr_1(accel_io_memStreams_gathers_0_cmd_bits_addr_1),
    .io_memStreams_gathers_0_cmd_bits_addr_2(accel_io_memStreams_gathers_0_cmd_bits_addr_2),
    .io_memStreams_gathers_0_cmd_bits_addr_3(accel_io_memStreams_gathers_0_cmd_bits_addr_3),
    .io_memStreams_gathers_0_cmd_bits_addr_4(accel_io_memStreams_gathers_0_cmd_bits_addr_4),
    .io_memStreams_gathers_0_cmd_bits_addr_5(accel_io_memStreams_gathers_0_cmd_bits_addr_5),
    .io_memStreams_gathers_0_cmd_bits_addr_6(accel_io_memStreams_gathers_0_cmd_bits_addr_6),
    .io_memStreams_gathers_0_cmd_bits_addr_7(accel_io_memStreams_gathers_0_cmd_bits_addr_7),
    .io_memStreams_gathers_0_cmd_bits_addr_8(accel_io_memStreams_gathers_0_cmd_bits_addr_8),
    .io_memStreams_gathers_0_cmd_bits_addr_9(accel_io_memStreams_gathers_0_cmd_bits_addr_9),
    .io_memStreams_gathers_0_cmd_bits_addr_10(accel_io_memStreams_gathers_0_cmd_bits_addr_10),
    .io_memStreams_gathers_0_cmd_bits_addr_11(accel_io_memStreams_gathers_0_cmd_bits_addr_11),
    .io_memStreams_gathers_0_cmd_bits_addr_12(accel_io_memStreams_gathers_0_cmd_bits_addr_12),
    .io_memStreams_gathers_0_cmd_bits_addr_13(accel_io_memStreams_gathers_0_cmd_bits_addr_13),
    .io_memStreams_gathers_0_cmd_bits_addr_14(accel_io_memStreams_gathers_0_cmd_bits_addr_14),
    .io_memStreams_gathers_0_cmd_bits_addr_15(accel_io_memStreams_gathers_0_cmd_bits_addr_15),
    .io_memStreams_gathers_0_data_ready(accel_io_memStreams_gathers_0_data_ready),
    .io_memStreams_gathers_0_data_valid(accel_io_memStreams_gathers_0_data_valid),
    .io_memStreams_gathers_0_data_bits_0(accel_io_memStreams_gathers_0_data_bits_0),
    .io_memStreams_gathers_0_data_bits_1(accel_io_memStreams_gathers_0_data_bits_1),
    .io_memStreams_gathers_0_data_bits_2(accel_io_memStreams_gathers_0_data_bits_2),
    .io_memStreams_gathers_0_data_bits_3(accel_io_memStreams_gathers_0_data_bits_3),
    .io_memStreams_gathers_0_data_bits_4(accel_io_memStreams_gathers_0_data_bits_4),
    .io_memStreams_gathers_0_data_bits_5(accel_io_memStreams_gathers_0_data_bits_5),
    .io_memStreams_gathers_0_data_bits_6(accel_io_memStreams_gathers_0_data_bits_6),
    .io_memStreams_gathers_0_data_bits_7(accel_io_memStreams_gathers_0_data_bits_7),
    .io_memStreams_gathers_0_data_bits_8(accel_io_memStreams_gathers_0_data_bits_8),
    .io_memStreams_gathers_0_data_bits_9(accel_io_memStreams_gathers_0_data_bits_9),
    .io_memStreams_gathers_0_data_bits_10(accel_io_memStreams_gathers_0_data_bits_10),
    .io_memStreams_gathers_0_data_bits_11(accel_io_memStreams_gathers_0_data_bits_11),
    .io_memStreams_gathers_0_data_bits_12(accel_io_memStreams_gathers_0_data_bits_12),
    .io_memStreams_gathers_0_data_bits_13(accel_io_memStreams_gathers_0_data_bits_13),
    .io_memStreams_gathers_0_data_bits_14(accel_io_memStreams_gathers_0_data_bits_14),
    .io_memStreams_gathers_0_data_bits_15(accel_io_memStreams_gathers_0_data_bits_15),
    .io_memStreams_scatters_0_cmd_ready(accel_io_memStreams_scatters_0_cmd_ready),
    .io_memStreams_scatters_0_cmd_valid(accel_io_memStreams_scatters_0_cmd_valid),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_0(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_1(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_2(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_3(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_4(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_5(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_6(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_7(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_8(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_9(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_10(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_11(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_12(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_13(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_14(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_15(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15),
    .io_memStreams_scatters_0_cmd_bits_wdata_0(accel_io_memStreams_scatters_0_cmd_bits_wdata_0),
    .io_memStreams_scatters_0_cmd_bits_wdata_1(accel_io_memStreams_scatters_0_cmd_bits_wdata_1),
    .io_memStreams_scatters_0_cmd_bits_wdata_2(accel_io_memStreams_scatters_0_cmd_bits_wdata_2),
    .io_memStreams_scatters_0_cmd_bits_wdata_3(accel_io_memStreams_scatters_0_cmd_bits_wdata_3),
    .io_memStreams_scatters_0_cmd_bits_wdata_4(accel_io_memStreams_scatters_0_cmd_bits_wdata_4),
    .io_memStreams_scatters_0_cmd_bits_wdata_5(accel_io_memStreams_scatters_0_cmd_bits_wdata_5),
    .io_memStreams_scatters_0_cmd_bits_wdata_6(accel_io_memStreams_scatters_0_cmd_bits_wdata_6),
    .io_memStreams_scatters_0_cmd_bits_wdata_7(accel_io_memStreams_scatters_0_cmd_bits_wdata_7),
    .io_memStreams_scatters_0_cmd_bits_wdata_8(accel_io_memStreams_scatters_0_cmd_bits_wdata_8),
    .io_memStreams_scatters_0_cmd_bits_wdata_9(accel_io_memStreams_scatters_0_cmd_bits_wdata_9),
    .io_memStreams_scatters_0_cmd_bits_wdata_10(accel_io_memStreams_scatters_0_cmd_bits_wdata_10),
    .io_memStreams_scatters_0_cmd_bits_wdata_11(accel_io_memStreams_scatters_0_cmd_bits_wdata_11),
    .io_memStreams_scatters_0_cmd_bits_wdata_12(accel_io_memStreams_scatters_0_cmd_bits_wdata_12),
    .io_memStreams_scatters_0_cmd_bits_wdata_13(accel_io_memStreams_scatters_0_cmd_bits_wdata_13),
    .io_memStreams_scatters_0_cmd_bits_wdata_14(accel_io_memStreams_scatters_0_cmd_bits_wdata_14),
    .io_memStreams_scatters_0_cmd_bits_wdata_15(accel_io_memStreams_scatters_0_cmd_bits_wdata_15),
    .io_memStreams_scatters_0_wresp_ready(accel_io_memStreams_scatters_0_wresp_ready),
    .io_memStreams_scatters_0_wresp_valid(accel_io_memStreams_scatters_0_wresp_valid),
    .io_memStreams_scatters_0_wresp_bits(accel_io_memStreams_scatters_0_wresp_bits),
    .io_axiStreamsIn_0_TVALID(accel_io_axiStreamsIn_0_TVALID),
    .io_axiStreamsIn_0_TREADY(accel_io_axiStreamsIn_0_TREADY),
    .io_axiStreamsIn_0_TDATA(accel_io_axiStreamsIn_0_TDATA),
    .io_axiStreamsIn_0_TSTRB(accel_io_axiStreamsIn_0_TSTRB),
    .io_axiStreamsIn_0_TKEEP(accel_io_axiStreamsIn_0_TKEEP),
    .io_axiStreamsIn_0_TLAST(accel_io_axiStreamsIn_0_TLAST),
    .io_axiStreamsIn_0_TID(accel_io_axiStreamsIn_0_TID),
    .io_axiStreamsIn_0_TDEST(accel_io_axiStreamsIn_0_TDEST),
    .io_axiStreamsOut_0_TVALID(accel_io_axiStreamsOut_0_TVALID),
    .io_axiStreamsOut_0_TREADY(accel_io_axiStreamsOut_0_TREADY),
    .io_axiStreamsOut_0_TDATA(accel_io_axiStreamsOut_0_TDATA),
    .io_axiStreamsOut_0_TSTRB(accel_io_axiStreamsOut_0_TSTRB),
    .io_axiStreamsOut_0_TKEEP(accel_io_axiStreamsOut_0_TKEEP),
    .io_axiStreamsOut_0_TLAST(accel_io_axiStreamsOut_0_TLAST),
    .io_axiStreamsOut_0_TID(accel_io_axiStreamsOut_0_TID),
    .io_axiStreamsOut_0_TDEST(accel_io_axiStreamsOut_0_TDEST),
    .io_heap_0_req_valid(accel_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(accel_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(accel_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(accel_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(accel_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(accel_io_heap_0_resp_bits_sizeAddr),
    .io_argIns_0(accel_io_argIns_0),
    .io_argOuts_0_port_ready(accel_io_argOuts_0_port_ready),
    .io_argOuts_0_port_valid(accel_io_argOuts_0_port_valid),
    .io_argOuts_0_port_bits(accel_io_argOuts_0_port_bits),
    .io_argOuts_0_echo(accel_io_argOuts_0_echo),
    .io_argOuts_1_port_ready(accel_io_argOuts_1_port_ready),
    .io_argOuts_1_port_valid(accel_io_argOuts_1_port_valid),
    .io_argOuts_1_port_bits(accel_io_argOuts_1_port_bits),
    .io_argOuts_1_echo(accel_io_argOuts_1_echo),
    .io_argOuts_2_port_ready(accel_io_argOuts_2_port_ready),
    .io_argOuts_2_port_valid(accel_io_argOuts_2_port_valid),
    .io_argOuts_2_port_bits(accel_io_argOuts_2_port_bits),
    .io_argOuts_2_echo(accel_io_argOuts_2_echo),
    .io_argOuts_3_port_ready(accel_io_argOuts_3_port_ready),
    .io_argOuts_3_port_valid(accel_io_argOuts_3_port_valid),
    .io_argOuts_3_port_bits(accel_io_argOuts_3_port_bits),
    .io_argOuts_3_echo(accel_io_argOuts_3_echo),
    .io_argOuts_4_port_ready(accel_io_argOuts_4_port_ready),
    .io_argOuts_4_port_valid(accel_io_argOuts_4_port_valid),
    .io_argOuts_4_port_bits(accel_io_argOuts_4_port_bits),
    .io_argOuts_4_echo(accel_io_argOuts_4_echo),
    .io_argOuts_5_port_ready(accel_io_argOuts_5_port_ready),
    .io_argOuts_5_port_valid(accel_io_argOuts_5_port_valid),
    .io_argOuts_5_port_bits(accel_io_argOuts_5_port_bits),
    .io_argOuts_5_echo(accel_io_argOuts_5_echo),
    .io_argOuts_6_port_ready(accel_io_argOuts_6_port_ready),
    .io_argOuts_6_port_valid(accel_io_argOuts_6_port_valid),
    .io_argOuts_6_port_bits(accel_io_argOuts_6_port_bits),
    .io_argOuts_6_echo(accel_io_argOuts_6_echo),
    .io_argOuts_7_port_ready(accel_io_argOuts_7_port_ready),
    .io_argOuts_7_port_valid(accel_io_argOuts_7_port_valid),
    .io_argOuts_7_port_bits(accel_io_argOuts_7_port_bits),
    .io_argOuts_7_echo(accel_io_argOuts_7_echo),
    .io_argOuts_8_port_ready(accel_io_argOuts_8_port_ready),
    .io_argOuts_8_port_valid(accel_io_argOuts_8_port_valid),
    .io_argOuts_8_port_bits(accel_io_argOuts_8_port_bits),
    .io_argOuts_8_echo(accel_io_argOuts_8_echo),
    .io_argOuts_9_port_ready(accel_io_argOuts_9_port_ready),
    .io_argOuts_9_port_valid(accel_io_argOuts_9_port_valid),
    .io_argOuts_9_port_bits(accel_io_argOuts_9_port_bits),
    .io_argOuts_9_echo(accel_io_argOuts_9_echo),
    .io_argOuts_10_port_ready(accel_io_argOuts_10_port_ready),
    .io_argOuts_10_port_valid(accel_io_argOuts_10_port_valid),
    .io_argOuts_10_port_bits(accel_io_argOuts_10_port_bits),
    .io_argOuts_10_echo(accel_io_argOuts_10_echo),
    .io_argOuts_11_port_ready(accel_io_argOuts_11_port_ready),
    .io_argOuts_11_port_valid(accel_io_argOuts_11_port_valid),
    .io_argOuts_11_port_bits(accel_io_argOuts_11_port_bits),
    .io_argOuts_11_echo(accel_io_argOuts_11_echo),
    .io_argOuts_12_port_ready(accel_io_argOuts_12_port_ready),
    .io_argOuts_12_port_valid(accel_io_argOuts_12_port_valid),
    .io_argOuts_12_port_bits(accel_io_argOuts_12_port_bits),
    .io_argOuts_12_echo(accel_io_argOuts_12_echo),
    .io_argOuts_13_port_ready(accel_io_argOuts_13_port_ready),
    .io_argOuts_13_port_valid(accel_io_argOuts_13_port_valid),
    .io_argOuts_13_port_bits(accel_io_argOuts_13_port_bits),
    .io_argOuts_13_echo(accel_io_argOuts_13_echo),
    .io_argOuts_14_port_ready(accel_io_argOuts_14_port_ready),
    .io_argOuts_14_port_valid(accel_io_argOuts_14_port_valid),
    .io_argOuts_14_port_bits(accel_io_argOuts_14_port_bits),
    .io_argOuts_14_echo(accel_io_argOuts_14_echo),
    .io_argOuts_15_port_ready(accel_io_argOuts_15_port_ready),
    .io_argOuts_15_port_valid(accel_io_argOuts_15_port_valid),
    .io_argOuts_15_port_bits(accel_io_argOuts_15_port_bits),
    .io_argOuts_15_echo(accel_io_argOuts_15_echo),
    .io_argOuts_16_port_ready(accel_io_argOuts_16_port_ready),
    .io_argOuts_16_port_valid(accel_io_argOuts_16_port_valid),
    .io_argOuts_16_port_bits(accel_io_argOuts_16_port_bits),
    .io_argOuts_16_echo(accel_io_argOuts_16_echo),
    .io_argOuts_17_port_ready(accel_io_argOuts_17_port_ready),
    .io_argOuts_17_port_valid(accel_io_argOuts_17_port_valid),
    .io_argOuts_17_port_bits(accel_io_argOuts_17_port_bits),
    .io_argOuts_17_echo(accel_io_argOuts_17_echo),
    .io_argOuts_18_port_ready(accel_io_argOuts_18_port_ready),
    .io_argOuts_18_port_valid(accel_io_argOuts_18_port_valid),
    .io_argOuts_18_port_bits(accel_io_argOuts_18_port_bits),
    .io_argOuts_18_echo(accel_io_argOuts_18_echo),
    .io_argOuts_19_port_ready(accel_io_argOuts_19_port_ready),
    .io_argOuts_19_port_valid(accel_io_argOuts_19_port_valid),
    .io_argOuts_19_port_bits(accel_io_argOuts_19_port_bits),
    .io_argOuts_19_echo(accel_io_argOuts_19_echo),
    .io_argOuts_20_port_ready(accel_io_argOuts_20_port_ready),
    .io_argOuts_20_port_valid(accel_io_argOuts_20_port_valid),
    .io_argOuts_20_port_bits(accel_io_argOuts_20_port_bits),
    .io_argOuts_20_echo(accel_io_argOuts_20_echo),
    .io_argOuts_21_port_ready(accel_io_argOuts_21_port_ready),
    .io_argOuts_21_port_valid(accel_io_argOuts_21_port_valid),
    .io_argOuts_21_port_bits(accel_io_argOuts_21_port_bits),
    .io_argOuts_21_echo(accel_io_argOuts_21_echo),
    .io_argOuts_22_port_ready(accel_io_argOuts_22_port_ready),
    .io_argOuts_22_port_valid(accel_io_argOuts_22_port_valid),
    .io_argOuts_22_port_bits(accel_io_argOuts_22_port_bits),
    .io_argOuts_22_echo(accel_io_argOuts_22_echo),
    .io_argOuts_23_port_ready(accel_io_argOuts_23_port_ready),
    .io_argOuts_23_port_valid(accel_io_argOuts_23_port_valid),
    .io_argOuts_23_port_bits(accel_io_argOuts_23_port_bits),
    .io_argOuts_23_echo(accel_io_argOuts_23_echo),
    .io_argOuts_24_port_ready(accel_io_argOuts_24_port_ready),
    .io_argOuts_24_port_valid(accel_io_argOuts_24_port_valid),
    .io_argOuts_24_port_bits(accel_io_argOuts_24_port_bits),
    .io_argOuts_24_echo(accel_io_argOuts_24_echo),
    .io_argOuts_25_port_ready(accel_io_argOuts_25_port_ready),
    .io_argOuts_25_port_valid(accel_io_argOuts_25_port_valid),
    .io_argOuts_25_port_bits(accel_io_argOuts_25_port_bits),
    .io_argOuts_25_echo(accel_io_argOuts_25_echo),
    .io_argOuts_26_port_ready(accel_io_argOuts_26_port_ready),
    .io_argOuts_26_port_valid(accel_io_argOuts_26_port_valid),
    .io_argOuts_26_port_bits(accel_io_argOuts_26_port_bits),
    .io_argOuts_26_echo(accel_io_argOuts_26_echo),
    .io_argOuts_27_port_ready(accel_io_argOuts_27_port_ready),
    .io_argOuts_27_port_valid(accel_io_argOuts_27_port_valid),
    .io_argOuts_27_port_bits(accel_io_argOuts_27_port_bits),
    .io_argOuts_27_echo(accel_io_argOuts_27_echo),
    .io_argOuts_28_port_ready(accel_io_argOuts_28_port_ready),
    .io_argOuts_28_port_valid(accel_io_argOuts_28_port_valid),
    .io_argOuts_28_port_bits(accel_io_argOuts_28_port_bits),
    .io_argOuts_28_echo(accel_io_argOuts_28_echo),
    .io_argOuts_29_port_ready(accel_io_argOuts_29_port_ready),
    .io_argOuts_29_port_valid(accel_io_argOuts_29_port_valid),
    .io_argOuts_29_port_bits(accel_io_argOuts_29_port_bits),
    .io_argOuts_29_echo(accel_io_argOuts_29_echo),
    .io_argOuts_30_port_ready(accel_io_argOuts_30_port_ready),
    .io_argOuts_30_port_valid(accel_io_argOuts_30_port_valid),
    .io_argOuts_30_port_bits(accel_io_argOuts_30_port_bits),
    .io_argOuts_30_echo(accel_io_argOuts_30_echo),
    .io_argOuts_31_port_ready(accel_io_argOuts_31_port_ready),
    .io_argOuts_31_port_valid(accel_io_argOuts_31_port_valid),
    .io_argOuts_31_port_bits(accel_io_argOuts_31_port_bits),
    .io_argOuts_31_echo(accel_io_argOuts_31_echo)
  );
  FringeZynq FringeZynq ( // @[KCU1500.scala 21:24:@57496.4]
    .clock(FringeZynq_clock),
    .reset(FringeZynq_reset),
    .io_S_AXI_AWADDR(FringeZynq_io_S_AXI_AWADDR),
    .io_S_AXI_AWPROT(FringeZynq_io_S_AXI_AWPROT),
    .io_S_AXI_AWVALID(FringeZynq_io_S_AXI_AWVALID),
    .io_S_AXI_AWREADY(FringeZynq_io_S_AXI_AWREADY),
    .io_S_AXI_ARADDR(FringeZynq_io_S_AXI_ARADDR),
    .io_S_AXI_ARPROT(FringeZynq_io_S_AXI_ARPROT),
    .io_S_AXI_ARVALID(FringeZynq_io_S_AXI_ARVALID),
    .io_S_AXI_ARREADY(FringeZynq_io_S_AXI_ARREADY),
    .io_S_AXI_WDATA(FringeZynq_io_S_AXI_WDATA),
    .io_S_AXI_WSTRB(FringeZynq_io_S_AXI_WSTRB),
    .io_S_AXI_WVALID(FringeZynq_io_S_AXI_WVALID),
    .io_S_AXI_WREADY(FringeZynq_io_S_AXI_WREADY),
    .io_S_AXI_RDATA(FringeZynq_io_S_AXI_RDATA),
    .io_S_AXI_RRESP(FringeZynq_io_S_AXI_RRESP),
    .io_S_AXI_RVALID(FringeZynq_io_S_AXI_RVALID),
    .io_S_AXI_RREADY(FringeZynq_io_S_AXI_RREADY),
    .io_S_AXI_BRESP(FringeZynq_io_S_AXI_BRESP),
    .io_S_AXI_BVALID(FringeZynq_io_S_AXI_BVALID),
    .io_S_AXI_BREADY(FringeZynq_io_S_AXI_BREADY),
    .io_M_AXI_0_AWLEN(FringeZynq_io_M_AXI_0_AWLEN),
    .io_M_AXI_0_ARLEN(FringeZynq_io_M_AXI_0_ARLEN),
    .io_enable(FringeZynq_io_enable),
    .io_done(FringeZynq_io_done),
    .io_reset(FringeZynq_io_reset),
    .io_argIns_0(FringeZynq_io_argIns_0),
    .io_argOuts_0_valid(FringeZynq_io_argOuts_0_valid),
    .io_argOuts_0_bits(FringeZynq_io_argOuts_0_bits),
    .io_argOuts_1_valid(FringeZynq_io_argOuts_1_valid),
    .io_argOuts_1_bits(FringeZynq_io_argOuts_1_bits),
    .io_argOuts_2_valid(FringeZynq_io_argOuts_2_valid),
    .io_argOuts_2_bits(FringeZynq_io_argOuts_2_bits),
    .io_argOuts_3_valid(FringeZynq_io_argOuts_3_valid),
    .io_argOuts_3_bits(FringeZynq_io_argOuts_3_bits),
    .io_argOuts_4_valid(FringeZynq_io_argOuts_4_valid),
    .io_argOuts_4_bits(FringeZynq_io_argOuts_4_bits),
    .io_argOuts_5_valid(FringeZynq_io_argOuts_5_valid),
    .io_argOuts_5_bits(FringeZynq_io_argOuts_5_bits),
    .io_argOuts_6_valid(FringeZynq_io_argOuts_6_valid),
    .io_argOuts_6_bits(FringeZynq_io_argOuts_6_bits),
    .io_argOuts_7_valid(FringeZynq_io_argOuts_7_valid),
    .io_argOuts_7_bits(FringeZynq_io_argOuts_7_bits),
    .io_argOuts_8_valid(FringeZynq_io_argOuts_8_valid),
    .io_argOuts_8_bits(FringeZynq_io_argOuts_8_bits),
    .io_argOuts_9_valid(FringeZynq_io_argOuts_9_valid),
    .io_argOuts_9_bits(FringeZynq_io_argOuts_9_bits),
    .io_argOuts_10_valid(FringeZynq_io_argOuts_10_valid),
    .io_argOuts_10_bits(FringeZynq_io_argOuts_10_bits),
    .io_argOuts_11_valid(FringeZynq_io_argOuts_11_valid),
    .io_argOuts_11_bits(FringeZynq_io_argOuts_11_bits),
    .io_argOuts_12_valid(FringeZynq_io_argOuts_12_valid),
    .io_argOuts_12_bits(FringeZynq_io_argOuts_12_bits),
    .io_argOuts_13_valid(FringeZynq_io_argOuts_13_valid),
    .io_argOuts_13_bits(FringeZynq_io_argOuts_13_bits),
    .io_argOuts_14_valid(FringeZynq_io_argOuts_14_valid),
    .io_argOuts_14_bits(FringeZynq_io_argOuts_14_bits),
    .io_argOuts_15_valid(FringeZynq_io_argOuts_15_valid),
    .io_argOuts_15_bits(FringeZynq_io_argOuts_15_bits),
    .io_argOuts_16_valid(FringeZynq_io_argOuts_16_valid),
    .io_argOuts_16_bits(FringeZynq_io_argOuts_16_bits),
    .io_argOuts_17_valid(FringeZynq_io_argOuts_17_valid),
    .io_argOuts_17_bits(FringeZynq_io_argOuts_17_bits),
    .io_argOuts_18_valid(FringeZynq_io_argOuts_18_valid),
    .io_argOuts_18_bits(FringeZynq_io_argOuts_18_bits),
    .io_argOuts_19_valid(FringeZynq_io_argOuts_19_valid),
    .io_argOuts_19_bits(FringeZynq_io_argOuts_19_bits),
    .io_argOuts_20_valid(FringeZynq_io_argOuts_20_valid),
    .io_argOuts_20_bits(FringeZynq_io_argOuts_20_bits),
    .io_argOuts_21_valid(FringeZynq_io_argOuts_21_valid),
    .io_argOuts_21_bits(FringeZynq_io_argOuts_21_bits),
    .io_argOuts_22_valid(FringeZynq_io_argOuts_22_valid),
    .io_argOuts_22_bits(FringeZynq_io_argOuts_22_bits),
    .io_argOuts_23_valid(FringeZynq_io_argOuts_23_valid),
    .io_argOuts_23_bits(FringeZynq_io_argOuts_23_bits),
    .io_argOuts_24_valid(FringeZynq_io_argOuts_24_valid),
    .io_argOuts_24_bits(FringeZynq_io_argOuts_24_bits),
    .io_argOuts_25_valid(FringeZynq_io_argOuts_25_valid),
    .io_argOuts_25_bits(FringeZynq_io_argOuts_25_bits),
    .io_argOuts_26_valid(FringeZynq_io_argOuts_26_valid),
    .io_argOuts_26_bits(FringeZynq_io_argOuts_26_bits),
    .io_argOuts_27_valid(FringeZynq_io_argOuts_27_valid),
    .io_argOuts_27_bits(FringeZynq_io_argOuts_27_bits),
    .io_argOuts_28_valid(FringeZynq_io_argOuts_28_valid),
    .io_argOuts_28_bits(FringeZynq_io_argOuts_28_bits),
    .io_argOuts_29_valid(FringeZynq_io_argOuts_29_valid),
    .io_argOuts_29_bits(FringeZynq_io_argOuts_29_bits),
    .io_argOuts_30_valid(FringeZynq_io_argOuts_30_valid),
    .io_argOuts_30_bits(FringeZynq_io_argOuts_30_bits),
    .io_argOuts_31_valid(FringeZynq_io_argOuts_31_valid),
    .io_argOuts_31_bits(FringeZynq_io_argOuts_31_bits),
    .io_heap_0_req_valid(FringeZynq_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(FringeZynq_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(FringeZynq_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(FringeZynq_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(FringeZynq_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(FringeZynq_io_heap_0_resp_bits_sizeAddr)
  );
  assign io_rdata = 1'h0;
  assign io_S_AXI_AWREADY = FringeZynq_io_S_AXI_AWREADY; // @[KCU1500.scala 24:21:@57514.4]
  assign io_S_AXI_ARREADY = FringeZynq_io_S_AXI_ARREADY; // @[KCU1500.scala 24:21:@57510.4]
  assign io_S_AXI_WREADY = FringeZynq_io_S_AXI_WREADY; // @[KCU1500.scala 24:21:@57506.4]
  assign io_S_AXI_RDATA = FringeZynq_io_S_AXI_RDATA; // @[KCU1500.scala 24:21:@57505.4]
  assign io_S_AXI_RRESP = FringeZynq_io_S_AXI_RRESP; // @[KCU1500.scala 24:21:@57504.4]
  assign io_S_AXI_RVALID = FringeZynq_io_S_AXI_RVALID; // @[KCU1500.scala 24:21:@57503.4]
  assign io_S_AXI_BRESP = FringeZynq_io_S_AXI_BRESP; // @[KCU1500.scala 24:21:@57501.4]
  assign io_S_AXI_BVALID = FringeZynq_io_S_AXI_BVALID; // @[KCU1500.scala 24:21:@57500.4]
  assign io_M_AXI_0_AWID = 4'h0; // @[KCU1500.scala 31:14:@57574.4]
  assign io_M_AXI_0_AWUSER = 4'h0; // @[KCU1500.scala 31:14:@57573.4]
  assign io_M_AXI_0_AWADDR = 32'h0; // @[KCU1500.scala 31:14:@57572.4]
  assign io_M_AXI_0_AWLEN = FringeZynq_io_M_AXI_0_AWLEN; // @[KCU1500.scala 31:14:@57571.4]
  assign io_M_AXI_0_AWSIZE = 3'h6; // @[KCU1500.scala 31:14:@57570.4]
  assign io_M_AXI_0_AWBURST = 2'h1; // @[KCU1500.scala 31:14:@57569.4]
  assign io_M_AXI_0_AWLOCK = 1'h0; // @[KCU1500.scala 31:14:@57568.4]
  assign io_M_AXI_0_AWCACHE = 4'h3; // @[KCU1500.scala 31:14:@57567.4]
  assign io_M_AXI_0_AWPROT = 3'h0; // @[KCU1500.scala 31:14:@57566.4]
  assign io_M_AXI_0_AWQOS = 4'h0; // @[KCU1500.scala 31:14:@57565.4]
  assign io_M_AXI_0_AWVALID = 1'h0; // @[KCU1500.scala 31:14:@57564.4]
  assign io_M_AXI_0_ARID = 4'h0; // @[KCU1500.scala 31:14:@57562.4]
  assign io_M_AXI_0_ARUSER = 4'h0; // @[KCU1500.scala 31:14:@57561.4]
  assign io_M_AXI_0_ARADDR = 32'h0; // @[KCU1500.scala 31:14:@57560.4]
  assign io_M_AXI_0_ARLEN = FringeZynq_io_M_AXI_0_ARLEN; // @[KCU1500.scala 31:14:@57559.4]
  assign io_M_AXI_0_ARSIZE = 3'h6; // @[KCU1500.scala 31:14:@57558.4]
  assign io_M_AXI_0_ARBURST = 2'h1; // @[KCU1500.scala 31:14:@57557.4]
  assign io_M_AXI_0_ARLOCK = 1'h0; // @[KCU1500.scala 31:14:@57556.4]
  assign io_M_AXI_0_ARCACHE = 4'h3; // @[KCU1500.scala 31:14:@57555.4]
  assign io_M_AXI_0_ARPROT = 3'h0; // @[KCU1500.scala 31:14:@57554.4]
  assign io_M_AXI_0_ARQOS = 4'h0; // @[KCU1500.scala 31:14:@57553.4]
  assign io_M_AXI_0_ARVALID = 1'h0; // @[KCU1500.scala 31:14:@57552.4]
  assign io_M_AXI_0_WDATA = 512'h0; // @[KCU1500.scala 31:14:@57550.4]
  assign io_M_AXI_0_WSTRB = 64'h0; // @[KCU1500.scala 31:14:@57549.4]
  assign io_M_AXI_0_WLAST = 1'h0; // @[KCU1500.scala 31:14:@57548.4]
  assign io_M_AXI_0_WVALID = 1'h0; // @[KCU1500.scala 31:14:@57547.4]
  assign io_M_AXI_0_RREADY = 1'h0; // @[KCU1500.scala 31:14:@57539.4]
  assign io_M_AXI_0_BREADY = 1'h0; // @[KCU1500.scala 31:14:@57534.4]
  assign io_AXIS_IN_TREADY = accel_io_axiStreamsIn_0_TREADY; // @[KCU1500.scala 27:16:@57524.4]
  assign io_AXIS_OUT_TVALID = accel_io_axiStreamsOut_0_TVALID; // @[KCU1500.scala 28:17:@57533.4]
  assign io_AXIS_OUT_TDATA = accel_io_axiStreamsOut_0_TDATA; // @[KCU1500.scala 28:17:@57531.4]
  assign io_AXIS_OUT_TSTRB = accel_io_axiStreamsOut_0_TSTRB; // @[KCU1500.scala 28:17:@57530.4]
  assign io_AXIS_OUT_TKEEP = accel_io_axiStreamsOut_0_TKEEP; // @[KCU1500.scala 28:17:@57529.4]
  assign io_AXIS_OUT_TLAST = accel_io_axiStreamsOut_0_TLAST; // @[KCU1500.scala 28:17:@57528.4]
  assign io_AXIS_OUT_TID = accel_io_axiStreamsOut_0_TID[3:0]; // @[KCU1500.scala 28:17:@57527.4]
  assign io_AXIS_OUT_TDEST = accel_io_axiStreamsOut_0_TDEST[3:0]; // @[KCU1500.scala 28:17:@57526.4]
  assign accel_clock = clock; // @[:@57219.4]
  assign accel_reset = FringeZynq_io_reset; // @[:@57220.4 KCU1500.scala 61:17:@57969.4]
  assign accel_io_enable = FringeZynq_io_enable; // @[KCU1500.scala 58:21:@57965.4]
  assign accel_io_reset = 1'h0;
  assign accel_io_memStreams_loads_0_cmd_ready = 1'h0; // @[KCU1500.scala 56:26:@57958.4]
  assign accel_io_memStreams_loads_0_data_valid = 1'h0; // @[KCU1500.scala 56:26:@57953.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_0 = 32'h0; // @[KCU1500.scala 56:26:@57937.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_1 = 32'h0; // @[KCU1500.scala 56:26:@57938.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_2 = 32'h0; // @[KCU1500.scala 56:26:@57939.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_3 = 32'h0; // @[KCU1500.scala 56:26:@57940.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_4 = 32'h0; // @[KCU1500.scala 56:26:@57941.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_5 = 32'h0; // @[KCU1500.scala 56:26:@57942.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_6 = 32'h0; // @[KCU1500.scala 56:26:@57943.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_7 = 32'h0; // @[KCU1500.scala 56:26:@57944.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_8 = 32'h0; // @[KCU1500.scala 56:26:@57945.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_9 = 32'h0; // @[KCU1500.scala 56:26:@57946.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_10 = 32'h0; // @[KCU1500.scala 56:26:@57947.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_11 = 32'h0; // @[KCU1500.scala 56:26:@57948.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_12 = 32'h0; // @[KCU1500.scala 56:26:@57949.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_13 = 32'h0; // @[KCU1500.scala 56:26:@57950.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_14 = 32'h0; // @[KCU1500.scala 56:26:@57951.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_15 = 32'h0; // @[KCU1500.scala 56:26:@57952.4]
  assign accel_io_memStreams_stores_0_cmd_ready = 1'h0; // @[KCU1500.scala 56:26:@57936.4]
  assign accel_io_memStreams_stores_0_data_ready = 1'h0; // @[KCU1500.scala 56:26:@57932.4]
  assign accel_io_memStreams_stores_0_wresp_valid = 1'h0; // @[KCU1500.scala 56:26:@57912.4]
  assign accel_io_memStreams_stores_0_wresp_bits = 1'h0; // @[KCU1500.scala 56:26:@57911.4]
  assign accel_io_memStreams_gathers_0_cmd_ready = 1'h0; // @[KCU1500.scala 56:26:@57910.4]
  assign accel_io_memStreams_gathers_0_data_valid = 1'h0; // @[KCU1500.scala 56:26:@57891.4]
  assign accel_io_memStreams_gathers_0_data_bits_0 = 32'h0; // @[KCU1500.scala 56:26:@57875.4]
  assign accel_io_memStreams_gathers_0_data_bits_1 = 32'h0; // @[KCU1500.scala 56:26:@57876.4]
  assign accel_io_memStreams_gathers_0_data_bits_2 = 32'h0; // @[KCU1500.scala 56:26:@57877.4]
  assign accel_io_memStreams_gathers_0_data_bits_3 = 32'h0; // @[KCU1500.scala 56:26:@57878.4]
  assign accel_io_memStreams_gathers_0_data_bits_4 = 32'h0; // @[KCU1500.scala 56:26:@57879.4]
  assign accel_io_memStreams_gathers_0_data_bits_5 = 32'h0; // @[KCU1500.scala 56:26:@57880.4]
  assign accel_io_memStreams_gathers_0_data_bits_6 = 32'h0; // @[KCU1500.scala 56:26:@57881.4]
  assign accel_io_memStreams_gathers_0_data_bits_7 = 32'h0; // @[KCU1500.scala 56:26:@57882.4]
  assign accel_io_memStreams_gathers_0_data_bits_8 = 32'h0; // @[KCU1500.scala 56:26:@57883.4]
  assign accel_io_memStreams_gathers_0_data_bits_9 = 32'h0; // @[KCU1500.scala 56:26:@57884.4]
  assign accel_io_memStreams_gathers_0_data_bits_10 = 32'h0; // @[KCU1500.scala 56:26:@57885.4]
  assign accel_io_memStreams_gathers_0_data_bits_11 = 32'h0; // @[KCU1500.scala 56:26:@57886.4]
  assign accel_io_memStreams_gathers_0_data_bits_12 = 32'h0; // @[KCU1500.scala 56:26:@57887.4]
  assign accel_io_memStreams_gathers_0_data_bits_13 = 32'h0; // @[KCU1500.scala 56:26:@57888.4]
  assign accel_io_memStreams_gathers_0_data_bits_14 = 32'h0; // @[KCU1500.scala 56:26:@57889.4]
  assign accel_io_memStreams_gathers_0_data_bits_15 = 32'h0; // @[KCU1500.scala 56:26:@57890.4]
  assign accel_io_memStreams_scatters_0_cmd_ready = 1'h0; // @[KCU1500.scala 56:26:@57874.4]
  assign accel_io_memStreams_scatters_0_wresp_valid = 1'h0; // @[KCU1500.scala 56:26:@57839.4]
  assign accel_io_memStreams_scatters_0_wresp_bits = 1'h0; // @[KCU1500.scala 56:26:@57838.4]
  assign accel_io_axiStreamsIn_0_TVALID = io_AXIS_IN_TVALID; // @[KCU1500.scala 27:16:@57525.4]
  assign accel_io_axiStreamsIn_0_TDATA = io_AXIS_IN_TDATA; // @[KCU1500.scala 27:16:@57523.4]
  assign accel_io_axiStreamsIn_0_TSTRB = io_AXIS_IN_TSTRB; // @[KCU1500.scala 27:16:@57522.4]
  assign accel_io_axiStreamsIn_0_TKEEP = io_AXIS_IN_TKEEP; // @[KCU1500.scala 27:16:@57521.4]
  assign accel_io_axiStreamsIn_0_TLAST = io_AXIS_IN_TLAST; // @[KCU1500.scala 27:16:@57520.4]
  assign accel_io_axiStreamsIn_0_TID = {{4'd0}, io_AXIS_IN_TID}; // @[KCU1500.scala 27:16:@57519.4]
  assign accel_io_axiStreamsIn_0_TDEST = {{4'd0}, io_AXIS_IN_TDEST}; // @[KCU1500.scala 27:16:@57518.4]
  assign accel_io_axiStreamsOut_0_TREADY = io_AXIS_OUT_TREADY; // @[KCU1500.scala 28:17:@57532.4]
  assign accel_io_heap_0_resp_valid = FringeZynq_io_heap_0_resp_valid; // @[KCU1500.scala 57:20:@57961.4]
  assign accel_io_heap_0_resp_bits_allocDealloc = FringeZynq_io_heap_0_resp_bits_allocDealloc; // @[KCU1500.scala 57:20:@57960.4]
  assign accel_io_heap_0_resp_bits_sizeAddr = FringeZynq_io_heap_0_resp_bits_sizeAddr; // @[KCU1500.scala 57:20:@57959.4]
  assign accel_io_argIns_0 = FringeZynq_io_argIns_0; // @[KCU1500.scala 41:21:@57740.4]
  assign accel_io_argOuts_0_port_ready = 1'h0;
  assign accel_io_argOuts_0_echo = 64'h0; // @[KCU1500.scala 47:24:@57805.4]
  assign accel_io_argOuts_1_port_ready = 1'h0;
  assign accel_io_argOuts_1_echo = 64'h0; // @[KCU1500.scala 47:24:@57806.4]
  assign accel_io_argOuts_2_port_ready = 1'h0;
  assign accel_io_argOuts_2_echo = 64'h0; // @[KCU1500.scala 47:24:@57807.4]
  assign accel_io_argOuts_3_port_ready = 1'h0;
  assign accel_io_argOuts_3_echo = 64'h0; // @[KCU1500.scala 47:24:@57808.4]
  assign accel_io_argOuts_4_port_ready = 1'h0;
  assign accel_io_argOuts_4_echo = 64'h0; // @[KCU1500.scala 47:24:@57809.4]
  assign accel_io_argOuts_5_port_ready = 1'h0;
  assign accel_io_argOuts_5_echo = 64'h0; // @[KCU1500.scala 47:24:@57810.4]
  assign accel_io_argOuts_6_port_ready = 1'h0;
  assign accel_io_argOuts_6_echo = 64'h0; // @[KCU1500.scala 47:24:@57811.4]
  assign accel_io_argOuts_7_port_ready = 1'h0;
  assign accel_io_argOuts_7_echo = 64'h0; // @[KCU1500.scala 47:24:@57812.4]
  assign accel_io_argOuts_8_port_ready = 1'h0;
  assign accel_io_argOuts_8_echo = 64'h0; // @[KCU1500.scala 47:24:@57813.4]
  assign accel_io_argOuts_9_port_ready = 1'h0;
  assign accel_io_argOuts_9_echo = 64'h0; // @[KCU1500.scala 47:24:@57814.4]
  assign accel_io_argOuts_10_port_ready = 1'h0;
  assign accel_io_argOuts_10_echo = 64'h0; // @[KCU1500.scala 47:24:@57815.4]
  assign accel_io_argOuts_11_port_ready = 1'h0;
  assign accel_io_argOuts_11_echo = 64'h0; // @[KCU1500.scala 47:24:@57816.4]
  assign accel_io_argOuts_12_port_ready = 1'h0;
  assign accel_io_argOuts_12_echo = 64'h0; // @[KCU1500.scala 47:24:@57817.4]
  assign accel_io_argOuts_13_port_ready = 1'h0;
  assign accel_io_argOuts_13_echo = 64'h0; // @[KCU1500.scala 47:24:@57818.4]
  assign accel_io_argOuts_14_port_ready = 1'h0;
  assign accel_io_argOuts_14_echo = 64'h0; // @[KCU1500.scala 47:24:@57819.4]
  assign accel_io_argOuts_15_port_ready = 1'h0;
  assign accel_io_argOuts_15_echo = 64'h0; // @[KCU1500.scala 47:24:@57820.4]
  assign accel_io_argOuts_16_port_ready = 1'h0;
  assign accel_io_argOuts_16_echo = 64'h0; // @[KCU1500.scala 47:24:@57821.4]
  assign accel_io_argOuts_17_port_ready = 1'h0;
  assign accel_io_argOuts_17_echo = 64'h0; // @[KCU1500.scala 47:24:@57822.4]
  assign accel_io_argOuts_18_port_ready = 1'h0;
  assign accel_io_argOuts_18_echo = 64'h0; // @[KCU1500.scala 47:24:@57823.4]
  assign accel_io_argOuts_19_port_ready = 1'h0;
  assign accel_io_argOuts_19_echo = 64'h0; // @[KCU1500.scala 47:24:@57824.4]
  assign accel_io_argOuts_20_port_ready = 1'h0;
  assign accel_io_argOuts_20_echo = 64'h0; // @[KCU1500.scala 47:24:@57825.4]
  assign accel_io_argOuts_21_port_ready = 1'h0;
  assign accel_io_argOuts_21_echo = 64'h0; // @[KCU1500.scala 47:24:@57826.4]
  assign accel_io_argOuts_22_port_ready = 1'h0;
  assign accel_io_argOuts_22_echo = 64'h0; // @[KCU1500.scala 47:24:@57827.4]
  assign accel_io_argOuts_23_port_ready = 1'h0;
  assign accel_io_argOuts_23_echo = 64'h0; // @[KCU1500.scala 47:24:@57828.4]
  assign accel_io_argOuts_24_port_ready = 1'h0;
  assign accel_io_argOuts_24_echo = 64'h0; // @[KCU1500.scala 47:24:@57829.4]
  assign accel_io_argOuts_25_port_ready = 1'h0;
  assign accel_io_argOuts_25_echo = 64'h0; // @[KCU1500.scala 47:24:@57830.4]
  assign accel_io_argOuts_26_port_ready = 1'h0;
  assign accel_io_argOuts_26_echo = 64'h0; // @[KCU1500.scala 47:24:@57831.4]
  assign accel_io_argOuts_27_port_ready = 1'h0;
  assign accel_io_argOuts_27_echo = 64'h0; // @[KCU1500.scala 47:24:@57832.4]
  assign accel_io_argOuts_28_port_ready = 1'h0;
  assign accel_io_argOuts_28_echo = 64'h0; // @[KCU1500.scala 47:24:@57833.4]
  assign accel_io_argOuts_29_port_ready = 1'h0;
  assign accel_io_argOuts_29_echo = 64'h0; // @[KCU1500.scala 47:24:@57834.4]
  assign accel_io_argOuts_30_port_ready = 1'h0;
  assign accel_io_argOuts_30_echo = 64'h0; // @[KCU1500.scala 47:24:@57835.4]
  assign accel_io_argOuts_31_port_ready = 1'h0;
  assign accel_io_argOuts_31_echo = 64'h0; // @[KCU1500.scala 47:24:@57836.4]
  assign FringeZynq_clock = clock; // @[:@57497.4]
  assign FringeZynq_reset = reset; // @[:@57498.4 KCU1500.scala 60:18:@57968.4]
  assign FringeZynq_io_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[KCU1500.scala 24:21:@57517.4]
  assign FringeZynq_io_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[KCU1500.scala 24:21:@57516.4]
  assign FringeZynq_io_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[KCU1500.scala 24:21:@57515.4]
  assign FringeZynq_io_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[KCU1500.scala 24:21:@57513.4]
  assign FringeZynq_io_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[KCU1500.scala 24:21:@57512.4]
  assign FringeZynq_io_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[KCU1500.scala 24:21:@57511.4]
  assign FringeZynq_io_S_AXI_WDATA = io_S_AXI_WDATA; // @[KCU1500.scala 24:21:@57509.4]
  assign FringeZynq_io_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[KCU1500.scala 24:21:@57508.4]
  assign FringeZynq_io_S_AXI_WVALID = io_S_AXI_WVALID; // @[KCU1500.scala 24:21:@57507.4]
  assign FringeZynq_io_S_AXI_RREADY = io_S_AXI_RREADY; // @[KCU1500.scala 24:21:@57502.4]
  assign FringeZynq_io_S_AXI_BREADY = io_S_AXI_BREADY; // @[KCU1500.scala 24:21:@57499.4]
  assign FringeZynq_io_done = accel_io_done; // @[KCU1500.scala 59:20:@57966.4]
  assign FringeZynq_io_argOuts_0_valid = accel_io_argOuts_0_port_valid; // @[KCU1500.scala 44:26:@57742.4]
  assign FringeZynq_io_argOuts_0_bits = accel_io_argOuts_0_port_bits; // @[KCU1500.scala 43:25:@57741.4]
  assign FringeZynq_io_argOuts_1_valid = accel_io_argOuts_1_port_valid; // @[KCU1500.scala 44:26:@57744.4]
  assign FringeZynq_io_argOuts_1_bits = accel_io_argOuts_1_port_bits; // @[KCU1500.scala 43:25:@57743.4]
  assign FringeZynq_io_argOuts_2_valid = accel_io_argOuts_2_port_valid; // @[KCU1500.scala 44:26:@57746.4]
  assign FringeZynq_io_argOuts_2_bits = accel_io_argOuts_2_port_bits; // @[KCU1500.scala 43:25:@57745.4]
  assign FringeZynq_io_argOuts_3_valid = accel_io_argOuts_3_port_valid; // @[KCU1500.scala 44:26:@57748.4]
  assign FringeZynq_io_argOuts_3_bits = accel_io_argOuts_3_port_bits; // @[KCU1500.scala 43:25:@57747.4]
  assign FringeZynq_io_argOuts_4_valid = accel_io_argOuts_4_port_valid; // @[KCU1500.scala 44:26:@57750.4]
  assign FringeZynq_io_argOuts_4_bits = accel_io_argOuts_4_port_bits; // @[KCU1500.scala 43:25:@57749.4]
  assign FringeZynq_io_argOuts_5_valid = accel_io_argOuts_5_port_valid; // @[KCU1500.scala 44:26:@57752.4]
  assign FringeZynq_io_argOuts_5_bits = accel_io_argOuts_5_port_bits; // @[KCU1500.scala 43:25:@57751.4]
  assign FringeZynq_io_argOuts_6_valid = accel_io_argOuts_6_port_valid; // @[KCU1500.scala 44:26:@57754.4]
  assign FringeZynq_io_argOuts_6_bits = accel_io_argOuts_6_port_bits; // @[KCU1500.scala 43:25:@57753.4]
  assign FringeZynq_io_argOuts_7_valid = accel_io_argOuts_7_port_valid; // @[KCU1500.scala 44:26:@57756.4]
  assign FringeZynq_io_argOuts_7_bits = accel_io_argOuts_7_port_bits; // @[KCU1500.scala 43:25:@57755.4]
  assign FringeZynq_io_argOuts_8_valid = accel_io_argOuts_8_port_valid; // @[KCU1500.scala 44:26:@57758.4]
  assign FringeZynq_io_argOuts_8_bits = accel_io_argOuts_8_port_bits; // @[KCU1500.scala 43:25:@57757.4]
  assign FringeZynq_io_argOuts_9_valid = accel_io_argOuts_9_port_valid; // @[KCU1500.scala 44:26:@57760.4]
  assign FringeZynq_io_argOuts_9_bits = accel_io_argOuts_9_port_bits; // @[KCU1500.scala 43:25:@57759.4]
  assign FringeZynq_io_argOuts_10_valid = accel_io_argOuts_10_port_valid; // @[KCU1500.scala 44:26:@57762.4]
  assign FringeZynq_io_argOuts_10_bits = accel_io_argOuts_10_port_bits; // @[KCU1500.scala 43:25:@57761.4]
  assign FringeZynq_io_argOuts_11_valid = accel_io_argOuts_11_port_valid; // @[KCU1500.scala 44:26:@57764.4]
  assign FringeZynq_io_argOuts_11_bits = accel_io_argOuts_11_port_bits; // @[KCU1500.scala 43:25:@57763.4]
  assign FringeZynq_io_argOuts_12_valid = accel_io_argOuts_12_port_valid; // @[KCU1500.scala 44:26:@57766.4]
  assign FringeZynq_io_argOuts_12_bits = accel_io_argOuts_12_port_bits; // @[KCU1500.scala 43:25:@57765.4]
  assign FringeZynq_io_argOuts_13_valid = accel_io_argOuts_13_port_valid; // @[KCU1500.scala 44:26:@57768.4]
  assign FringeZynq_io_argOuts_13_bits = accel_io_argOuts_13_port_bits; // @[KCU1500.scala 43:25:@57767.4]
  assign FringeZynq_io_argOuts_14_valid = accel_io_argOuts_14_port_valid; // @[KCU1500.scala 44:26:@57770.4]
  assign FringeZynq_io_argOuts_14_bits = accel_io_argOuts_14_port_bits; // @[KCU1500.scala 43:25:@57769.4]
  assign FringeZynq_io_argOuts_15_valid = accel_io_argOuts_15_port_valid; // @[KCU1500.scala 44:26:@57772.4]
  assign FringeZynq_io_argOuts_15_bits = accel_io_argOuts_15_port_bits; // @[KCU1500.scala 43:25:@57771.4]
  assign FringeZynq_io_argOuts_16_valid = accel_io_argOuts_16_port_valid; // @[KCU1500.scala 44:26:@57774.4]
  assign FringeZynq_io_argOuts_16_bits = accel_io_argOuts_16_port_bits; // @[KCU1500.scala 43:25:@57773.4]
  assign FringeZynq_io_argOuts_17_valid = accel_io_argOuts_17_port_valid; // @[KCU1500.scala 44:26:@57776.4]
  assign FringeZynq_io_argOuts_17_bits = accel_io_argOuts_17_port_bits; // @[KCU1500.scala 43:25:@57775.4]
  assign FringeZynq_io_argOuts_18_valid = accel_io_argOuts_18_port_valid; // @[KCU1500.scala 44:26:@57778.4]
  assign FringeZynq_io_argOuts_18_bits = accel_io_argOuts_18_port_bits; // @[KCU1500.scala 43:25:@57777.4]
  assign FringeZynq_io_argOuts_19_valid = accel_io_argOuts_19_port_valid; // @[KCU1500.scala 44:26:@57780.4]
  assign FringeZynq_io_argOuts_19_bits = accel_io_argOuts_19_port_bits; // @[KCU1500.scala 43:25:@57779.4]
  assign FringeZynq_io_argOuts_20_valid = accel_io_argOuts_20_port_valid; // @[KCU1500.scala 44:26:@57782.4]
  assign FringeZynq_io_argOuts_20_bits = accel_io_argOuts_20_port_bits; // @[KCU1500.scala 43:25:@57781.4]
  assign FringeZynq_io_argOuts_21_valid = accel_io_argOuts_21_port_valid; // @[KCU1500.scala 44:26:@57784.4]
  assign FringeZynq_io_argOuts_21_bits = accel_io_argOuts_21_port_bits; // @[KCU1500.scala 43:25:@57783.4]
  assign FringeZynq_io_argOuts_22_valid = accel_io_argOuts_22_port_valid; // @[KCU1500.scala 44:26:@57786.4]
  assign FringeZynq_io_argOuts_22_bits = accel_io_argOuts_22_port_bits; // @[KCU1500.scala 43:25:@57785.4]
  assign FringeZynq_io_argOuts_23_valid = accel_io_argOuts_23_port_valid; // @[KCU1500.scala 44:26:@57788.4]
  assign FringeZynq_io_argOuts_23_bits = accel_io_argOuts_23_port_bits; // @[KCU1500.scala 43:25:@57787.4]
  assign FringeZynq_io_argOuts_24_valid = accel_io_argOuts_24_port_valid; // @[KCU1500.scala 44:26:@57790.4]
  assign FringeZynq_io_argOuts_24_bits = accel_io_argOuts_24_port_bits; // @[KCU1500.scala 43:25:@57789.4]
  assign FringeZynq_io_argOuts_25_valid = accel_io_argOuts_25_port_valid; // @[KCU1500.scala 44:26:@57792.4]
  assign FringeZynq_io_argOuts_25_bits = accel_io_argOuts_25_port_bits; // @[KCU1500.scala 43:25:@57791.4]
  assign FringeZynq_io_argOuts_26_valid = accel_io_argOuts_26_port_valid; // @[KCU1500.scala 44:26:@57794.4]
  assign FringeZynq_io_argOuts_26_bits = accel_io_argOuts_26_port_bits; // @[KCU1500.scala 43:25:@57793.4]
  assign FringeZynq_io_argOuts_27_valid = accel_io_argOuts_27_port_valid; // @[KCU1500.scala 44:26:@57796.4]
  assign FringeZynq_io_argOuts_27_bits = accel_io_argOuts_27_port_bits; // @[KCU1500.scala 43:25:@57795.4]
  assign FringeZynq_io_argOuts_28_valid = accel_io_argOuts_28_port_valid; // @[KCU1500.scala 44:26:@57798.4]
  assign FringeZynq_io_argOuts_28_bits = accel_io_argOuts_28_port_bits; // @[KCU1500.scala 43:25:@57797.4]
  assign FringeZynq_io_argOuts_29_valid = accel_io_argOuts_29_port_valid; // @[KCU1500.scala 44:26:@57800.4]
  assign FringeZynq_io_argOuts_29_bits = accel_io_argOuts_29_port_bits; // @[KCU1500.scala 43:25:@57799.4]
  assign FringeZynq_io_argOuts_30_valid = accel_io_argOuts_30_port_valid; // @[KCU1500.scala 44:26:@57802.4]
  assign FringeZynq_io_argOuts_30_bits = accel_io_argOuts_30_port_bits; // @[KCU1500.scala 43:25:@57801.4]
  assign FringeZynq_io_argOuts_31_valid = accel_io_argOuts_31_port_valid; // @[KCU1500.scala 44:26:@57804.4]
  assign FringeZynq_io_argOuts_31_bits = accel_io_argOuts_31_port_bits; // @[KCU1500.scala 43:25:@57803.4]
  assign FringeZynq_io_heap_0_req_valid = accel_io_heap_0_req_valid; // @[KCU1500.scala 57:20:@57964.4]
  assign FringeZynq_io_heap_0_req_bits_allocDealloc = accel_io_heap_0_req_bits_allocDealloc; // @[KCU1500.scala 57:20:@57963.4]
  assign FringeZynq_io_heap_0_req_bits_sizeAddr = accel_io_heap_0_req_bits_sizeAddr; // @[KCU1500.scala 57:20:@57962.4]
endmodule
module SRAMVerilogAWS
#(
    parameter WORDS = 1024,
    parameter AWIDTH = 10,
    parameter DWIDTH = 32)
(
    input clk,
    input [AWIDTH-1:0] raddr,
    input [AWIDTH-1:0] waddr,
    input raddrEn,
    input waddrEn,
    input wen,
    input [DWIDTH-1:0] wdata,
    input backpressure,
    output reg [DWIDTH-1:0] rdata
);

    reg [DWIDTH-1:0] mem [0:WORDS-1];

    always @(posedge clk) begin
      if (wen) mem[waddr] <= wdata;
      if (backpressure) rdata <= mem[raddr];
    end

endmodule
