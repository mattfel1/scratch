module FF( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  output [31:0] io_rPort_0_output_0, // @[:@6.4]
  input  [31:0] io_wPort_0_data_0, // @[:@6.4]
  input         io_wPort_0_reset, // @[:@6.4]
  input         io_wPort_0_en_0 // @[:@6.4]
);
  reg [31:0] ff; // @[MemPrimitives.scala 173:19:@21.4]
  reg [31:0] _RAND_0;
  wire [31:0] _T_68; // @[MemPrimitives.scala 177:32:@23.4]
  wire [31:0] _T_69; // @[MemPrimitives.scala 177:12:@24.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 177:32:@23.4]
  assign _T_69 = io_wPort_0_reset ? 32'h0 : _T_68; // @[MemPrimitives.scala 177:12:@24.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 178:34:@26.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 32'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 32'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SRFF( // @[:@28.2]
  input   clock, // @[:@29.4]
  input   reset, // @[:@30.4]
  input   io_input_set, // @[:@31.4]
  input   io_input_reset, // @[:@31.4]
  input   io_input_asyn_reset, // @[:@31.4]
  output  io_output // @[:@31.4]
);
  reg  _T_15; // @[SRFF.scala 20:21:@33.4]
  reg [31:0] _RAND_0;
  wire  _T_19; // @[SRFF.scala 21:74:@34.4]
  wire  _T_20; // @[SRFF.scala 21:48:@35.4]
  wire  _T_21; // @[SRFF.scala 21:14:@36.4]
  assign _T_19 = io_input_reset ? 1'h0 : _T_15; // @[SRFF.scala 21:74:@34.4]
  assign _T_20 = io_input_set ? 1'h1 : _T_19; // @[SRFF.scala 21:48:@35.4]
  assign _T_21 = io_input_asyn_reset ? 1'h0 : _T_20; // @[SRFF.scala 21:14:@36.4]
  assign io_output = io_input_asyn_reset ? 1'h0 : _T_15; // @[SRFF.scala 22:15:@39.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_15 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_15 <= 1'h0;
    end else begin
      if (io_input_asyn_reset) begin
        _T_15 <= 1'h0;
      end else begin
        if (io_input_set) begin
          _T_15 <= 1'h1;
        end else begin
          if (io_input_reset) begin
            _T_15 <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module SingleCounter( // @[:@41.2]
  input   clock, // @[:@42.4]
  input   reset, // @[:@43.4]
  input   io_input_reset, // @[:@44.4]
  output  io_output_done // @[:@44.4]
);
  wire  bases_0_clock; // @[Counter.scala 253:53:@57.4]
  wire  bases_0_reset; // @[Counter.scala 253:53:@57.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 253:53:@57.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 253:53:@57.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 253:53:@57.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 253:53:@57.4]
  wire  SRFF_clock; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_reset; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_input_set; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_output; // @[Counter.scala 255:22:@73.4]
  wire [31:0] _T_48; // @[Counter.scala 279:52:@101.4]
  wire [32:0] _T_50; // @[Counter.scala 283:33:@102.4]
  wire [31:0] _T_51; // @[Counter.scala 283:33:@103.4]
  wire [31:0] _T_52; // @[Counter.scala 283:33:@104.4]
  wire  _T_57; // @[Counter.scala 285:18:@106.4]
  wire [31:0] _T_68; // @[Counter.scala 291:115:@114.4]
  wire [31:0] _T_71; // @[Counter.scala 291:152:@117.4]
  wire [31:0] _T_72; // @[Counter.scala 291:74:@118.4]
  FF bases_0 ( // @[Counter.scala 253:53:@57.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 255:22:@73.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 279:52:@101.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@102.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@103.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 283:33:@104.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh3); // @[Counter.scala 285:18:@106.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 291:115:@114.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 291:152:@117.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 291:74:@118.4]
  assign io_output_done = $signed(_T_52) >= $signed(32'sh3); // @[Counter.scala 325:20:@127.4]
  assign bases_0_clock = clock; // @[:@58.4]
  assign bases_0_reset = reset; // @[:@59.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 291:31:@120.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 273:27:@99.4]
  assign bases_0_io_wPort_0_en_0 = 1'h1; // @[Counter.scala 276:29:@100.4]
  assign SRFF_clock = clock; // @[:@74.4]
  assign SRFF_reset = reset; // @[:@75.4]
  assign SRFF_io_input_set = io_input_reset == 1'h0; // @[Counter.scala 256:23:@78.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 257:25:@80.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 258:30:@81.4]
endmodule
module RetimeWrapper( // @[:@144.2]
  input   clock, // @[:@145.4]
  input   reset, // @[:@146.4]
  input   io_flow, // @[:@147.4]
  input   io_in, // @[:@147.4]
  output  io_out // @[:@147.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@149.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@149.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@162.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@161.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@160.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@159.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@158.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@156.4]
endmodule
module RootController_sm( // @[:@312.2]
  input   clock, // @[:@313.4]
  input   reset, // @[:@314.4]
  input   io_enable, // @[:@315.4]
  output  io_done, // @[:@315.4]
  input   io_rst, // @[:@315.4]
  input   io_ctrDone, // @[:@315.4]
  output  io_ctrInc, // @[:@315.4]
  input   io_doneIn_0, // @[:@315.4]
  output  io_enableOut_0, // @[:@315.4]
  output  io_childAck_0 // @[:@315.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@318.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@321.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@338.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@433.4]
  wire  finished; // @[Controllers.scala 81:26:@324.4]
  wire  synchronize; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  wire  _T_122; // @[Controllers.scala 128:33:@371.4]
  wire  _T_124; // @[Controllers.scala 128:54:@372.4]
  wire  _T_125; // @[Controllers.scala 128:52:@373.4]
  wire  _T_126; // @[Controllers.scala 128:66:@374.4]
  wire  _T_128; // @[Controllers.scala 128:98:@376.4]
  wire  _T_129; // @[Controllers.scala 128:96:@377.4]
  wire  _T_131; // @[Controllers.scala 128:123:@378.4]
  wire  _T_133; // @[Controllers.scala 129:48:@381.4]
  wire  _T_138; // @[Controllers.scala 130:52:@386.4]
  wire  _T_139; // @[Controllers.scala 130:50:@387.4]
  wire  _T_147; // @[Controllers.scala 130:129:@393.4]
  wire  _T_150; // @[Controllers.scala 131:45:@396.4]
  wire  _T_154; // @[Controllers.scala 213:68:@402.4]
  wire  _T_156; // @[Controllers.scala 213:90:@404.4]
  wire  _T_158; // @[Controllers.scala 213:132:@406.4]
  wire  _T_159; // @[Controllers.scala 213:130:@407.4]
  wire  _T_160; // @[Controllers.scala 213:156:@408.4]
  reg  _T_166; // @[package.scala 48:56:@412.4]
  reg [31:0] _RAND_0;
  reg  _T_180; // @[package.scala 48:56:@430.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@318.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@321.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@338.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@357.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@416.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@433.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  assign finished = done_0_io_output | io_done; // @[Controllers.scala 81:26:@324.4]
  assign synchronize = RetimeWrapper_io_out; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  assign _T_122 = done_0_io_output == 1'h0; // @[Controllers.scala 128:33:@371.4]
  assign _T_124 = io_ctrDone == 1'h0; // @[Controllers.scala 128:54:@372.4]
  assign _T_125 = _T_122 & _T_124; // @[Controllers.scala 128:52:@373.4]
  assign _T_126 = _T_125 & io_enable; // @[Controllers.scala 128:66:@374.4]
  assign _T_128 = ~ iterDone_0_io_output; // @[Controllers.scala 128:98:@376.4]
  assign _T_129 = _T_126 & _T_128; // @[Controllers.scala 128:96:@377.4]
  assign _T_131 = io_doneIn_0 == 1'h0; // @[Controllers.scala 128:123:@378.4]
  assign _T_133 = io_doneIn_0 | io_rst; // @[Controllers.scala 129:48:@381.4]
  assign _T_138 = synchronize == 1'h0; // @[Controllers.scala 130:52:@386.4]
  assign _T_139 = io_doneIn_0 & _T_138; // @[Controllers.scala 130:50:@387.4]
  assign _T_147 = finished == 1'h0; // @[Controllers.scala 130:129:@393.4]
  assign _T_150 = io_rst == 1'h0; // @[Controllers.scala 131:45:@396.4]
  assign _T_154 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@402.4]
  assign _T_156 = _T_154 & _T_128; // @[Controllers.scala 213:90:@404.4]
  assign _T_158 = ~ done_0_io_output; // @[Controllers.scala 213:132:@406.4]
  assign _T_159 = _T_156 & _T_158; // @[Controllers.scala 213:130:@407.4]
  assign _T_160 = ~ io_ctrDone; // @[Controllers.scala 213:156:@408.4]
  assign io_done = RetimeWrapper_2_io_out; // @[Controllers.scala 245:13:@440.4]
  assign io_ctrInc = io_doneIn_0; // @[Controllers.scala 122:17:@356.4]
  assign io_enableOut_0 = _T_159 & _T_160; // @[Controllers.scala 213:55:@410.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@401.4]
  assign active_0_clock = clock; // @[:@319.4]
  assign active_0_reset = reset; // @[:@320.4]
  assign active_0_io_input_set = _T_129 & _T_131; // @[Controllers.scala 128:30:@380.4]
  assign active_0_io_input_reset = _T_133 | done_0_io_output; // @[Controllers.scala 129:32:@385.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@326.4]
  assign done_0_clock = clock; // @[:@322.4]
  assign done_0_reset = reset; // @[:@323.4]
  assign done_0_io_input_set = io_ctrDone & _T_150; // @[Controllers.scala 131:28:@399.4]
  assign done_0_io_input_reset = io_rst | done_0_io_output; // @[Controllers.scala 86:33:@336.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@327.4]
  assign iterDone_0_clock = clock; // @[:@339.4]
  assign iterDone_0_reset = reset; // @[:@340.4]
  assign iterDone_0_io_input_set = _T_139 & _T_147; // @[Controllers.scala 130:32:@395.4]
  assign iterDone_0_io_input_reset = synchronize | io_rst; // @[Controllers.scala 92:37:@350.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@341.4]
  assign RetimeWrapper_clock = clock; // @[:@358.4]
  assign RetimeWrapper_reset = reset; // @[:@359.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@361.4]
  assign RetimeWrapper_io_in = io_doneIn_0; // @[package.scala 94:16:@360.4]
  assign RetimeWrapper_1_clock = clock; // @[:@417.4]
  assign RetimeWrapper_1_reset = reset; // @[:@418.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@420.4]
  assign RetimeWrapper_1_io_in = done_0_io_output & _T_166; // @[package.scala 94:16:@419.4]
  assign RetimeWrapper_2_clock = clock; // @[:@434.4]
  assign RetimeWrapper_2_reset = reset; // @[:@435.4]
  assign RetimeWrapper_2_io_flow = io_enable; // @[package.scala 95:18:@437.4]
  assign RetimeWrapper_2_io_in = done_0_io_output & _T_180; // @[package.scala 94:16:@436.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_166 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_180 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_166 <= 1'h0;
    end else begin
      _T_166 <= _T_122;
    end
    if (reset) begin
      _T_180 <= 1'h0;
    end else begin
      _T_180 <= _T_122;
    end
  end
endmodule
module InstrumentationCounter( // @[:@490.2]
  input         clock, // @[:@491.4]
  input         reset, // @[:@492.4]
  input         io_enable, // @[:@493.4]
  output [63:0] io_count // @[:@493.4]
);
  reg [63:0] ff; // @[Counter.scala 214:19:@495.4]
  reg [63:0] _RAND_0;
  wire [64:0] _T_12; // @[Counter.scala 215:27:@496.4]
  wire [63:0] _T_13; // @[Counter.scala 215:27:@497.4]
  wire [63:0] _T_14; // @[Counter.scala 215:12:@498.4]
  assign _T_12 = ff + 64'h1; // @[Counter.scala 215:27:@496.4]
  assign _T_13 = ff + 64'h1; // @[Counter.scala 215:27:@497.4]
  assign _T_14 = io_enable ? _T_13 : ff; // @[Counter.scala 215:12:@498.4]
  assign io_count = ff; // @[Counter.scala 216:12:@500.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  ff = _RAND_0[63:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 64'h0;
    end else begin
      if (io_enable) begin
        ff <= _T_13;
      end
    end
  end
endmodule
module x132_outr_UnitPipe_sm( // @[:@983.2]
  input   clock, // @[:@984.4]
  input   reset, // @[:@985.4]
  input   io_enable, // @[:@986.4]
  output  io_done, // @[:@986.4]
  input   io_parentAck, // @[:@986.4]
  input   io_doneIn_0, // @[:@986.4]
  input   io_doneIn_1, // @[:@986.4]
  input   io_doneIn_2, // @[:@986.4]
  output  io_enableOut_0, // @[:@986.4]
  output  io_enableOut_1, // @[:@986.4]
  output  io_enableOut_2, // @[:@986.4]
  output  io_childAck_0, // @[:@986.4]
  output  io_childAck_1, // @[:@986.4]
  output  io_childAck_2, // @[:@986.4]
  input   io_ctrCopyDone_0, // @[:@986.4]
  input   io_ctrCopyDone_1, // @[:@986.4]
  input   io_ctrCopyDone_2 // @[:@986.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@989.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@989.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@989.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@989.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@989.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@989.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@992.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@992.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@992.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@992.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@992.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@992.4]
  wire  active_2_clock; // @[Controllers.scala 76:50:@995.4]
  wire  active_2_reset; // @[Controllers.scala 76:50:@995.4]
  wire  active_2_io_input_set; // @[Controllers.scala 76:50:@995.4]
  wire  active_2_io_input_reset; // @[Controllers.scala 76:50:@995.4]
  wire  active_2_io_input_asyn_reset; // @[Controllers.scala 76:50:@995.4]
  wire  active_2_io_output; // @[Controllers.scala 76:50:@995.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@998.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@998.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@998.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@998.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@998.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@998.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@1001.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@1001.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@1001.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@1001.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@1001.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@1001.4]
  wire  done_2_clock; // @[Controllers.scala 77:48:@1004.4]
  wire  done_2_reset; // @[Controllers.scala 77:48:@1004.4]
  wire  done_2_io_input_set; // @[Controllers.scala 77:48:@1004.4]
  wire  done_2_io_input_reset; // @[Controllers.scala 77:48:@1004.4]
  wire  done_2_io_input_asyn_reset; // @[Controllers.scala 77:48:@1004.4]
  wire  done_2_io_output; // @[Controllers.scala 77:48:@1004.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@1045.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@1045.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@1045.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@1045.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@1045.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@1045.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@1048.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@1048.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@1048.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@1048.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@1048.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@1048.4]
  wire  iterDone_2_clock; // @[Controllers.scala 90:52:@1051.4]
  wire  iterDone_2_reset; // @[Controllers.scala 90:52:@1051.4]
  wire  iterDone_2_io_input_set; // @[Controllers.scala 90:52:@1051.4]
  wire  iterDone_2_io_input_reset; // @[Controllers.scala 90:52:@1051.4]
  wire  iterDone_2_io_input_asyn_reset; // @[Controllers.scala 90:52:@1051.4]
  wire  iterDone_2_io_output; // @[Controllers.scala 90:52:@1051.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@1102.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@1102.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@1102.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@1102.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@1102.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@1116.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@1116.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@1116.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@1116.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@1116.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@1134.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@1134.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@1134.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@1134.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@1134.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@1171.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@1171.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@1171.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@1171.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@1171.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@1185.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@1185.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@1185.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@1185.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@1185.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@1203.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@1203.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@1203.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@1203.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@1203.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@1240.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@1240.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@1240.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@1240.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@1240.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@1254.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@1254.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@1254.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@1254.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@1254.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@1272.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@1272.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@1272.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@1272.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@1272.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@1329.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@1329.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@1329.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@1329.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@1329.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@1346.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@1346.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@1346.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@1346.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@1346.4]
  wire  _T_77; // @[Controllers.scala 80:47:@1007.4]
  wire  allDone; // @[Controllers.scala 80:47:@1008.4]
  wire  _T_151; // @[Controllers.scala 165:35:@1086.4]
  wire  _T_153; // @[Controllers.scala 165:60:@1087.4]
  wire  _T_154; // @[Controllers.scala 165:58:@1088.4]
  wire  _T_156; // @[Controllers.scala 165:76:@1089.4]
  wire  _T_157; // @[Controllers.scala 165:74:@1090.4]
  wire  _T_161; // @[Controllers.scala 165:109:@1093.4]
  wire  _T_164; // @[Controllers.scala 165:141:@1095.4]
  wire  _T_172; // @[package.scala 96:25:@1107.4 package.scala 96:25:@1108.4]
  wire  _T_176; // @[Controllers.scala 167:54:@1110.4]
  wire  _T_177; // @[Controllers.scala 167:52:@1111.4]
  wire  _T_184; // @[package.scala 96:25:@1121.4 package.scala 96:25:@1122.4]
  wire  _T_202; // @[package.scala 96:25:@1139.4 package.scala 96:25:@1140.4]
  wire  _T_206; // @[Controllers.scala 169:67:@1142.4]
  wire  _T_207; // @[Controllers.scala 169:86:@1143.4]
  wire  _T_219; // @[Controllers.scala 165:35:@1155.4]
  wire  _T_221; // @[Controllers.scala 165:60:@1156.4]
  wire  _T_222; // @[Controllers.scala 165:58:@1157.4]
  wire  _T_224; // @[Controllers.scala 165:76:@1158.4]
  wire  _T_225; // @[Controllers.scala 165:74:@1159.4]
  wire  _T_229; // @[Controllers.scala 165:109:@1162.4]
  wire  _T_232; // @[Controllers.scala 165:141:@1164.4]
  wire  _T_240; // @[package.scala 96:25:@1176.4 package.scala 96:25:@1177.4]
  wire  _T_244; // @[Controllers.scala 167:54:@1179.4]
  wire  _T_245; // @[Controllers.scala 167:52:@1180.4]
  wire  _T_252; // @[package.scala 96:25:@1190.4 package.scala 96:25:@1191.4]
  wire  _T_270; // @[package.scala 96:25:@1208.4 package.scala 96:25:@1209.4]
  wire  _T_274; // @[Controllers.scala 169:67:@1211.4]
  wire  _T_275; // @[Controllers.scala 169:86:@1212.4]
  wire  _T_287; // @[Controllers.scala 165:35:@1224.4]
  wire  _T_289; // @[Controllers.scala 165:60:@1225.4]
  wire  _T_290; // @[Controllers.scala 165:58:@1226.4]
  wire  _T_292; // @[Controllers.scala 165:76:@1227.4]
  wire  _T_293; // @[Controllers.scala 165:74:@1228.4]
  wire  _T_297; // @[Controllers.scala 165:109:@1231.4]
  wire  _T_300; // @[Controllers.scala 165:141:@1233.4]
  wire  _T_308; // @[package.scala 96:25:@1245.4 package.scala 96:25:@1246.4]
  wire  _T_312; // @[Controllers.scala 167:54:@1248.4]
  wire  _T_313; // @[Controllers.scala 167:52:@1249.4]
  wire  _T_320; // @[package.scala 96:25:@1259.4 package.scala 96:25:@1260.4]
  wire  _T_338; // @[package.scala 96:25:@1277.4 package.scala 96:25:@1278.4]
  wire  _T_342; // @[Controllers.scala 169:67:@1280.4]
  wire  _T_343; // @[Controllers.scala 169:86:@1281.4]
  wire  _T_358; // @[Controllers.scala 213:68:@1299.4]
  wire  _T_360; // @[Controllers.scala 213:90:@1301.4]
  wire  _T_362; // @[Controllers.scala 213:132:@1303.4]
  wire  _T_366; // @[Controllers.scala 213:68:@1308.4]
  wire  _T_368; // @[Controllers.scala 213:90:@1310.4]
  wire  _T_374; // @[Controllers.scala 213:68:@1316.4]
  wire  _T_376; // @[Controllers.scala 213:90:@1318.4]
  wire  _T_383; // @[package.scala 100:49:@1324.4]
  reg  _T_386; // @[package.scala 48:56:@1325.4]
  reg [31:0] _RAND_0;
  wire  _T_387; // @[package.scala 100:41:@1327.4]
  reg  _T_400; // @[package.scala 48:56:@1343.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@989.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@992.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF active_2 ( // @[Controllers.scala 76:50:@995.4]
    .clock(active_2_clock),
    .reset(active_2_reset),
    .io_input_set(active_2_io_input_set),
    .io_input_reset(active_2_io_input_reset),
    .io_input_asyn_reset(active_2_io_input_asyn_reset),
    .io_output(active_2_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@998.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@1001.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF done_2 ( // @[Controllers.scala 77:48:@1004.4]
    .clock(done_2_clock),
    .reset(done_2_reset),
    .io_input_set(done_2_io_input_set),
    .io_input_reset(done_2_io_input_reset),
    .io_input_asyn_reset(done_2_io_input_asyn_reset),
    .io_output(done_2_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@1045.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@1048.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  SRFF iterDone_2 ( // @[Controllers.scala 90:52:@1051.4]
    .clock(iterDone_2_clock),
    .reset(iterDone_2_reset),
    .io_input_set(iterDone_2_io_input_set),
    .io_input_reset(iterDone_2_io_input_reset),
    .io_input_asyn_reset(iterDone_2_io_input_asyn_reset),
    .io_output(iterDone_2_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@1102.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@1116.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@1134.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@1171.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@1185.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@1203.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@1240.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@1254.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper RetimeWrapper_8 ( // @[package.scala 93:22:@1272.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper RetimeWrapper_9 ( // @[package.scala 93:22:@1329.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper RetimeWrapper_10 ( // @[package.scala 93:22:@1346.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  assign _T_77 = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@1007.4]
  assign allDone = _T_77 & done_2_io_output; // @[Controllers.scala 80:47:@1008.4]
  assign _T_151 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@1086.4]
  assign _T_153 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@1087.4]
  assign _T_154 = _T_151 & _T_153; // @[Controllers.scala 165:58:@1088.4]
  assign _T_156 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@1089.4]
  assign _T_157 = _T_154 & _T_156; // @[Controllers.scala 165:74:@1090.4]
  assign _T_161 = _T_157 & io_enable; // @[Controllers.scala 165:109:@1093.4]
  assign _T_164 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@1095.4]
  assign _T_172 = RetimeWrapper_io_out; // @[package.scala 96:25:@1107.4 package.scala 96:25:@1108.4]
  assign _T_176 = _T_172 == 1'h0; // @[Controllers.scala 167:54:@1110.4]
  assign _T_177 = io_doneIn_0 | _T_176; // @[Controllers.scala 167:52:@1111.4]
  assign _T_184 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@1121.4 package.scala 96:25:@1122.4]
  assign _T_202 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@1139.4 package.scala 96:25:@1140.4]
  assign _T_206 = _T_202 == 1'h0; // @[Controllers.scala 169:67:@1142.4]
  assign _T_207 = _T_206 & io_enable; // @[Controllers.scala 169:86:@1143.4]
  assign _T_219 = ~ iterDone_1_io_output; // @[Controllers.scala 165:35:@1155.4]
  assign _T_221 = io_doneIn_1 == 1'h0; // @[Controllers.scala 165:60:@1156.4]
  assign _T_222 = _T_219 & _T_221; // @[Controllers.scala 165:58:@1157.4]
  assign _T_224 = done_1_io_output == 1'h0; // @[Controllers.scala 165:76:@1158.4]
  assign _T_225 = _T_222 & _T_224; // @[Controllers.scala 165:74:@1159.4]
  assign _T_229 = _T_225 & io_enable; // @[Controllers.scala 165:109:@1162.4]
  assign _T_232 = io_ctrCopyDone_1 == 1'h0; // @[Controllers.scala 165:141:@1164.4]
  assign _T_240 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@1176.4 package.scala 96:25:@1177.4]
  assign _T_244 = _T_240 == 1'h0; // @[Controllers.scala 167:54:@1179.4]
  assign _T_245 = io_doneIn_1 | _T_244; // @[Controllers.scala 167:52:@1180.4]
  assign _T_252 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@1190.4 package.scala 96:25:@1191.4]
  assign _T_270 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@1208.4 package.scala 96:25:@1209.4]
  assign _T_274 = _T_270 == 1'h0; // @[Controllers.scala 169:67:@1211.4]
  assign _T_275 = _T_274 & io_enable; // @[Controllers.scala 169:86:@1212.4]
  assign _T_287 = ~ iterDone_2_io_output; // @[Controllers.scala 165:35:@1224.4]
  assign _T_289 = io_doneIn_2 == 1'h0; // @[Controllers.scala 165:60:@1225.4]
  assign _T_290 = _T_287 & _T_289; // @[Controllers.scala 165:58:@1226.4]
  assign _T_292 = done_2_io_output == 1'h0; // @[Controllers.scala 165:76:@1227.4]
  assign _T_293 = _T_290 & _T_292; // @[Controllers.scala 165:74:@1228.4]
  assign _T_297 = _T_293 & io_enable; // @[Controllers.scala 165:109:@1231.4]
  assign _T_300 = io_ctrCopyDone_2 == 1'h0; // @[Controllers.scala 165:141:@1233.4]
  assign _T_308 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@1245.4 package.scala 96:25:@1246.4]
  assign _T_312 = _T_308 == 1'h0; // @[Controllers.scala 167:54:@1248.4]
  assign _T_313 = io_doneIn_2 | _T_312; // @[Controllers.scala 167:52:@1249.4]
  assign _T_320 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@1259.4 package.scala 96:25:@1260.4]
  assign _T_338 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@1277.4 package.scala 96:25:@1278.4]
  assign _T_342 = _T_338 == 1'h0; // @[Controllers.scala 169:67:@1280.4]
  assign _T_343 = _T_342 & io_enable; // @[Controllers.scala 169:86:@1281.4]
  assign _T_358 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@1299.4]
  assign _T_360 = _T_358 & _T_151; // @[Controllers.scala 213:90:@1301.4]
  assign _T_362 = ~ allDone; // @[Controllers.scala 213:132:@1303.4]
  assign _T_366 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@1308.4]
  assign _T_368 = _T_366 & _T_219; // @[Controllers.scala 213:90:@1310.4]
  assign _T_374 = io_enable & active_2_io_output; // @[Controllers.scala 213:68:@1316.4]
  assign _T_376 = _T_374 & _T_287; // @[Controllers.scala 213:90:@1318.4]
  assign _T_383 = allDone == 1'h0; // @[package.scala 100:49:@1324.4]
  assign _T_387 = allDone & _T_386; // @[package.scala 100:41:@1327.4]
  assign io_done = RetimeWrapper_10_io_out; // @[Controllers.scala 245:13:@1353.4]
  assign io_enableOut_0 = _T_360 & _T_362; // @[Controllers.scala 213:55:@1307.4]
  assign io_enableOut_1 = _T_368 & _T_362; // @[Controllers.scala 213:55:@1315.4]
  assign io_enableOut_2 = _T_376 & _T_362; // @[Controllers.scala 213:55:@1323.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@1294.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@1296.4]
  assign io_childAck_2 = iterDone_2_io_output; // @[Controllers.scala 212:58:@1298.4]
  assign active_0_clock = clock; // @[:@990.4]
  assign active_0_reset = reset; // @[:@991.4]
  assign active_0_io_input_set = _T_161 & _T_164; // @[Controllers.scala 165:32:@1097.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@1101.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@1011.4]
  assign active_1_clock = clock; // @[:@993.4]
  assign active_1_reset = reset; // @[:@994.4]
  assign active_1_io_input_set = _T_229 & _T_232; // @[Controllers.scala 165:32:@1166.4]
  assign active_1_io_input_reset = io_ctrCopyDone_1 | io_parentAck; // @[Controllers.scala 166:34:@1170.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@1012.4]
  assign active_2_clock = clock; // @[:@996.4]
  assign active_2_reset = reset; // @[:@997.4]
  assign active_2_io_input_set = _T_297 & _T_300; // @[Controllers.scala 165:32:@1235.4]
  assign active_2_io_input_reset = io_ctrCopyDone_2 | io_parentAck; // @[Controllers.scala 166:34:@1239.4]
  assign active_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@1013.4]
  assign done_0_clock = clock; // @[:@999.4]
  assign done_0_reset = reset; // @[:@1000.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_207; // @[Controllers.scala 169:30:@1147.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@1025.4 Controllers.scala 170:32:@1154.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@1014.4]
  assign done_1_clock = clock; // @[:@1002.4]
  assign done_1_reset = reset; // @[:@1003.4]
  assign done_1_io_input_set = io_ctrCopyDone_1 | _T_275; // @[Controllers.scala 169:30:@1216.4]
  assign done_1_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@1034.4 Controllers.scala 170:32:@1223.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@1015.4]
  assign done_2_clock = clock; // @[:@1005.4]
  assign done_2_reset = reset; // @[:@1006.4]
  assign done_2_io_input_set = io_ctrCopyDone_2 | _T_343; // @[Controllers.scala 169:30:@1285.4]
  assign done_2_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@1043.4 Controllers.scala 170:32:@1292.4]
  assign done_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@1016.4]
  assign iterDone_0_clock = clock; // @[:@1046.4]
  assign iterDone_0_reset = reset; // @[:@1047.4]
  assign iterDone_0_io_input_set = _T_177 & io_enable; // @[Controllers.scala 167:34:@1115.4]
  assign iterDone_0_io_input_reset = _T_184 | io_parentAck; // @[Controllers.scala 92:37:@1065.4 Controllers.scala 168:36:@1131.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@1054.4]
  assign iterDone_1_clock = clock; // @[:@1049.4]
  assign iterDone_1_reset = reset; // @[:@1050.4]
  assign iterDone_1_io_input_set = _T_245 & io_enable; // @[Controllers.scala 167:34:@1184.4]
  assign iterDone_1_io_input_reset = _T_252 | io_parentAck; // @[Controllers.scala 92:37:@1074.4 Controllers.scala 168:36:@1200.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@1055.4]
  assign iterDone_2_clock = clock; // @[:@1052.4]
  assign iterDone_2_reset = reset; // @[:@1053.4]
  assign iterDone_2_io_input_set = _T_313 & io_enable; // @[Controllers.scala 167:34:@1253.4]
  assign iterDone_2_io_input_reset = _T_320 | io_parentAck; // @[Controllers.scala 92:37:@1083.4 Controllers.scala 168:36:@1269.4]
  assign iterDone_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@1056.4]
  assign RetimeWrapper_clock = clock; // @[:@1103.4]
  assign RetimeWrapper_reset = reset; // @[:@1104.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@1106.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@1105.4]
  assign RetimeWrapper_1_clock = clock; // @[:@1117.4]
  assign RetimeWrapper_1_reset = reset; // @[:@1118.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@1120.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@1119.4]
  assign RetimeWrapper_2_clock = clock; // @[:@1135.4]
  assign RetimeWrapper_2_reset = reset; // @[:@1136.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@1138.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@1137.4]
  assign RetimeWrapper_3_clock = clock; // @[:@1172.4]
  assign RetimeWrapper_3_reset = reset; // @[:@1173.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@1175.4]
  assign RetimeWrapper_3_io_in = 1'h1; // @[package.scala 94:16:@1174.4]
  assign RetimeWrapper_4_clock = clock; // @[:@1186.4]
  assign RetimeWrapper_4_reset = reset; // @[:@1187.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@1189.4]
  assign RetimeWrapper_4_io_in = io_doneIn_1; // @[package.scala 94:16:@1188.4]
  assign RetimeWrapper_5_clock = clock; // @[:@1204.4]
  assign RetimeWrapper_5_reset = reset; // @[:@1205.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@1207.4]
  assign RetimeWrapper_5_io_in = 1'h1; // @[package.scala 94:16:@1206.4]
  assign RetimeWrapper_6_clock = clock; // @[:@1241.4]
  assign RetimeWrapper_6_reset = reset; // @[:@1242.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@1244.4]
  assign RetimeWrapper_6_io_in = 1'h1; // @[package.scala 94:16:@1243.4]
  assign RetimeWrapper_7_clock = clock; // @[:@1255.4]
  assign RetimeWrapper_7_reset = reset; // @[:@1256.4]
  assign RetimeWrapper_7_io_flow = 1'h1; // @[package.scala 95:18:@1258.4]
  assign RetimeWrapper_7_io_in = io_doneIn_2; // @[package.scala 94:16:@1257.4]
  assign RetimeWrapper_8_clock = clock; // @[:@1273.4]
  assign RetimeWrapper_8_reset = reset; // @[:@1274.4]
  assign RetimeWrapper_8_io_flow = 1'h1; // @[package.scala 95:18:@1276.4]
  assign RetimeWrapper_8_io_in = 1'h1; // @[package.scala 94:16:@1275.4]
  assign RetimeWrapper_9_clock = clock; // @[:@1330.4]
  assign RetimeWrapper_9_reset = reset; // @[:@1331.4]
  assign RetimeWrapper_9_io_flow = 1'h1; // @[package.scala 95:18:@1333.4]
  assign RetimeWrapper_9_io_in = _T_387 | io_parentAck; // @[package.scala 94:16:@1332.4]
  assign RetimeWrapper_10_clock = clock; // @[:@1347.4]
  assign RetimeWrapper_10_reset = reset; // @[:@1348.4]
  assign RetimeWrapper_10_io_flow = io_enable; // @[package.scala 95:18:@1350.4]
  assign RetimeWrapper_10_io_in = allDone & _T_400; // @[package.scala 94:16:@1349.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_386 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_400 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_386 <= 1'h0;
    end else begin
      _T_386 <= _T_383;
    end
    if (reset) begin
      _T_400 <= 1'h0;
    end else begin
      _T_400 <= _T_383;
    end
  end
endmodule
module FF_1( // @[:@1459.2]
  input        clock, // @[:@1460.4]
  input        reset, // @[:@1461.4]
  output [5:0] io_rPort_0_output_0, // @[:@1462.4]
  input  [5:0] io_wPort_0_data_0, // @[:@1462.4]
  input        io_wPort_0_reset, // @[:@1462.4]
  input  [5:0] io_wPort_0_init, // @[:@1462.4]
  input        io_wPort_0_en_0, // @[:@1462.4]
  input        io_reset // @[:@1462.4]
);
  reg [5:0] ff; // @[MemPrimitives.scala 173:19:@1477.4]
  reg [31:0] _RAND_0;
  wire  anyReset; // @[MemPrimitives.scala 174:65:@1478.4]
  wire [5:0] _T_68; // @[MemPrimitives.scala 177:32:@1479.4]
  wire [5:0] _T_69; // @[MemPrimitives.scala 177:12:@1480.4]
  assign anyReset = io_wPort_0_reset | io_reset; // @[MemPrimitives.scala 174:65:@1478.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 177:32:@1479.4]
  assign _T_69 = anyReset ? io_wPort_0_init : _T_68; // @[MemPrimitives.scala 177:12:@1480.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 178:34:@1482.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[5:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= io_wPort_0_init;
    end else begin
      if (anyReset) begin
        ff <= io_wPort_0_init;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module CompactingCounter( // @[:@1484.2]
  input        clock, // @[:@1485.4]
  input        reset, // @[:@1486.4]
  input        io_input_dir, // @[:@1487.4]
  input        io_input_reset, // @[:@1487.4]
  input        io_input_enables_0, // @[:@1487.4]
  output [5:0] io_output_count // @[:@1487.4]
);
  wire  base_clock; // @[Counter.scala 191:20:@1489.4]
  wire  base_reset; // @[Counter.scala 191:20:@1489.4]
  wire [5:0] base_io_rPort_0_output_0; // @[Counter.scala 191:20:@1489.4]
  wire [5:0] base_io_wPort_0_data_0; // @[Counter.scala 191:20:@1489.4]
  wire  base_io_wPort_0_reset; // @[Counter.scala 191:20:@1489.4]
  wire [5:0] base_io_wPort_0_init; // @[Counter.scala 191:20:@1489.4]
  wire  base_io_wPort_0_en_0; // @[Counter.scala 191:20:@1489.4]
  wire  base_io_reset; // @[Counter.scala 191:20:@1489.4]
  wire [5:0] count; // @[Counter.scala 197:42:@1508.4]
  wire [5:0] num_enabled; // @[Counter.scala 198:56:@1509.4]
  wire [6:0] _T_23; // @[Counter.scala 199:55:@1510.4]
  wire [5:0] _T_24; // @[Counter.scala 199:55:@1511.4]
  wire [5:0] _T_25; // @[Counter.scala 199:55:@1512.4]
  wire [5:0] _T_26; // @[Counter.scala 199:27:@1513.4]
  wire [6:0] _T_27; // @[Counter.scala 199:22:@1514.4]
  wire [5:0] _T_28; // @[Counter.scala 199:22:@1515.4]
  wire [5:0] newval; // @[Counter.scala 199:22:@1516.4]
  wire  _T_30; // @[Counter.scala 200:40:@1517.4]
  wire  _T_32; // @[Counter.scala 200:59:@1518.4]
  wire  isMax; // @[Counter.scala 200:18:@1519.4]
  wire [6:0] _T_34; // @[Counter.scala 201:32:@1520.4]
  wire [5:0] _T_35; // @[Counter.scala 201:32:@1521.4]
  wire [5:0] _T_36; // @[Counter.scala 201:32:@1522.4]
  wire [5:0] next; // @[Counter.scala 201:17:@1523.4]
  wire [5:0] _T_38; // @[Counter.scala 202:68:@1524.4]
  FF_1 base ( // @[Counter.scala 191:20:@1489.4]
    .clock(base_clock),
    .reset(base_reset),
    .io_rPort_0_output_0(base_io_rPort_0_output_0),
    .io_wPort_0_data_0(base_io_wPort_0_data_0),
    .io_wPort_0_reset(base_io_wPort_0_reset),
    .io_wPort_0_init(base_io_wPort_0_init),
    .io_wPort_0_en_0(base_io_wPort_0_en_0),
    .io_reset(base_io_reset)
  );
  assign count = $signed(base_io_rPort_0_output_0); // @[Counter.scala 197:42:@1508.4]
  assign num_enabled = io_input_enables_0 ? $signed(6'sh1) : $signed(6'sh0); // @[Counter.scala 198:56:@1509.4]
  assign _T_23 = $signed(6'sh0) - $signed(num_enabled); // @[Counter.scala 199:55:@1510.4]
  assign _T_24 = $signed(6'sh0) - $signed(num_enabled); // @[Counter.scala 199:55:@1511.4]
  assign _T_25 = $signed(_T_24); // @[Counter.scala 199:55:@1512.4]
  assign _T_26 = io_input_dir ? $signed(num_enabled) : $signed(_T_25); // @[Counter.scala 199:27:@1513.4]
  assign _T_27 = $signed(count) + $signed(_T_26); // @[Counter.scala 199:22:@1514.4]
  assign _T_28 = $signed(count) + $signed(_T_26); // @[Counter.scala 199:22:@1515.4]
  assign newval = $signed(_T_28); // @[Counter.scala 199:22:@1516.4]
  assign _T_30 = $signed(newval) >= $signed(6'sh8); // @[Counter.scala 200:40:@1517.4]
  assign _T_32 = $signed(newval) <= $signed(6'sh0); // @[Counter.scala 200:59:@1518.4]
  assign isMax = io_input_dir ? _T_30 : _T_32; // @[Counter.scala 200:18:@1519.4]
  assign _T_34 = $signed(newval) - $signed(6'sh8); // @[Counter.scala 201:32:@1520.4]
  assign _T_35 = $signed(newval) - $signed(6'sh8); // @[Counter.scala 201:32:@1521.4]
  assign _T_36 = $signed(_T_35); // @[Counter.scala 201:32:@1522.4]
  assign next = isMax ? $signed(_T_36) : $signed(newval); // @[Counter.scala 201:17:@1523.4]
  assign _T_38 = $unsigned(next); // @[Counter.scala 202:68:@1524.4]
  assign io_output_count = $signed(base_io_rPort_0_output_0); // @[Counter.scala 204:19:@1528.4]
  assign base_clock = clock; // @[:@1490.4]
  assign base_reset = reset; // @[:@1491.4]
  assign base_io_wPort_0_data_0 = io_input_reset ? 6'h0 : _T_38; // @[Counter.scala 202:30:@1526.4]
  assign base_io_wPort_0_reset = io_input_reset; // @[Counter.scala 194:26:@1506.4]
  assign base_io_wPort_0_init = 6'h0; // @[Counter.scala 193:25:@1505.4]
  assign base_io_wPort_0_en_0 = io_input_enables_0; // @[Counter.scala 195:28:@1507.4]
  assign base_io_reset = 1'h0;
endmodule
module CompactingIncDincCtr( // @[:@1605.2]
  input   clock, // @[:@1606.4]
  input   reset, // @[:@1607.4]
  input   io_input_inc_en_0, // @[:@1608.4]
  input   io_input_dinc_en_0, // @[:@1608.4]
  output  io_output_empty, // @[:@1608.4]
  output  io_output_full // @[:@1608.4]
);
  reg [31:0] cnt; // @[Counter.scala 162:20:@1610.4]
  reg [31:0] _RAND_0;
  wire [5:0] numPushed; // @[Counter.scala 164:47:@1611.4]
  wire [5:0] numPopped; // @[Counter.scala 165:48:@1612.4]
  wire [31:0] _GEN_0; // @[Counter.scala 166:14:@1613.4]
  wire [32:0] _T_37; // @[Counter.scala 166:14:@1613.4]
  wire [31:0] _T_38; // @[Counter.scala 166:14:@1614.4]
  wire [31:0] _T_39; // @[Counter.scala 166:14:@1615.4]
  wire [31:0] _GEN_1; // @[Counter.scala 166:26:@1616.4]
  wire [32:0] _T_40; // @[Counter.scala 166:26:@1616.4]
  wire [31:0] _T_41; // @[Counter.scala 166:26:@1617.4]
  wire [31:0] _T_42; // @[Counter.scala 166:26:@1618.4]
  assign numPushed = io_input_inc_en_0 ? $signed(6'sh1) : $signed(6'sh0); // @[Counter.scala 164:47:@1611.4]
  assign numPopped = io_input_dinc_en_0 ? $signed(6'sh1) : $signed(6'sh0); // @[Counter.scala 165:48:@1612.4]
  assign _GEN_0 = {{26{numPushed[5]}},numPushed}; // @[Counter.scala 166:14:@1613.4]
  assign _T_37 = $signed(cnt) + $signed(_GEN_0); // @[Counter.scala 166:14:@1613.4]
  assign _T_38 = $signed(cnt) + $signed(_GEN_0); // @[Counter.scala 166:14:@1614.4]
  assign _T_39 = $signed(_T_38); // @[Counter.scala 166:14:@1615.4]
  assign _GEN_1 = {{26{numPopped[5]}},numPopped}; // @[Counter.scala 166:26:@1616.4]
  assign _T_40 = $signed(_T_39) - $signed(_GEN_1); // @[Counter.scala 166:26:@1616.4]
  assign _T_41 = $signed(_T_39) - $signed(_GEN_1); // @[Counter.scala 166:26:@1617.4]
  assign _T_42 = $signed(_T_41); // @[Counter.scala 166:26:@1618.4]
  assign io_output_empty = $signed(cnt) == $signed(32'sh0); // @[Counter.scala 170:19:@1625.4]
  assign io_output_full = $signed(cnt) > $signed(32'sh7); // @[Counter.scala 172:18:@1632.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      cnt <= 32'sh0;
    end else begin
      cnt <= _T_42;
    end
  end
endmodule
module Mem1D( // @[:@1640.2]
  input         clock, // @[:@1641.4]
  input  [3:0]  io_r_ofs_0, // @[:@1643.4]
  input  [3:0]  io_w_ofs_0, // @[:@1643.4]
  input  [31:0] io_w_data_0, // @[:@1643.4]
  input         io_w_en_0, // @[:@1643.4]
  output [31:0] io_output // @[:@1643.4]
);
  reg [31:0] _T_127 [0:7]; // @[MemPrimitives.scala 585:18:@1647.4]
  reg [31:0] _RAND_0;
  wire [31:0] _T_127__T_132_data; // @[MemPrimitives.scala 585:18:@1647.4]
  wire [2:0] _T_127__T_132_addr; // @[MemPrimitives.scala 585:18:@1647.4]
  wire [31:0] _T_127__T_130_data; // @[MemPrimitives.scala 585:18:@1647.4]
  wire [2:0] _T_127__T_130_addr; // @[MemPrimitives.scala 585:18:@1647.4]
  wire  _T_127__T_130_mask; // @[MemPrimitives.scala 585:18:@1647.4]
  wire  _T_127__T_130_en; // @[MemPrimitives.scala 585:18:@1647.4]
  wire  wInBound; // @[MemPrimitives.scala 554:32:@1645.4]
  assign _T_127__T_132_addr = io_r_ofs_0[2:0];
  assign _T_127__T_132_data = _T_127[_T_127__T_132_addr]; // @[MemPrimitives.scala 585:18:@1647.4]
  assign _T_127__T_130_data = io_w_data_0;
  assign _T_127__T_130_addr = io_w_ofs_0[2:0];
  assign _T_127__T_130_mask = 1'h1;
  assign _T_127__T_130_en = io_w_en_0 & wInBound;
  assign wInBound = io_w_ofs_0 <= 4'h8; // @[MemPrimitives.scala 554:32:@1645.4]
  assign io_output = _T_127__T_132_data; // @[MemPrimitives.scala 587:17:@1656.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    _T_127[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(_T_127__T_130_en & _T_127__T_130_mask) begin
      _T_127[_T_127__T_130_addr] <= _T_127__T_130_data; // @[MemPrimitives.scala 585:18:@1647.4]
    end
  end
endmodule
module Compactor( // @[:@1658.2]
  input  [31:0] io_in_0_data, // @[:@1661.4]
  output [31:0] io_out_0_data // @[:@1661.4]
);
  assign io_out_0_data = io_in_0_data; // @[MemPrimitives.scala 616:22:@1665.4]
endmodule
module CompactingEnqNetwork( // @[:@1669.2]
  input  [5:0]  io_headCnt, // @[:@1672.4]
  input  [31:0] io_in_0_data, // @[:@1672.4]
  input         io_in_0_en, // @[:@1672.4]
  output [31:0] io_out_0_data, // @[:@1672.4]
  output        io_out_0_en // @[:@1672.4]
);
  wire [31:0] compactor_io_in_0_data; // @[MemPrimitives.scala 638:25:@1675.4]
  wire [31:0] compactor_io_out_0_data; // @[MemPrimitives.scala 638:25:@1675.4]
  wire [5:0] numEnabled; // @[MemPrimitives.scala 634:38:@1674.4]
  wire [5:0] _GEN_0; // @[Math.scala 53:59:@1681.4]
  wire [5:0] current_base_bank; // @[Math.scala 53:59:@1681.4]
  wire [5:0] _T_22; // @[MemPrimitives.scala 644:46:@1682.4]
  wire [6:0] _T_23; // @[MemPrimitives.scala 644:33:@1683.4]
  wire [5:0] _T_24; // @[MemPrimitives.scala 644:33:@1684.4]
  wire [5:0] _T_25; // @[MemPrimitives.scala 644:33:@1685.4]
  wire [6:0] _T_27; // @[MemPrimitives.scala 644:53:@1686.4]
  wire [5:0] _T_28; // @[MemPrimitives.scala 644:53:@1687.4]
  wire [5:0] upper; // @[MemPrimitives.scala 644:53:@1688.4]
  wire  _T_30; // @[MemPrimitives.scala 645:34:@1689.4]
  wire [5:0] num_straddling; // @[MemPrimitives.scala 645:27:@1690.4]
  wire [6:0] _T_33; // @[MemPrimitives.scala 646:42:@1692.4]
  wire [5:0] _T_34; // @[MemPrimitives.scala 646:42:@1693.4]
  wire [5:0] num_straight; // @[MemPrimitives.scala 646:42:@1694.4]
  wire  _T_36; // @[MemPrimitives.scala 648:40:@1695.4]
  wire  _T_38; // @[MemPrimitives.scala 648:73:@1696.4]
  wire  _T_44; // @[MemPrimitives.scala 648:109:@1701.4]
  wire  _T_45; // @[MemPrimitives.scala 648:94:@1702.4]
  wire [6:0] _T_53; // @[MemPrimitives.scala 649:72:@1706.4]
  wire [5:0] _T_54; // @[MemPrimitives.scala 649:72:@1707.4]
  wire [5:0] _T_55; // @[MemPrimitives.scala 649:72:@1708.4]
  wire [6:0] _T_57; // @[MemPrimitives.scala 649:101:@1709.4]
  wire [5:0] _T_58; // @[MemPrimitives.scala 649:101:@1710.4]
  wire [5:0] _T_59; // @[MemPrimitives.scala 649:101:@1711.4]
  wire [5:0] _T_60; // @[MemPrimitives.scala 649:27:@1712.4]
  wire [5:0] _T_62; // @[MemPrimitives.scala 653:57:@1713.4]
  wire  _T_64; // @[Mux.scala 46:19:@1714.4]
  Compactor compactor ( // @[MemPrimitives.scala 638:25:@1675.4]
    .io_in_0_data(compactor_io_in_0_data),
    .io_out_0_data(compactor_io_out_0_data)
  );
  assign numEnabled = io_in_0_en ? 6'h1 : 6'h0; // @[MemPrimitives.scala 634:38:@1674.4]
  assign _GEN_0 = $signed(io_headCnt) % $signed(6'sh1); // @[Math.scala 53:59:@1681.4]
  assign current_base_bank = _GEN_0[5:0]; // @[Math.scala 53:59:@1681.4]
  assign _T_22 = $signed(numEnabled); // @[MemPrimitives.scala 644:46:@1682.4]
  assign _T_23 = $signed(current_base_bank) + $signed(_T_22); // @[MemPrimitives.scala 644:33:@1683.4]
  assign _T_24 = $signed(current_base_bank) + $signed(_T_22); // @[MemPrimitives.scala 644:33:@1684.4]
  assign _T_25 = $signed(_T_24); // @[MemPrimitives.scala 644:33:@1685.4]
  assign _T_27 = $signed(_T_25) - $signed(6'sh1); // @[MemPrimitives.scala 644:53:@1686.4]
  assign _T_28 = $signed(_T_25) - $signed(6'sh1); // @[MemPrimitives.scala 644:53:@1687.4]
  assign upper = $signed(_T_28); // @[MemPrimitives.scala 644:53:@1688.4]
  assign _T_30 = $signed(upper) < $signed(6'sh0); // @[MemPrimitives.scala 645:34:@1689.4]
  assign num_straddling = _T_30 ? $signed(6'sh0) : $signed(upper); // @[MemPrimitives.scala 645:27:@1690.4]
  assign _T_33 = $signed(_T_22) - $signed(num_straddling); // @[MemPrimitives.scala 646:42:@1692.4]
  assign _T_34 = $signed(_T_22) - $signed(num_straddling); // @[MemPrimitives.scala 646:42:@1693.4]
  assign num_straight = $signed(_T_34); // @[MemPrimitives.scala 646:42:@1694.4]
  assign _T_36 = $signed(6'sh0) < $signed(num_straddling); // @[MemPrimitives.scala 648:40:@1695.4]
  assign _T_38 = $signed(6'sh0) >= $signed(current_base_bank); // @[MemPrimitives.scala 648:73:@1696.4]
  assign _T_44 = $signed(6'sh0) < $signed(_T_25); // @[MemPrimitives.scala 648:109:@1701.4]
  assign _T_45 = _T_38 & _T_44; // @[MemPrimitives.scala 648:94:@1702.4]
  assign _T_53 = {{1{num_straight[5]}},num_straight}; // @[MemPrimitives.scala 649:72:@1706.4]
  assign _T_54 = _T_53[5:0]; // @[MemPrimitives.scala 649:72:@1707.4]
  assign _T_55 = $signed(_T_54); // @[MemPrimitives.scala 649:72:@1708.4]
  assign _T_57 = $signed(6'sh0) - $signed(current_base_bank); // @[MemPrimitives.scala 649:101:@1709.4]
  assign _T_58 = $signed(6'sh0) - $signed(current_base_bank); // @[MemPrimitives.scala 649:101:@1710.4]
  assign _T_59 = $signed(_T_58); // @[MemPrimitives.scala 649:101:@1711.4]
  assign _T_60 = _T_36 ? $signed(_T_55) : $signed(_T_59); // @[MemPrimitives.scala 649:27:@1712.4]
  assign _T_62 = $unsigned(_T_60); // @[MemPrimitives.scala 653:57:@1713.4]
  assign _T_64 = 6'h0 == _T_62; // @[Mux.scala 46:19:@1714.4]
  assign io_out_0_data = _T_64 ? compactor_io_out_0_data : 32'h0; // @[MemPrimitives.scala 658:63:@1716.4]
  assign io_out_0_en = _T_36 | _T_45; // @[MemPrimitives.scala 659:63:@1717.4]
  assign compactor_io_in_0_data = io_in_0_data; // @[MemPrimitives.scala 639:19:@1679.4]
endmodule
module CompactingDeqNetwork( // @[:@1719.2]
  input  [5:0]  io_tailCnt, // @[:@1722.4]
  input  [31:0] io_input_data_0, // @[:@1722.4]
  output [31:0] io_output_0 // @[:@1722.4]
);
  wire [5:0] _GEN_0; // @[Math.scala 53:59:@1726.4]
  wire [5:0] current_base_bank; // @[Math.scala 53:59:@1726.4]
  wire [5:0] _T_55; // @[MemPrimitives.scala 685:65:@1749.4]
  wire [6:0] _T_56; // @[MemPrimitives.scala 685:72:@1750.4]
  wire [5:0] _T_57; // @[MemPrimitives.scala 685:72:@1751.4]
  wire [5:0] _GEN_1; // @[Math.scala 55:59:@1752.4]
  wire [5:0] _T_59; // @[Math.scala 55:59:@1752.4]
  wire  _T_62; // @[Mux.scala 46:19:@1753.4]
  assign _GEN_0 = $signed(io_tailCnt) % $signed(6'sh1); // @[Math.scala 53:59:@1726.4]
  assign current_base_bank = _GEN_0[5:0]; // @[Math.scala 53:59:@1726.4]
  assign _T_55 = $unsigned(current_base_bank); // @[MemPrimitives.scala 685:65:@1749.4]
  assign _T_56 = {{1'd0}, _T_55}; // @[MemPrimitives.scala 685:72:@1750.4]
  assign _T_57 = _T_56[5:0]; // @[MemPrimitives.scala 685:72:@1751.4]
  assign _GEN_1 = _T_57 % 6'h1; // @[Math.scala 55:59:@1752.4]
  assign _T_59 = _GEN_1[5:0]; // @[Math.scala 55:59:@1752.4]
  assign _T_62 = 6'h0 == _T_59; // @[Mux.scala 46:19:@1753.4]
  assign io_output_0 = _T_62 ? io_input_data_0 : 32'h0; // @[MemPrimitives.scala 689:18:@1755.4]
endmodule
module x97_a_0( // @[:@1757.2]
  input         clock, // @[:@1758.4]
  input         reset, // @[:@1759.4]
  input         io_rPort_0_en_0, // @[:@1760.4]
  output [31:0] io_rPort_0_output_0, // @[:@1760.4]
  input  [31:0] io_wPort_0_data_0, // @[:@1760.4]
  input         io_wPort_0_en_0, // @[:@1760.4]
  output        io_full, // @[:@1760.4]
  output        io_empty, // @[:@1760.4]
  output        io_accessActivesOut_0, // @[:@1760.4]
  output        io_accessActivesOut_1, // @[:@1760.4]
  input         io_accessActivesIn_0, // @[:@1760.4]
  input         io_accessActivesIn_1 // @[:@1760.4]
);
  wire  headCtr_clock; // @[MemPrimitives.scala 233:23:@1784.4]
  wire  headCtr_reset; // @[MemPrimitives.scala 233:23:@1784.4]
  wire  headCtr_io_input_dir; // @[MemPrimitives.scala 233:23:@1784.4]
  wire  headCtr_io_input_reset; // @[MemPrimitives.scala 233:23:@1784.4]
  wire  headCtr_io_input_enables_0; // @[MemPrimitives.scala 233:23:@1784.4]
  wire [5:0] headCtr_io_output_count; // @[MemPrimitives.scala 233:23:@1784.4]
  wire  tailCtr_clock; // @[MemPrimitives.scala 234:23:@1792.4]
  wire  tailCtr_reset; // @[MemPrimitives.scala 234:23:@1792.4]
  wire  tailCtr_io_input_dir; // @[MemPrimitives.scala 234:23:@1792.4]
  wire  tailCtr_io_input_reset; // @[MemPrimitives.scala 234:23:@1792.4]
  wire  tailCtr_io_input_enables_0; // @[MemPrimitives.scala 234:23:@1792.4]
  wire [5:0] tailCtr_io_output_count; // @[MemPrimitives.scala 234:23:@1792.4]
  wire  elements_clock; // @[MemPrimitives.scala 244:24:@1806.4]
  wire  elements_reset; // @[MemPrimitives.scala 244:24:@1806.4]
  wire  elements_io_input_inc_en_0; // @[MemPrimitives.scala 244:24:@1806.4]
  wire  elements_io_input_dinc_en_0; // @[MemPrimitives.scala 244:24:@1806.4]
  wire  elements_io_output_empty; // @[MemPrimitives.scala 244:24:@1806.4]
  wire  elements_io_output_full; // @[MemPrimitives.scala 244:24:@1806.4]
  wire  m_0_clock; // @[MemPrimitives.scala 250:56:@1820.4]
  wire [3:0] m_0_io_r_ofs_0; // @[MemPrimitives.scala 250:56:@1820.4]
  wire [3:0] m_0_io_w_ofs_0; // @[MemPrimitives.scala 250:56:@1820.4]
  wire [31:0] m_0_io_w_data_0; // @[MemPrimitives.scala 250:56:@1820.4]
  wire  m_0_io_w_en_0; // @[MemPrimitives.scala 250:56:@1820.4]
  wire [31:0] m_0_io_output; // @[MemPrimitives.scala 250:56:@1820.4]
  wire [5:0] enqCompactor_io_headCnt; // @[MemPrimitives.scala 254:28:@1836.4]
  wire [31:0] enqCompactor_io_in_0_data; // @[MemPrimitives.scala 254:28:@1836.4]
  wire  enqCompactor_io_in_0_en; // @[MemPrimitives.scala 254:28:@1836.4]
  wire [31:0] enqCompactor_io_out_0_data; // @[MemPrimitives.scala 254:28:@1836.4]
  wire  enqCompactor_io_out_0_en; // @[MemPrimitives.scala 254:28:@1836.4]
  wire [5:0] deqCompactor_io_tailCnt; // @[MemPrimitives.scala 273:28:@1858.4]
  wire [31:0] deqCompactor_io_input_data_0; // @[MemPrimitives.scala 273:28:@1858.4]
  wire [31:0] deqCompactor_io_output_0; // @[MemPrimitives.scala 273:28:@1858.4]
  wire [5:0] _GEN_0; // @[Math.scala 53:59:@1847.4]
  wire [5:0] active_w_bank; // @[Math.scala 53:59:@1847.4]
  wire [6:0] active_w_addr; // @[Math.scala 52:59:@1848.4]
  wire  _T_94; // @[MemPrimitives.scala 266:38:@1849.4]
  wire [7:0] _T_96; // @[MemPrimitives.scala 266:69:@1850.4]
  wire [6:0] _T_97; // @[MemPrimitives.scala 266:69:@1851.4]
  wire [6:0] _T_98; // @[MemPrimitives.scala 266:69:@1852.4]
  wire [6:0] _T_99; // @[MemPrimitives.scala 266:19:@1853.4]
  wire [6:0] _T_100; // @[MemPrimitives.scala 267:32:@1854.4]
  wire [5:0] _GEN_1; // @[Math.scala 53:59:@1866.4]
  wire [5:0] active_r_bank; // @[Math.scala 53:59:@1866.4]
  wire [6:0] active_r_addr; // @[Math.scala 52:59:@1867.4]
  wire  _T_104; // @[MemPrimitives.scala 279:38:@1868.4]
  wire [7:0] _T_106; // @[MemPrimitives.scala 279:69:@1869.4]
  wire [6:0] _T_107; // @[MemPrimitives.scala 279:69:@1870.4]
  wire [6:0] _T_108; // @[MemPrimitives.scala 279:69:@1871.4]
  wire [6:0] _T_109; // @[MemPrimitives.scala 279:19:@1872.4]
  wire [6:0] _T_110; // @[MemPrimitives.scala 280:32:@1873.4]
  CompactingCounter headCtr ( // @[MemPrimitives.scala 233:23:@1784.4]
    .clock(headCtr_clock),
    .reset(headCtr_reset),
    .io_input_dir(headCtr_io_input_dir),
    .io_input_reset(headCtr_io_input_reset),
    .io_input_enables_0(headCtr_io_input_enables_0),
    .io_output_count(headCtr_io_output_count)
  );
  CompactingCounter tailCtr ( // @[MemPrimitives.scala 234:23:@1792.4]
    .clock(tailCtr_clock),
    .reset(tailCtr_reset),
    .io_input_dir(tailCtr_io_input_dir),
    .io_input_reset(tailCtr_io_input_reset),
    .io_input_enables_0(tailCtr_io_input_enables_0),
    .io_output_count(tailCtr_io_output_count)
  );
  CompactingIncDincCtr elements ( // @[MemPrimitives.scala 244:24:@1806.4]
    .clock(elements_clock),
    .reset(elements_reset),
    .io_input_inc_en_0(elements_io_input_inc_en_0),
    .io_input_dinc_en_0(elements_io_input_dinc_en_0),
    .io_output_empty(elements_io_output_empty),
    .io_output_full(elements_io_output_full)
  );
  Mem1D m_0 ( // @[MemPrimitives.scala 250:56:@1820.4]
    .clock(m_0_clock),
    .io_r_ofs_0(m_0_io_r_ofs_0),
    .io_w_ofs_0(m_0_io_w_ofs_0),
    .io_w_data_0(m_0_io_w_data_0),
    .io_w_en_0(m_0_io_w_en_0),
    .io_output(m_0_io_output)
  );
  CompactingEnqNetwork enqCompactor ( // @[MemPrimitives.scala 254:28:@1836.4]
    .io_headCnt(enqCompactor_io_headCnt),
    .io_in_0_data(enqCompactor_io_in_0_data),
    .io_in_0_en(enqCompactor_io_in_0_en),
    .io_out_0_data(enqCompactor_io_out_0_data),
    .io_out_0_en(enqCompactor_io_out_0_en)
  );
  CompactingDeqNetwork deqCompactor ( // @[MemPrimitives.scala 273:28:@1858.4]
    .io_tailCnt(deqCompactor_io_tailCnt),
    .io_input_data_0(deqCompactor_io_input_data_0),
    .io_output_0(deqCompactor_io_output_0)
  );
  assign _GEN_0 = $signed(headCtr_io_output_count) % $signed(6'sh1); // @[Math.scala 53:59:@1847.4]
  assign active_w_bank = _GEN_0[5:0]; // @[Math.scala 53:59:@1847.4]
  assign active_w_addr = $signed(headCtr_io_output_count) / $signed(6'sh1); // @[Math.scala 52:59:@1848.4]
  assign _T_94 = $signed(6'sh0) < $signed(active_w_bank); // @[MemPrimitives.scala 266:38:@1849.4]
  assign _T_96 = $signed(active_w_addr) + $signed(7'sh1); // @[MemPrimitives.scala 266:69:@1850.4]
  assign _T_97 = $signed(active_w_addr) + $signed(7'sh1); // @[MemPrimitives.scala 266:69:@1851.4]
  assign _T_98 = $signed(_T_97); // @[MemPrimitives.scala 266:69:@1852.4]
  assign _T_99 = _T_94 ? $signed(_T_98) : $signed(active_w_addr); // @[MemPrimitives.scala 266:19:@1853.4]
  assign _T_100 = $unsigned(_T_99); // @[MemPrimitives.scala 267:32:@1854.4]
  assign _GEN_1 = $signed(tailCtr_io_output_count) % $signed(6'sh1); // @[Math.scala 53:59:@1866.4]
  assign active_r_bank = _GEN_1[5:0]; // @[Math.scala 53:59:@1866.4]
  assign active_r_addr = $signed(tailCtr_io_output_count) / $signed(6'sh1); // @[Math.scala 52:59:@1867.4]
  assign _T_104 = $signed(6'sh0) < $signed(active_r_bank); // @[MemPrimitives.scala 279:38:@1868.4]
  assign _T_106 = $signed(active_r_addr) + $signed(7'sh1); // @[MemPrimitives.scala 279:69:@1869.4]
  assign _T_107 = $signed(active_r_addr) + $signed(7'sh1); // @[MemPrimitives.scala 279:69:@1870.4]
  assign _T_108 = $signed(_T_107); // @[MemPrimitives.scala 279:69:@1871.4]
  assign _T_109 = _T_104 ? $signed(_T_108) : $signed(active_r_addr); // @[MemPrimitives.scala 279:19:@1872.4]
  assign _T_110 = $unsigned(_T_109); // @[MemPrimitives.scala 280:32:@1873.4]
  assign io_rPort_0_output_0 = deqCompactor_io_output_0; // @[MemPrimitives.scala 284:82:@1877.4]
  assign io_full = elements_io_output_full; // @[MemPrimitives.scala 291:39:@1881.4]
  assign io_empty = elements_io_output_empty; // @[MemPrimitives.scala 290:40:@1880.4]
  assign io_accessActivesOut_0 = io_accessActivesIn_0; // @[MemPrimitives.scala 289:127:@1878.4]
  assign io_accessActivesOut_1 = io_accessActivesIn_1; // @[MemPrimitives.scala 289:127:@1879.4]
  assign headCtr_clock = clock; // @[:@1785.4]
  assign headCtr_reset = reset; // @[:@1786.4]
  assign headCtr_io_input_dir = 1'h1; // @[MemPrimitives.scala 239:24:@1804.4]
  assign headCtr_io_input_reset = reset; // @[MemPrimitives.scala 237:26:@1802.4]
  assign headCtr_io_input_enables_0 = io_wPort_0_en_0; // @[MemPrimitives.scala 235:129:@1800.4]
  assign tailCtr_clock = clock; // @[:@1793.4]
  assign tailCtr_reset = reset; // @[:@1794.4]
  assign tailCtr_io_input_dir = 1'h1; // @[MemPrimitives.scala 240:24:@1805.4]
  assign tailCtr_io_input_reset = reset; // @[MemPrimitives.scala 238:26:@1803.4]
  assign tailCtr_io_input_enables_0 = io_rPort_0_en_0; // @[MemPrimitives.scala 236:129:@1801.4]
  assign elements_clock = clock; // @[:@1807.4]
  assign elements_reset = reset; // @[:@1808.4]
  assign elements_io_input_inc_en_0 = io_wPort_0_en_0; // @[MemPrimitives.scala 246:79:@1818.4]
  assign elements_io_input_dinc_en_0 = io_rPort_0_en_0; // @[MemPrimitives.scala 247:80:@1819.4]
  assign m_0_clock = clock; // @[:@1821.4]
  assign m_0_io_r_ofs_0 = _T_110[3:0]; // @[MemPrimitives.scala 280:24:@1874.4]
  assign m_0_io_w_ofs_0 = _T_100[3:0]; // @[MemPrimitives.scala 267:24:@1855.4]
  assign m_0_io_w_data_0 = enqCompactor_io_out_0_data; // @[MemPrimitives.scala 268:25:@1856.4]
  assign m_0_io_w_en_0 = enqCompactor_io_out_0_en; // @[MemPrimitives.scala 269:25:@1857.4]
  assign enqCompactor_io_headCnt = headCtr_io_output_count; // @[MemPrimitives.scala 256:27:@1844.4]
  assign enqCompactor_io_in_0_data = io_wPort_0_data_0; // @[MemPrimitives.scala 258:90:@1845.4]
  assign enqCompactor_io_in_0_en = io_wPort_0_en_0; // @[MemPrimitives.scala 259:85:@1846.4]
  assign deqCompactor_io_tailCnt = tailCtr_io_output_count; // @[MemPrimitives.scala 275:27:@1865.4]
  assign deqCompactor_io_input_data_0 = m_0_io_output; // @[MemPrimitives.scala 281:35:@1875.4]
endmodule
module x106_outr_UnitPipe_sm( // @[:@2086.2]
  input   clock, // @[:@2087.4]
  input   reset, // @[:@2088.4]
  input   io_enable, // @[:@2089.4]
  output  io_done, // @[:@2089.4]
  input   io_parentAck, // @[:@2089.4]
  input   io_doneIn_0, // @[:@2089.4]
  output  io_enableOut_0, // @[:@2089.4]
  output  io_childAck_0, // @[:@2089.4]
  input   io_ctrCopyDone_0 // @[:@2089.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@2092.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@2092.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@2092.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@2092.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@2092.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@2092.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@2095.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@2095.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@2095.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@2095.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@2095.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@2095.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@2112.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@2112.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@2112.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@2112.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@2112.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@2112.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@2143.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@2143.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@2143.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@2143.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@2143.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@2157.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@2157.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@2157.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@2157.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@2157.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@2175.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@2175.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@2175.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@2175.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@2175.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@2212.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@2212.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@2212.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@2212.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@2212.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@2229.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@2229.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@2229.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@2229.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@2229.4]
  wire  _T_105; // @[Controllers.scala 165:35:@2127.4]
  wire  _T_107; // @[Controllers.scala 165:60:@2128.4]
  wire  _T_108; // @[Controllers.scala 165:58:@2129.4]
  wire  _T_110; // @[Controllers.scala 165:76:@2130.4]
  wire  _T_111; // @[Controllers.scala 165:74:@2131.4]
  wire  _T_115; // @[Controllers.scala 165:109:@2134.4]
  wire  _T_118; // @[Controllers.scala 165:141:@2136.4]
  wire  _T_126; // @[package.scala 96:25:@2148.4 package.scala 96:25:@2149.4]
  wire  _T_130; // @[Controllers.scala 167:54:@2151.4]
  wire  _T_131; // @[Controllers.scala 167:52:@2152.4]
  wire  _T_138; // @[package.scala 96:25:@2162.4 package.scala 96:25:@2163.4]
  wire  _T_156; // @[package.scala 96:25:@2180.4 package.scala 96:25:@2181.4]
  wire  _T_160; // @[Controllers.scala 169:67:@2183.4]
  wire  _T_161; // @[Controllers.scala 169:86:@2184.4]
  wire  _T_174; // @[Controllers.scala 213:68:@2198.4]
  wire  _T_176; // @[Controllers.scala 213:90:@2200.4]
  wire  _T_178; // @[Controllers.scala 213:132:@2202.4]
  reg  _T_186; // @[package.scala 48:56:@2208.4]
  reg [31:0] _RAND_0;
  wire  _T_187; // @[package.scala 100:41:@2210.4]
  reg  _T_200; // @[package.scala 48:56:@2226.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@2092.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@2095.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@2112.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@2143.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@2157.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@2175.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@2212.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@2229.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_105 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@2127.4]
  assign _T_107 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@2128.4]
  assign _T_108 = _T_105 & _T_107; // @[Controllers.scala 165:58:@2129.4]
  assign _T_110 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@2130.4]
  assign _T_111 = _T_108 & _T_110; // @[Controllers.scala 165:74:@2131.4]
  assign _T_115 = _T_111 & io_enable; // @[Controllers.scala 165:109:@2134.4]
  assign _T_118 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@2136.4]
  assign _T_126 = RetimeWrapper_io_out; // @[package.scala 96:25:@2148.4 package.scala 96:25:@2149.4]
  assign _T_130 = _T_126 == 1'h0; // @[Controllers.scala 167:54:@2151.4]
  assign _T_131 = io_doneIn_0 | _T_130; // @[Controllers.scala 167:52:@2152.4]
  assign _T_138 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@2162.4 package.scala 96:25:@2163.4]
  assign _T_156 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@2180.4 package.scala 96:25:@2181.4]
  assign _T_160 = _T_156 == 1'h0; // @[Controllers.scala 169:67:@2183.4]
  assign _T_161 = _T_160 & io_enable; // @[Controllers.scala 169:86:@2184.4]
  assign _T_174 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@2198.4]
  assign _T_176 = _T_174 & _T_105; // @[Controllers.scala 213:90:@2200.4]
  assign _T_178 = ~ done_0_io_output; // @[Controllers.scala 213:132:@2202.4]
  assign _T_187 = done_0_io_output & _T_186; // @[package.scala 100:41:@2210.4]
  assign io_done = RetimeWrapper_4_io_out; // @[Controllers.scala 245:13:@2236.4]
  assign io_enableOut_0 = _T_176 & _T_178; // @[Controllers.scala 213:55:@2206.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@2197.4]
  assign active_0_clock = clock; // @[:@2093.4]
  assign active_0_reset = reset; // @[:@2094.4]
  assign active_0_io_input_set = _T_115 & _T_118; // @[Controllers.scala 165:32:@2138.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@2142.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@2100.4]
  assign done_0_clock = clock; // @[:@2096.4]
  assign done_0_reset = reset; // @[:@2097.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_161; // @[Controllers.scala 169:30:@2188.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@2110.4 Controllers.scala 170:32:@2195.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@2101.4]
  assign iterDone_0_clock = clock; // @[:@2113.4]
  assign iterDone_0_reset = reset; // @[:@2114.4]
  assign iterDone_0_io_input_set = _T_131 & io_enable; // @[Controllers.scala 167:34:@2156.4]
  assign iterDone_0_io_input_reset = _T_138 | io_parentAck; // @[Controllers.scala 92:37:@2124.4 Controllers.scala 168:36:@2172.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@2115.4]
  assign RetimeWrapper_clock = clock; // @[:@2144.4]
  assign RetimeWrapper_reset = reset; // @[:@2145.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@2147.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@2146.4]
  assign RetimeWrapper_1_clock = clock; // @[:@2158.4]
  assign RetimeWrapper_1_reset = reset; // @[:@2159.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@2161.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@2160.4]
  assign RetimeWrapper_2_clock = clock; // @[:@2176.4]
  assign RetimeWrapper_2_reset = reset; // @[:@2177.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@2179.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@2178.4]
  assign RetimeWrapper_3_clock = clock; // @[:@2213.4]
  assign RetimeWrapper_3_reset = reset; // @[:@2214.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@2216.4]
  assign RetimeWrapper_3_io_in = _T_187 | io_parentAck; // @[package.scala 94:16:@2215.4]
  assign RetimeWrapper_4_clock = clock; // @[:@2230.4]
  assign RetimeWrapper_4_reset = reset; // @[:@2231.4]
  assign RetimeWrapper_4_io_flow = io_enable; // @[package.scala 95:18:@2233.4]
  assign RetimeWrapper_4_io_in = done_0_io_output & _T_200; // @[package.scala 94:16:@2232.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_186 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_200 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_186 <= 1'h0;
    end else begin
      _T_186 <= _T_110;
    end
    if (reset) begin
      _T_200 <= 1'h0;
    end else begin
      _T_200 <= _T_110;
    end
  end
endmodule
module SingleCounter_1( // @[:@2380.2]
  input         clock, // @[:@2381.4]
  input         reset, // @[:@2382.4]
  input         io_setup_saturate, // @[:@2383.4]
  input         io_input_reset, // @[:@2383.4]
  input         io_input_enable, // @[:@2383.4]
  output [31:0] io_output_count_0, // @[:@2383.4]
  output        io_output_oobs_0, // @[:@2383.4]
  output        io_output_done // @[:@2383.4]
);
  wire  bases_0_clock; // @[Counter.scala 253:53:@2396.4]
  wire  bases_0_reset; // @[Counter.scala 253:53:@2396.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 253:53:@2396.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 253:53:@2396.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 253:53:@2396.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 253:53:@2396.4]
  wire  SRFF_clock; // @[Counter.scala 255:22:@2412.4]
  wire  SRFF_reset; // @[Counter.scala 255:22:@2412.4]
  wire  SRFF_io_input_set; // @[Counter.scala 255:22:@2412.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 255:22:@2412.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 255:22:@2412.4]
  wire  SRFF_io_output; // @[Counter.scala 255:22:@2412.4]
  wire  _T_36; // @[Counter.scala 256:45:@2415.4]
  wire [31:0] _T_48; // @[Counter.scala 279:52:@2440.4]
  wire [32:0] _T_50; // @[Counter.scala 283:33:@2441.4]
  wire [31:0] _T_51; // @[Counter.scala 283:33:@2442.4]
  wire [31:0] _T_52; // @[Counter.scala 283:33:@2443.4]
  wire  _T_57; // @[Counter.scala 285:18:@2445.4]
  wire [31:0] _T_68; // @[Counter.scala 291:115:@2453.4]
  wire [31:0] _T_70; // @[Counter.scala 291:85:@2455.4]
  wire [31:0] _T_71; // @[Counter.scala 291:152:@2456.4]
  wire [31:0] _T_72; // @[Counter.scala 291:74:@2457.4]
  wire  _T_75; // @[Counter.scala 314:102:@2461.4]
  wire  _T_77; // @[Counter.scala 314:130:@2462.4]
  FF bases_0 ( // @[Counter.scala 253:53:@2396.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 255:22:@2412.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 256:45:@2415.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 279:52:@2440.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@2441.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@2442.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 283:33:@2443.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh40); // @[Counter.scala 285:18:@2445.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 291:115:@2453.4]
  assign _T_70 = io_setup_saturate ? _T_68 : 32'h0; // @[Counter.scala 291:85:@2455.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 291:152:@2456.4]
  assign _T_72 = _T_57 ? _T_70 : _T_71; // @[Counter.scala 291:74:@2457.4]
  assign _T_75 = $signed(_T_48) < $signed(32'sh0); // @[Counter.scala 314:102:@2461.4]
  assign _T_77 = $signed(_T_48) >= $signed(32'sh40); // @[Counter.scala 314:130:@2462.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 296:28:@2460.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 314:60:@2464.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 325:20:@2466.4]
  assign bases_0_clock = clock; // @[:@2397.4]
  assign bases_0_reset = reset; // @[:@2398.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 291:31:@2459.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 273:27:@2438.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 276:29:@2439.4]
  assign SRFF_clock = clock; // @[:@2413.4]
  assign SRFF_reset = reset; // @[:@2414.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 256:23:@2417.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 257:25:@2419.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 258:30:@2420.4]
endmodule
module x99_ctrchain( // @[:@2471.2]
  input         clock, // @[:@2472.4]
  input         reset, // @[:@2473.4]
  input         io_input_reset, // @[:@2474.4]
  input         io_input_enable, // @[:@2474.4]
  output [31:0] io_output_counts_0, // @[:@2474.4]
  output        io_output_oobs_0, // @[:@2474.4]
  output        io_output_done // @[:@2474.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 505:46:@2476.4]
  wire  ctrs_0_reset; // @[Counter.scala 505:46:@2476.4]
  wire  ctrs_0_io_setup_saturate; // @[Counter.scala 505:46:@2476.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 505:46:@2476.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 505:46:@2476.4]
  wire [31:0] ctrs_0_io_output_count_0; // @[Counter.scala 505:46:@2476.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 505:46:@2476.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 505:46:@2476.4]
  reg  wasDone; // @[Counter.scala 534:24:@2485.4]
  reg [31:0] _RAND_0;
  wire  _T_45; // @[Counter.scala 538:69:@2491.4]
  wire  _T_47; // @[Counter.scala 538:80:@2492.4]
  reg  doneLatch; // @[Counter.scala 542:26:@2497.4]
  reg [31:0] _RAND_1;
  wire  _T_54; // @[Counter.scala 543:48:@2498.4]
  wire  _T_55; // @[Counter.scala 543:19:@2499.4]
  SingleCounter_1 ctrs_0 ( // @[Counter.scala 505:46:@2476.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_setup_saturate(ctrs_0_io_setup_saturate),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done)
  );
  assign _T_45 = io_input_enable & ctrs_0_io_output_done; // @[Counter.scala 538:69:@2491.4]
  assign _T_47 = wasDone == 1'h0; // @[Counter.scala 538:80:@2492.4]
  assign _T_54 = ctrs_0_io_output_done ? 1'h1 : doneLatch; // @[Counter.scala 543:48:@2498.4]
  assign _T_55 = io_input_reset ? 1'h0 : _T_54; // @[Counter.scala 543:19:@2499.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 549:32:@2501.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 550:30:@2503.4]
  assign io_output_done = _T_45 & _T_47; // @[Counter.scala 538:18:@2494.4]
  assign ctrs_0_clock = clock; // @[:@2477.4]
  assign ctrs_0_reset = reset; // @[:@2478.4]
  assign ctrs_0_io_setup_saturate = 1'h1; // @[Counter.scala 522:29:@2484.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 512:24:@2482.4]
  assign ctrs_0_io_input_enable = io_input_enable; // @[Counter.scala 516:33:@2483.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= ctrs_0_io_output_done;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (ctrs_0_io_output_done) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module RetimeWrapper_25( // @[:@2543.2]
  input   clock, // @[:@2544.4]
  input   reset, // @[:@2545.4]
  input   io_flow, // @[:@2546.4]
  input   io_in, // @[:@2546.4]
  output  io_out // @[:@2546.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@2548.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@2548.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@2548.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@2548.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@2548.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@2548.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@2548.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@2561.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@2560.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@2559.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@2558.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@2557.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@2555.4]
endmodule
module x105_inr_Foreach_sm( // @[:@2691.2]
  input   clock, // @[:@2692.4]
  input   reset, // @[:@2693.4]
  input   io_enable, // @[:@2694.4]
  output  io_done, // @[:@2694.4]
  output  io_doneLatch, // @[:@2694.4]
  input   io_ctrDone, // @[:@2694.4]
  output  io_datapathEn, // @[:@2694.4]
  output  io_ctrInc, // @[:@2694.4]
  output  io_ctrRst, // @[:@2694.4]
  input   io_parentAck, // @[:@2694.4]
  input   io_backpressure, // @[:@2694.4]
  input   io_break // @[:@2694.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@2696.4]
  wire  active_reset; // @[Controllers.scala 261:22:@2696.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@2696.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@2696.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@2696.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@2696.4]
  wire  done_clock; // @[Controllers.scala 262:20:@2699.4]
  wire  done_reset; // @[Controllers.scala 262:20:@2699.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@2699.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@2699.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@2699.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@2699.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@2733.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@2733.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@2733.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@2733.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@2733.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@2755.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@2755.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@2755.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@2755.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@2755.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@2767.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@2767.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@2767.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@2767.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@2767.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@2775.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@2775.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@2775.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@2775.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@2775.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@2791.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@2791.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@2791.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@2791.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@2791.4]
  wire  _T_80; // @[Controllers.scala 264:48:@2704.4]
  wire  _T_81; // @[Controllers.scala 264:46:@2705.4]
  wire  _T_82; // @[Controllers.scala 264:62:@2706.4]
  wire  _T_83; // @[Controllers.scala 264:60:@2707.4]
  wire  _T_100; // @[package.scala 100:49:@2724.4]
  reg  _T_103; // @[package.scala 48:56:@2725.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@2738.4 package.scala 96:25:@2739.4]
  wire  _T_110; // @[package.scala 100:49:@2740.4]
  reg  _T_113; // @[package.scala 48:56:@2741.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@2743.4]
  wire  _T_118; // @[Controllers.scala 283:41:@2748.4]
  wire  _T_119; // @[Controllers.scala 283:59:@2749.4]
  wire  _T_121; // @[Controllers.scala 284:37:@2752.4]
  wire  _T_124; // @[package.scala 96:25:@2760.4 package.scala 96:25:@2761.4]
  wire  _T_126; // @[package.scala 100:49:@2762.4]
  reg  _T_129; // @[package.scala 48:56:@2763.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@2785.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@2787.4]
  reg  _T_153; // @[package.scala 48:56:@2788.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@2796.4 package.scala 96:25:@2797.4]
  wire  _T_158; // @[Controllers.scala 292:61:@2798.4]
  wire  _T_159; // @[Controllers.scala 292:24:@2799.4]
  SRFF active ( // @[Controllers.scala 261:22:@2696.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@2699.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_25 RetimeWrapper ( // @[package.scala 93:22:@2733.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_1 ( // @[package.scala 93:22:@2755.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@2767.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@2775.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@2791.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@2704.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@2705.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@2706.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@2707.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@2724.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@2738.4 package.scala 96:25:@2739.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@2740.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@2743.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@2748.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@2749.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@2752.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@2760.4 package.scala 96:25:@2761.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@2762.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@2787.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@2796.4 package.scala 96:25:@2797.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@2798.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@2799.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@2766.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@2801.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@2751.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@2754.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@2746.4]
  assign active_clock = clock; // @[:@2697.4]
  assign active_reset = reset; // @[:@2698.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@2709.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@2713.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@2714.4]
  assign done_clock = clock; // @[:@2700.4]
  assign done_reset = reset; // @[:@2701.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@2729.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@2722.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@2723.4]
  assign RetimeWrapper_clock = clock; // @[:@2734.4]
  assign RetimeWrapper_reset = reset; // @[:@2735.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@2737.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@2736.4]
  assign RetimeWrapper_1_clock = clock; // @[:@2756.4]
  assign RetimeWrapper_1_reset = reset; // @[:@2757.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@2759.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@2758.4]
  assign RetimeWrapper_2_clock = clock; // @[:@2768.4]
  assign RetimeWrapper_2_reset = reset; // @[:@2769.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@2771.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@2770.4]
  assign RetimeWrapper_3_clock = clock; // @[:@2776.4]
  assign RetimeWrapper_3_reset = reset; // @[:@2777.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@2779.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@2778.4]
  assign RetimeWrapper_4_clock = clock; // @[:@2792.4]
  assign RetimeWrapper_4_reset = reset; // @[:@2793.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@2795.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@2794.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module fix2fixBox( // @[:@2955.2]
  input  [31:0] io_a, // @[:@2958.4]
  output [31:0] io_b // @[:@2958.4]
);
  assign io_b = io_a; // @[Converter.scala 95:38:@2968.4]
endmodule
module _( // @[:@2970.2]
  input  [31:0] io_b, // @[:@2973.4]
  output [31:0] io_result // @[:@2973.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@2978.4]
  wire [31:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@2978.4]
  fix2fixBox fix2fixBox ( // @[BigIPZynq.scala 219:30:@2978.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 706:17:@2986.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@2981.4]
endmodule
module RetimeWrapper_33( // @[:@3000.2]
  input         clock, // @[:@3001.4]
  input         reset, // @[:@3002.4]
  input         io_flow, // @[:@3003.4]
  input  [31:0] io_in, // @[:@3003.4]
  output [31:0] io_out // @[:@3003.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@3005.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@3005.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@3005.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3005.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3005.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3005.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@3005.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3018.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3017.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@3016.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3015.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3014.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3012.4]
endmodule
module x105_inr_Foreach_kernelx105_inr_Foreach_concrete1( // @[:@3084.2]
  input         clock, // @[:@3085.4]
  input         reset, // @[:@3086.4]
  output [31:0] io_in_x97_a_0_wPort_0_data_0, // @[:@3087.4]
  output        io_in_x97_a_0_wPort_0_en_0, // @[:@3087.4]
  input         io_in_x97_a_0_full, // @[:@3087.4]
  input         io_in_x97_a_0_accessActivesOut_0, // @[:@3087.4]
  output        io_in_x97_a_0_accessActivesIn_0, // @[:@3087.4]
  input         io_in_x90_TVALID, // @[:@3087.4]
  output        io_in_x90_TREADY, // @[:@3087.4]
  input  [63:0] io_in_x90_TDATA, // @[:@3087.4]
  input  [7:0]  io_in_x90_TID, // @[:@3087.4]
  input  [7:0]  io_in_x90_TDEST, // @[:@3087.4]
  output [63:0] io_in_instrctrs_3_cycs, // @[:@3087.4]
  output [63:0] io_in_instrctrs_3_iters, // @[:@3087.4]
  output [63:0] io_in_instrctrs_3_stalls, // @[:@3087.4]
  output [63:0] io_in_instrctrs_3_idles, // @[:@3087.4]
  input         io_sigsIn_done, // @[:@3087.4]
  input         io_sigsIn_backpressure, // @[:@3087.4]
  input         io_sigsIn_datapathEn, // @[:@3087.4]
  input         io_sigsIn_baseEn, // @[:@3087.4]
  input         io_sigsIn_break, // @[:@3087.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@3087.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@3087.4]
  input         io_rr // @[:@3087.4]
);
  wire  cycles_clock; // @[sm_x105_inr_Foreach.scala 63:26:@3147.4]
  wire  cycles_reset; // @[sm_x105_inr_Foreach.scala 63:26:@3147.4]
  wire  cycles_io_enable; // @[sm_x105_inr_Foreach.scala 63:26:@3147.4]
  wire [63:0] cycles_io_count; // @[sm_x105_inr_Foreach.scala 63:26:@3147.4]
  wire  iters_clock; // @[sm_x105_inr_Foreach.scala 64:25:@3150.4]
  wire  iters_reset; // @[sm_x105_inr_Foreach.scala 64:25:@3150.4]
  wire  iters_io_enable; // @[sm_x105_inr_Foreach.scala 64:25:@3150.4]
  wire [63:0] iters_io_count; // @[sm_x105_inr_Foreach.scala 64:25:@3150.4]
  wire  stalls_clock; // @[sm_x105_inr_Foreach.scala 67:26:@3159.4]
  wire  stalls_reset; // @[sm_x105_inr_Foreach.scala 67:26:@3159.4]
  wire  stalls_io_enable; // @[sm_x105_inr_Foreach.scala 67:26:@3159.4]
  wire [63:0] stalls_io_count; // @[sm_x105_inr_Foreach.scala 67:26:@3159.4]
  wire  idles_clock; // @[sm_x105_inr_Foreach.scala 68:25:@3162.4]
  wire  idles_reset; // @[sm_x105_inr_Foreach.scala 68:25:@3162.4]
  wire  idles_io_enable; // @[sm_x105_inr_Foreach.scala 68:25:@3162.4]
  wire [63:0] idles_io_count; // @[sm_x105_inr_Foreach.scala 68:25:@3162.4]
  wire [31:0] __io_b; // @[Math.scala 709:24:@3182.4]
  wire [31:0] __io_result; // @[Math.scala 709:24:@3182.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3202.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3202.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3202.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@3202.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@3202.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@3213.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@3213.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@3213.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@3213.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@3213.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@3224.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@3224.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@3224.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@3224.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@3224.4]
  wire  _T_312; // @[package.scala 100:49:@3154.4]
  reg  _T_315; // @[package.scala 48:56:@3155.4]
  reg [31:0] _RAND_0;
  wire  _T_317; // @[sm_x105_inr_Foreach.scala 69:49:@3165.4]
  wire  _T_318; // @[sm_x105_inr_Foreach.scala 69:65:@3166.4]
  wire  _T_319; // @[sm_x105_inr_Foreach.scala 69:63:@3167.4]
  wire  _T_320; // @[sm_x105_inr_Foreach.scala 69:46:@3168.4]
  wire  _T_322; // @[sm_x105_inr_Foreach.scala 70:45:@3171.4]
  wire  b101; // @[sm_x105_inr_Foreach.scala 73:18:@3190.4]
  wire  _T_337; // @[sm_x105_inr_Foreach.scala 75:25:@3192.4]
  wire  _T_340; // @[sm_x105_inr_Foreach.scala 77:63:@3196.4]
  wire  _T_341; // @[sm_x105_inr_Foreach.scala 77:50:@3197.4]
  wire  _T_343; // @[sm_x105_inr_Foreach.scala 77:87:@3198.4]
  wire  _T_357; // @[sm_x105_inr_Foreach.scala 88:115:@3221.4]
  wire  _T_361; // @[package.scala 96:25:@3229.4 package.scala 96:25:@3230.4]
  wire  _T_363; // @[implicits.scala 55:10:@3231.4]
  wire  _T_364; // @[sm_x105_inr_Foreach.scala 88:132:@3232.4]
  wire  _T_366; // @[sm_x105_inr_Foreach.scala 88:219:@3234.4]
  wire  _T_367; // @[sm_x105_inr_Foreach.scala 88:238:@3235.4]
  wire  x167_b101_D1; // @[package.scala 96:25:@3218.4 package.scala 96:25:@3219.4]
  InstrumentationCounter cycles ( // @[sm_x105_inr_Foreach.scala 63:26:@3147.4]
    .clock(cycles_clock),
    .reset(cycles_reset),
    .io_enable(cycles_io_enable),
    .io_count(cycles_io_count)
  );
  InstrumentationCounter iters ( // @[sm_x105_inr_Foreach.scala 64:25:@3150.4]
    .clock(iters_clock),
    .reset(iters_reset),
    .io_enable(iters_io_enable),
    .io_count(iters_io_count)
  );
  InstrumentationCounter stalls ( // @[sm_x105_inr_Foreach.scala 67:26:@3159.4]
    .clock(stalls_clock),
    .reset(stalls_reset),
    .io_enable(stalls_io_enable),
    .io_count(stalls_io_count)
  );
  InstrumentationCounter idles ( // @[sm_x105_inr_Foreach.scala 68:25:@3162.4]
    .clock(idles_clock),
    .reset(idles_reset),
    .io_enable(idles_io_enable),
    .io_count(idles_io_count)
  );
  _ _ ( // @[Math.scala 709:24:@3182.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  RetimeWrapper_33 RetimeWrapper ( // @[package.scala 93:22:@3202.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@3213.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@3224.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  assign _T_312 = io_sigsIn_done == 1'h0; // @[package.scala 100:49:@3154.4]
  assign _T_317 = ~ io_in_x97_a_0_full; // @[sm_x105_inr_Foreach.scala 69:49:@3165.4]
  assign _T_318 = ~ io_in_x97_a_0_accessActivesOut_0; // @[sm_x105_inr_Foreach.scala 69:65:@3166.4]
  assign _T_319 = _T_317 | _T_318; // @[sm_x105_inr_Foreach.scala 69:63:@3167.4]
  assign _T_320 = ~ _T_319; // @[sm_x105_inr_Foreach.scala 69:46:@3168.4]
  assign _T_322 = ~ io_in_x90_TVALID; // @[sm_x105_inr_Foreach.scala 70:45:@3171.4]
  assign b101 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x105_inr_Foreach.scala 73:18:@3190.4]
  assign _T_337 = b101 & io_sigsIn_datapathEn; // @[sm_x105_inr_Foreach.scala 75:25:@3192.4]
  assign _T_340 = io_in_x90_TID == 8'h0; // @[sm_x105_inr_Foreach.scala 77:63:@3196.4]
  assign _T_341 = _T_337 & _T_340; // @[sm_x105_inr_Foreach.scala 77:50:@3197.4]
  assign _T_343 = io_in_x90_TDEST == 8'h0; // @[sm_x105_inr_Foreach.scala 77:87:@3198.4]
  assign _T_357 = ~ io_sigsIn_break; // @[sm_x105_inr_Foreach.scala 88:115:@3221.4]
  assign _T_361 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@3229.4 package.scala 96:25:@3230.4]
  assign _T_363 = io_rr ? _T_361 : 1'h0; // @[implicits.scala 55:10:@3231.4]
  assign _T_364 = _T_357 & _T_363; // @[sm_x105_inr_Foreach.scala 88:132:@3232.4]
  assign _T_366 = _T_364 & _T_357; // @[sm_x105_inr_Foreach.scala 88:219:@3234.4]
  assign _T_367 = _T_366 & io_sigsIn_backpressure; // @[sm_x105_inr_Foreach.scala 88:238:@3235.4]
  assign x167_b101_D1 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@3218.4 package.scala 96:25:@3219.4]
  assign io_in_x97_a_0_wPort_0_data_0 = RetimeWrapper_io_out; // @[MemInterfaceType.scala 90:56:@3237.4]
  assign io_in_x97_a_0_wPort_0_en_0 = _T_367 & x167_b101_D1; // @[MemInterfaceType.scala 93:57:@3239.4]
  assign io_in_x97_a_0_accessActivesIn_0 = RetimeWrapper_1_io_out; // @[MemInterfaceType.scala 148:24:@3240.4]
  assign io_in_x90_TREADY = _T_341 & _T_343; // @[sm_x105_inr_Foreach.scala 75:17:@3193.4 sm_x105_inr_Foreach.scala 77:17:@3200.4]
  assign io_in_instrctrs_3_cycs = cycles_io_count; // @[Ledger.scala 282:21:@3174.4]
  assign io_in_instrctrs_3_iters = iters_io_count; // @[Ledger.scala 283:22:@3175.4]
  assign io_in_instrctrs_3_stalls = stalls_io_count; // @[Ledger.scala 284:23:@3176.4]
  assign io_in_instrctrs_3_idles = idles_io_count; // @[Ledger.scala 285:22:@3177.4]
  assign cycles_clock = clock; // @[:@3148.4]
  assign cycles_reset = reset; // @[:@3149.4]
  assign cycles_io_enable = io_sigsIn_baseEn; // @[sm_x105_inr_Foreach.scala 65:24:@3153.4]
  assign iters_clock = clock; // @[:@3151.4]
  assign iters_reset = reset; // @[:@3152.4]
  assign iters_io_enable = io_sigsIn_done & _T_315; // @[sm_x105_inr_Foreach.scala 66:23:@3158.4]
  assign stalls_clock = clock; // @[:@3160.4]
  assign stalls_reset = reset; // @[:@3161.4]
  assign stalls_io_enable = io_sigsIn_baseEn & _T_320; // @[sm_x105_inr_Foreach.scala 69:24:@3170.4]
  assign idles_clock = clock; // @[:@3163.4]
  assign idles_reset = reset; // @[:@3164.4]
  assign idles_io_enable = io_sigsIn_baseEn & _T_322; // @[sm_x105_inr_Foreach.scala 70:23:@3173.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 710:17:@3185.4]
  assign RetimeWrapper_clock = clock; // @[:@3203.4]
  assign RetimeWrapper_reset = reset; // @[:@3204.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@3206.4]
  assign RetimeWrapper_io_in = io_in_x90_TDATA[31:0]; // @[package.scala 94:16:@3205.4]
  assign RetimeWrapper_1_clock = clock; // @[:@3214.4]
  assign RetimeWrapper_1_reset = reset; // @[:@3215.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@3217.4]
  assign RetimeWrapper_1_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@3216.4]
  assign RetimeWrapper_2_clock = clock; // @[:@3225.4]
  assign RetimeWrapper_2_reset = reset; // @[:@3226.4]
  assign RetimeWrapper_2_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@3228.4]
  assign RetimeWrapper_2_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@3227.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_315 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_315 <= 1'h0;
    end else begin
      _T_315 <= _T_312;
    end
  end
endmodule
module x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1( // @[:@3242.2]
  input         clock, // @[:@3243.4]
  input         reset, // @[:@3244.4]
  output [31:0] io_in_x97_a_0_wPort_0_data_0, // @[:@3245.4]
  output        io_in_x97_a_0_wPort_0_en_0, // @[:@3245.4]
  input         io_in_x97_a_0_full, // @[:@3245.4]
  input         io_in_x97_a_0_accessActivesOut_0, // @[:@3245.4]
  output        io_in_x97_a_0_accessActivesIn_0, // @[:@3245.4]
  input         io_in_x90_TVALID, // @[:@3245.4]
  output        io_in_x90_TREADY, // @[:@3245.4]
  input  [63:0] io_in_x90_TDATA, // @[:@3245.4]
  input  [7:0]  io_in_x90_TID, // @[:@3245.4]
  input  [7:0]  io_in_x90_TDEST, // @[:@3245.4]
  output [63:0] io_in_instrctrs_2_cycs, // @[:@3245.4]
  output [63:0] io_in_instrctrs_2_iters, // @[:@3245.4]
  output [63:0] io_in_instrctrs_3_cycs, // @[:@3245.4]
  output [63:0] io_in_instrctrs_3_iters, // @[:@3245.4]
  output [63:0] io_in_instrctrs_3_stalls, // @[:@3245.4]
  output [63:0] io_in_instrctrs_3_idles, // @[:@3245.4]
  input         io_sigsIn_done, // @[:@3245.4]
  input         io_sigsIn_baseEn, // @[:@3245.4]
  input         io_sigsIn_smEnableOuts_0, // @[:@3245.4]
  input         io_sigsIn_smChildAcks_0, // @[:@3245.4]
  output        io_sigsOut_smDoneIn_0, // @[:@3245.4]
  output        io_sigsOut_smCtrCopyDone_0, // @[:@3245.4]
  input         io_rr // @[:@3245.4]
);
  wire  cycles_clock; // @[sm_x106_outr_UnitPipe.scala 63:26:@3305.4]
  wire  cycles_reset; // @[sm_x106_outr_UnitPipe.scala 63:26:@3305.4]
  wire  cycles_io_enable; // @[sm_x106_outr_UnitPipe.scala 63:26:@3305.4]
  wire [63:0] cycles_io_count; // @[sm_x106_outr_UnitPipe.scala 63:26:@3305.4]
  wire  iters_clock; // @[sm_x106_outr_UnitPipe.scala 64:25:@3308.4]
  wire  iters_reset; // @[sm_x106_outr_UnitPipe.scala 64:25:@3308.4]
  wire  iters_io_enable; // @[sm_x106_outr_UnitPipe.scala 64:25:@3308.4]
  wire [63:0] iters_io_count; // @[sm_x106_outr_UnitPipe.scala 64:25:@3308.4]
  wire  x99_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@3321.4]
  wire  x99_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@3321.4]
  wire  x99_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@3321.4]
  wire  x99_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@3321.4]
  wire [31:0] x99_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@3321.4]
  wire  x99_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@3321.4]
  wire  x99_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@3321.4]
  wire  x105_inr_Foreach_sm_clock; // @[sm_x105_inr_Foreach.scala 33:18:@3373.4]
  wire  x105_inr_Foreach_sm_reset; // @[sm_x105_inr_Foreach.scala 33:18:@3373.4]
  wire  x105_inr_Foreach_sm_io_enable; // @[sm_x105_inr_Foreach.scala 33:18:@3373.4]
  wire  x105_inr_Foreach_sm_io_done; // @[sm_x105_inr_Foreach.scala 33:18:@3373.4]
  wire  x105_inr_Foreach_sm_io_doneLatch; // @[sm_x105_inr_Foreach.scala 33:18:@3373.4]
  wire  x105_inr_Foreach_sm_io_ctrDone; // @[sm_x105_inr_Foreach.scala 33:18:@3373.4]
  wire  x105_inr_Foreach_sm_io_datapathEn; // @[sm_x105_inr_Foreach.scala 33:18:@3373.4]
  wire  x105_inr_Foreach_sm_io_ctrInc; // @[sm_x105_inr_Foreach.scala 33:18:@3373.4]
  wire  x105_inr_Foreach_sm_io_ctrRst; // @[sm_x105_inr_Foreach.scala 33:18:@3373.4]
  wire  x105_inr_Foreach_sm_io_parentAck; // @[sm_x105_inr_Foreach.scala 33:18:@3373.4]
  wire  x105_inr_Foreach_sm_io_backpressure; // @[sm_x105_inr_Foreach.scala 33:18:@3373.4]
  wire  x105_inr_Foreach_sm_io_break; // @[sm_x105_inr_Foreach.scala 33:18:@3373.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3401.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3401.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3401.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@3401.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@3401.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@3444.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@3444.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@3444.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@3444.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@3444.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@3452.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@3452.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@3452.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@3452.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@3452.4]
  wire  x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_clock; // @[sm_x105_inr_Foreach.scala 91:24:@3484.4]
  wire  x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_reset; // @[sm_x105_inr_Foreach.scala 91:24:@3484.4]
  wire [31:0] x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_in_x97_a_0_wPort_0_data_0; // @[sm_x105_inr_Foreach.scala 91:24:@3484.4]
  wire  x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_in_x97_a_0_wPort_0_en_0; // @[sm_x105_inr_Foreach.scala 91:24:@3484.4]
  wire  x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_in_x97_a_0_full; // @[sm_x105_inr_Foreach.scala 91:24:@3484.4]
  wire  x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_in_x97_a_0_accessActivesOut_0; // @[sm_x105_inr_Foreach.scala 91:24:@3484.4]
  wire  x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_in_x97_a_0_accessActivesIn_0; // @[sm_x105_inr_Foreach.scala 91:24:@3484.4]
  wire  x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_in_x90_TVALID; // @[sm_x105_inr_Foreach.scala 91:24:@3484.4]
  wire  x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_in_x90_TREADY; // @[sm_x105_inr_Foreach.scala 91:24:@3484.4]
  wire [63:0] x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_in_x90_TDATA; // @[sm_x105_inr_Foreach.scala 91:24:@3484.4]
  wire [7:0] x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_in_x90_TID; // @[sm_x105_inr_Foreach.scala 91:24:@3484.4]
  wire [7:0] x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_in_x90_TDEST; // @[sm_x105_inr_Foreach.scala 91:24:@3484.4]
  wire [63:0] x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_in_instrctrs_3_cycs; // @[sm_x105_inr_Foreach.scala 91:24:@3484.4]
  wire [63:0] x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_in_instrctrs_3_iters; // @[sm_x105_inr_Foreach.scala 91:24:@3484.4]
  wire [63:0] x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_in_instrctrs_3_stalls; // @[sm_x105_inr_Foreach.scala 91:24:@3484.4]
  wire [63:0] x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_in_instrctrs_3_idles; // @[sm_x105_inr_Foreach.scala 91:24:@3484.4]
  wire  x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_sigsIn_done; // @[sm_x105_inr_Foreach.scala 91:24:@3484.4]
  wire  x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_sigsIn_backpressure; // @[sm_x105_inr_Foreach.scala 91:24:@3484.4]
  wire  x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x105_inr_Foreach.scala 91:24:@3484.4]
  wire  x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_sigsIn_baseEn; // @[sm_x105_inr_Foreach.scala 91:24:@3484.4]
  wire  x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x105_inr_Foreach.scala 91:24:@3484.4]
  wire [31:0] x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x105_inr_Foreach.scala 91:24:@3484.4]
  wire  x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x105_inr_Foreach.scala 91:24:@3484.4]
  wire  x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_rr; // @[sm_x105_inr_Foreach.scala 91:24:@3484.4]
  wire  _T_312; // @[package.scala 100:49:@3312.4]
  reg  _T_315; // @[package.scala 48:56:@3313.4]
  reg [31:0] _RAND_0;
  wire  _T_379; // @[package.scala 96:25:@3406.4 package.scala 96:25:@3407.4]
  wire  _T_382; // @[sm_x106_outr_UnitPipe.scala 74:41:@3410.4]
  wire  _T_383; // @[sm_x106_outr_UnitPipe.scala 74:57:@3411.4]
  wire  _T_384; // @[sm_x106_outr_UnitPipe.scala 74:55:@3412.4]
  wire  x105_inr_Foreach_sigsIn_forwardpressure; // @[sm_x106_outr_UnitPipe.scala 75:53:@3415.4]
  wire  _T_395; // @[package.scala 96:25:@3449.4 package.scala 96:25:@3450.4]
  wire  _T_401; // @[package.scala 96:25:@3457.4 package.scala 96:25:@3458.4]
  wire  _T_404; // @[SpatialBlocks.scala 110:93:@3460.4]
  wire  x105_inr_Foreach_sigsIn_baseEn; // @[SpatialBlocks.scala 110:90:@3461.4]
  wire  _T_406; // @[SpatialBlocks.scala 128:36:@3469.4]
  wire  _T_407; // @[SpatialBlocks.scala 128:78:@3470.4]
  wire  _T_412; // @[SpatialBlocks.scala 130:61:@3479.4]
  InstrumentationCounter cycles ( // @[sm_x106_outr_UnitPipe.scala 63:26:@3305.4]
    .clock(cycles_clock),
    .reset(cycles_reset),
    .io_enable(cycles_io_enable),
    .io_count(cycles_io_count)
  );
  InstrumentationCounter iters ( // @[sm_x106_outr_UnitPipe.scala 64:25:@3308.4]
    .clock(iters_clock),
    .reset(iters_reset),
    .io_enable(iters_io_enable),
    .io_count(iters_io_count)
  );
  x99_ctrchain x99_ctrchain ( // @[SpatialBlocks.scala 37:22:@3321.4]
    .clock(x99_ctrchain_clock),
    .reset(x99_ctrchain_reset),
    .io_input_reset(x99_ctrchain_io_input_reset),
    .io_input_enable(x99_ctrchain_io_input_enable),
    .io_output_counts_0(x99_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x99_ctrchain_io_output_oobs_0),
    .io_output_done(x99_ctrchain_io_output_done)
  );
  x105_inr_Foreach_sm x105_inr_Foreach_sm ( // @[sm_x105_inr_Foreach.scala 33:18:@3373.4]
    .clock(x105_inr_Foreach_sm_clock),
    .reset(x105_inr_Foreach_sm_reset),
    .io_enable(x105_inr_Foreach_sm_io_enable),
    .io_done(x105_inr_Foreach_sm_io_done),
    .io_doneLatch(x105_inr_Foreach_sm_io_doneLatch),
    .io_ctrDone(x105_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x105_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x105_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x105_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x105_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x105_inr_Foreach_sm_io_backpressure),
    .io_break(x105_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@3401.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@3444.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@3452.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x105_inr_Foreach_kernelx105_inr_Foreach_concrete1 x105_inr_Foreach_kernelx105_inr_Foreach_concrete1 ( // @[sm_x105_inr_Foreach.scala 91:24:@3484.4]
    .clock(x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_clock),
    .reset(x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_reset),
    .io_in_x97_a_0_wPort_0_data_0(x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_in_x97_a_0_wPort_0_data_0),
    .io_in_x97_a_0_wPort_0_en_0(x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_in_x97_a_0_wPort_0_en_0),
    .io_in_x97_a_0_full(x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_in_x97_a_0_full),
    .io_in_x97_a_0_accessActivesOut_0(x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_in_x97_a_0_accessActivesOut_0),
    .io_in_x97_a_0_accessActivesIn_0(x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_in_x97_a_0_accessActivesIn_0),
    .io_in_x90_TVALID(x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_in_x90_TVALID),
    .io_in_x90_TREADY(x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_in_x90_TREADY),
    .io_in_x90_TDATA(x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_in_x90_TDATA),
    .io_in_x90_TID(x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_in_x90_TID),
    .io_in_x90_TDEST(x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_in_x90_TDEST),
    .io_in_instrctrs_3_cycs(x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_in_instrctrs_3_cycs),
    .io_in_instrctrs_3_iters(x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_in_instrctrs_3_iters),
    .io_in_instrctrs_3_stalls(x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_in_instrctrs_3_stalls),
    .io_in_instrctrs_3_idles(x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_in_instrctrs_3_idles),
    .io_sigsIn_done(x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_sigsIn_done),
    .io_sigsIn_backpressure(x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_baseEn(x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_sigsIn_baseEn),
    .io_sigsIn_break(x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_0(x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_rr(x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_rr)
  );
  assign _T_312 = io_sigsIn_done == 1'h0; // @[package.scala 100:49:@3312.4]
  assign _T_379 = RetimeWrapper_io_out; // @[package.scala 96:25:@3406.4 package.scala 96:25:@3407.4]
  assign _T_382 = ~ io_in_x97_a_0_full; // @[sm_x106_outr_UnitPipe.scala 74:41:@3410.4]
  assign _T_383 = ~ io_in_x97_a_0_accessActivesOut_0; // @[sm_x106_outr_UnitPipe.scala 74:57:@3411.4]
  assign _T_384 = _T_382 | _T_383; // @[sm_x106_outr_UnitPipe.scala 74:55:@3412.4]
  assign x105_inr_Foreach_sigsIn_forwardpressure = io_in_x90_TVALID | x105_inr_Foreach_sm_io_doneLatch; // @[sm_x106_outr_UnitPipe.scala 75:53:@3415.4]
  assign _T_395 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@3449.4 package.scala 96:25:@3450.4]
  assign _T_401 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@3457.4 package.scala 96:25:@3458.4]
  assign _T_404 = ~ _T_401; // @[SpatialBlocks.scala 110:93:@3460.4]
  assign x105_inr_Foreach_sigsIn_baseEn = _T_395 & _T_404; // @[SpatialBlocks.scala 110:90:@3461.4]
  assign _T_406 = x105_inr_Foreach_sm_io_datapathEn; // @[SpatialBlocks.scala 128:36:@3469.4]
  assign _T_407 = ~ x105_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 128:78:@3470.4]
  assign _T_412 = x105_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 130:61:@3479.4]
  assign io_in_x97_a_0_wPort_0_data_0 = x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_in_x97_a_0_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@3584.4]
  assign io_in_x97_a_0_wPort_0_en_0 = x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_in_x97_a_0_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@3580.4]
  assign io_in_x97_a_0_accessActivesIn_0 = x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_in_x97_a_0_accessActivesIn_0; // @[MemInterfaceType.scala 69:92:@3587.4]
  assign io_in_x90_TREADY = x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_in_x90_TREADY; // @[sm_x105_inr_Foreach.scala 51:22:@3595.4]
  assign io_in_instrctrs_2_cycs = cycles_io_count; // @[Ledger.scala 282:21:@3317.4]
  assign io_in_instrctrs_2_iters = iters_io_count; // @[Ledger.scala 283:22:@3318.4]
  assign io_in_instrctrs_3_cycs = x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_in_instrctrs_3_cycs; // @[Ledger.scala 291:78:@3600.4]
  assign io_in_instrctrs_3_iters = x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_in_instrctrs_3_iters; // @[Ledger.scala 291:78:@3599.4]
  assign io_in_instrctrs_3_stalls = x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_in_instrctrs_3_stalls; // @[Ledger.scala 291:78:@3598.4]
  assign io_in_instrctrs_3_idles = x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_in_instrctrs_3_idles; // @[Ledger.scala 291:78:@3597.4]
  assign io_sigsOut_smDoneIn_0 = x105_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 127:53:@3467.4]
  assign io_sigsOut_smCtrCopyDone_0 = x105_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 139:125:@3483.4]
  assign cycles_clock = clock; // @[:@3306.4]
  assign cycles_reset = reset; // @[:@3307.4]
  assign cycles_io_enable = io_sigsIn_baseEn; // @[sm_x106_outr_UnitPipe.scala 65:24:@3311.4]
  assign iters_clock = clock; // @[:@3309.4]
  assign iters_reset = reset; // @[:@3310.4]
  assign iters_io_enable = io_sigsIn_done & _T_315; // @[sm_x106_outr_UnitPipe.scala 66:23:@3316.4]
  assign x99_ctrchain_clock = clock; // @[:@3322.4]
  assign x99_ctrchain_reset = reset; // @[:@3323.4]
  assign x99_ctrchain_io_input_reset = x105_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 130:103:@3482.4]
  assign x99_ctrchain_io_input_enable = _T_412 & x105_inr_Foreach_sigsIn_forwardpressure; // @[SpatialBlocks.scala 104:75:@3437.4 SpatialBlocks.scala 130:45:@3481.4]
  assign x105_inr_Foreach_sm_clock = clock; // @[:@3374.4]
  assign x105_inr_Foreach_sm_reset = reset; // @[:@3375.4]
  assign x105_inr_Foreach_sm_io_enable = x105_inr_Foreach_sigsIn_baseEn & x105_inr_Foreach_sigsIn_forwardpressure; // @[SpatialBlocks.scala 112:18:@3464.4]
  assign x105_inr_Foreach_sm_io_ctrDone = io_rr ? _T_379 : 1'h0; // @[sm_x106_outr_UnitPipe.scala 73:38:@3409.4]
  assign x105_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 114:21:@3466.4]
  assign x105_inr_Foreach_sm_io_backpressure = _T_384 | x105_inr_Foreach_sm_io_doneLatch; // @[SpatialBlocks.scala 105:24:@3438.4]
  assign x105_inr_Foreach_sm_io_break = 1'h0; // @[sm_x106_outr_UnitPipe.scala 77:36:@3418.4]
  assign RetimeWrapper_clock = clock; // @[:@3402.4]
  assign RetimeWrapper_reset = reset; // @[:@3403.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@3405.4]
  assign RetimeWrapper_io_in = x99_ctrchain_io_output_done; // @[package.scala 94:16:@3404.4]
  assign RetimeWrapper_1_clock = clock; // @[:@3445.4]
  assign RetimeWrapper_1_reset = reset; // @[:@3446.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@3448.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@3447.4]
  assign RetimeWrapper_2_clock = clock; // @[:@3453.4]
  assign RetimeWrapper_2_reset = reset; // @[:@3454.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@3456.4]
  assign RetimeWrapper_2_io_in = x105_inr_Foreach_sm_io_done; // @[package.scala 94:16:@3455.4]
  assign x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_clock = clock; // @[:@3485.4]
  assign x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_reset = reset; // @[:@3486.4]
  assign x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_in_x97_a_0_full = io_in_x97_a_0_full; // @[MemInterfaceType.scala 151:13:@3573.4]
  assign x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_in_x97_a_0_accessActivesOut_0 = io_in_x97_a_0_accessActivesOut_0; // @[MemInterfaceType.scala 156:25:@3578.4]
  assign x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_in_x90_TVALID = io_in_x90_TVALID; // @[sm_x105_inr_Foreach.scala 51:22:@3596.4]
  assign x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_in_x90_TDATA = io_in_x90_TDATA; // @[sm_x105_inr_Foreach.scala 51:22:@3594.4]
  assign x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_in_x90_TID = io_in_x90_TID; // @[sm_x105_inr_Foreach.scala 51:22:@3590.4]
  assign x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_in_x90_TDEST = io_in_x90_TDEST; // @[sm_x105_inr_Foreach.scala 51:22:@3589.4]
  assign x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_sigsIn_done = x105_inr_Foreach_sm_io_done; // @[sm_x105_inr_Foreach.scala 96:22:@3619.4]
  assign x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_sigsIn_backpressure = _T_384 | x105_inr_Foreach_sm_io_doneLatch; // @[sm_x105_inr_Foreach.scala 96:22:@3615.4]
  assign x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_406 & _T_407; // @[sm_x105_inr_Foreach.scala 96:22:@3613.4]
  assign x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_sigsIn_baseEn = _T_395 & _T_404; // @[sm_x105_inr_Foreach.scala 96:22:@3612.4]
  assign x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_sigsIn_break = x105_inr_Foreach_sm_io_break; // @[sm_x105_inr_Foreach.scala 96:22:@3611.4]
  assign x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = x99_ctrchain_io_output_counts_0; // @[sm_x105_inr_Foreach.scala 96:22:@3606.4]
  assign x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x99_ctrchain_io_output_oobs_0; // @[sm_x105_inr_Foreach.scala 96:22:@3605.4]
  assign x105_inr_Foreach_kernelx105_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x105_inr_Foreach.scala 95:18:@3601.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_315 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_315 <= 1'h0;
    end else begin
      _T_315 <= _T_312;
    end
  end
endmodule
module RetimeWrapper_36( // @[:@4257.2]
  input   clock, // @[:@4258.4]
  input   reset, // @[:@4259.4]
  input   io_flow, // @[:@4260.4]
  input   io_in, // @[:@4260.4]
  output  io_out // @[:@4260.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@4262.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@4262.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@4262.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@4262.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@4262.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@4262.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(4)) sr ( // @[RetimeShiftRegister.scala 15:20:@4262.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@4275.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@4274.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@4273.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@4272.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@4271.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@4269.4]
endmodule
module RetimeWrapper_40( // @[:@4385.2]
  input   clock, // @[:@4386.4]
  input   reset, // @[:@4387.4]
  input   io_flow, // @[:@4388.4]
  input   io_in, // @[:@4388.4]
  output  io_out // @[:@4388.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@4390.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@4390.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@4390.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@4390.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@4390.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@4390.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@4390.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@4403.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@4402.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@4401.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@4400.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@4399.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@4397.4]
endmodule
module x116_inr_Foreach_sm( // @[:@4405.2]
  input   clock, // @[:@4406.4]
  input   reset, // @[:@4407.4]
  input   io_enable, // @[:@4408.4]
  output  io_done, // @[:@4408.4]
  output  io_doneLatch, // @[:@4408.4]
  input   io_ctrDone, // @[:@4408.4]
  output  io_datapathEn, // @[:@4408.4]
  output  io_ctrInc, // @[:@4408.4]
  output  io_ctrRst, // @[:@4408.4]
  input   io_parentAck, // @[:@4408.4]
  input   io_backpressure, // @[:@4408.4]
  input   io_break // @[:@4408.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@4410.4]
  wire  active_reset; // @[Controllers.scala 261:22:@4410.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@4410.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@4410.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@4410.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@4410.4]
  wire  done_clock; // @[Controllers.scala 262:20:@4413.4]
  wire  done_reset; // @[Controllers.scala 262:20:@4413.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@4413.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@4413.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@4413.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@4413.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@4447.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@4447.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@4447.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@4447.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@4447.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@4469.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@4469.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@4469.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@4469.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@4469.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@4481.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@4481.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@4481.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@4481.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@4481.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@4489.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@4489.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@4489.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@4489.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@4489.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@4505.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@4505.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@4505.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@4505.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@4505.4]
  wire  _T_80; // @[Controllers.scala 264:48:@4418.4]
  wire  _T_81; // @[Controllers.scala 264:46:@4419.4]
  wire  _T_82; // @[Controllers.scala 264:62:@4420.4]
  wire  _T_83; // @[Controllers.scala 264:60:@4421.4]
  wire  _T_100; // @[package.scala 100:49:@4438.4]
  reg  _T_103; // @[package.scala 48:56:@4439.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@4452.4 package.scala 96:25:@4453.4]
  wire  _T_110; // @[package.scala 100:49:@4454.4]
  reg  _T_113; // @[package.scala 48:56:@4455.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@4457.4]
  wire  _T_118; // @[Controllers.scala 283:41:@4462.4]
  wire  _T_119; // @[Controllers.scala 283:59:@4463.4]
  wire  _T_121; // @[Controllers.scala 284:37:@4466.4]
  wire  _T_124; // @[package.scala 96:25:@4474.4 package.scala 96:25:@4475.4]
  wire  _T_126; // @[package.scala 100:49:@4476.4]
  reg  _T_129; // @[package.scala 48:56:@4477.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@4499.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@4501.4]
  reg  _T_153; // @[package.scala 48:56:@4502.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@4510.4 package.scala 96:25:@4511.4]
  wire  _T_158; // @[Controllers.scala 292:61:@4512.4]
  wire  _T_159; // @[Controllers.scala 292:24:@4513.4]
  SRFF active ( // @[Controllers.scala 261:22:@4410.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@4413.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_36 RetimeWrapper ( // @[package.scala 93:22:@4447.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_1 ( // @[package.scala 93:22:@4469.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@4481.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@4489.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_40 RetimeWrapper_4 ( // @[package.scala 93:22:@4505.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@4418.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@4419.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@4420.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@4421.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@4438.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@4452.4 package.scala 96:25:@4453.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@4454.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@4457.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@4462.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@4463.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@4466.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@4474.4 package.scala 96:25:@4475.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@4476.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@4501.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@4510.4 package.scala 96:25:@4511.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@4512.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@4513.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@4480.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@4515.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@4465.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@4468.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@4460.4]
  assign active_clock = clock; // @[:@4411.4]
  assign active_reset = reset; // @[:@4412.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@4423.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@4427.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@4428.4]
  assign done_clock = clock; // @[:@4414.4]
  assign done_reset = reset; // @[:@4415.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@4443.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@4436.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@4437.4]
  assign RetimeWrapper_clock = clock; // @[:@4448.4]
  assign RetimeWrapper_reset = reset; // @[:@4449.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@4451.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@4450.4]
  assign RetimeWrapper_1_clock = clock; // @[:@4470.4]
  assign RetimeWrapper_1_reset = reset; // @[:@4471.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@4473.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@4472.4]
  assign RetimeWrapper_2_clock = clock; // @[:@4482.4]
  assign RetimeWrapper_2_reset = reset; // @[:@4483.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@4485.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@4484.4]
  assign RetimeWrapper_3_clock = clock; // @[:@4490.4]
  assign RetimeWrapper_3_reset = reset; // @[:@4491.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@4493.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@4492.4]
  assign RetimeWrapper_4_clock = clock; // @[:@4506.4]
  assign RetimeWrapper_4_reset = reset; // @[:@4507.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@4509.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@4508.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module RetimeWrapper_44( // @[:@4714.2]
  input         clock, // @[:@4715.4]
  input         reset, // @[:@4716.4]
  input         io_flow, // @[:@4717.4]
  input  [31:0] io_in, // @[:@4717.4]
  output [31:0] io_out // @[:@4717.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@4719.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@4719.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@4719.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@4719.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@4719.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@4719.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@4719.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@4732.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@4731.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@4730.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@4729.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@4728.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@4726.4]
endmodule
module fix2fixBox_2( // @[:@4734.2]
  input  [31:0] io_a, // @[:@4737.4]
  output [32:0] io_b // @[:@4737.4]
);
  assign io_b = {1'h0,io_a}; // @[Converter.scala 95:38:@4748.4]
endmodule
module __2( // @[:@4750.2]
  input  [31:0] io_b, // @[:@4753.4]
  output [32:0] io_result // @[:@4753.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@4758.4]
  wire [32:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@4758.4]
  fix2fixBox_2 fix2fixBox ( // @[BigIPZynq.scala 219:30:@4758.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 706:17:@4766.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@4761.4]
endmodule
module fix2fixBox_4( // @[:@4834.2]
  input         clock, // @[:@4835.4]
  input         reset, // @[:@4836.4]
  input  [32:0] io_a, // @[:@4837.4]
  input         io_flow, // @[:@4837.4]
  output [31:0] io_b // @[:@4837.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@4847.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@4847.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@4847.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@4847.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@4847.4]
  RetimeWrapper_33 RetimeWrapper ( // @[package.scala 93:22:@4847.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@4854.4]
  assign RetimeWrapper_clock = clock; // @[:@4848.4]
  assign RetimeWrapper_reset = reset; // @[:@4849.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@4851.4]
  assign RetimeWrapper_io_in = io_a[31:0]; // @[package.scala 94:16:@4850.4]
endmodule
module x114_sum( // @[:@4856.2]
  input         clock, // @[:@4857.4]
  input         reset, // @[:@4858.4]
  input  [31:0] io_a, // @[:@4859.4]
  input         io_flow, // @[:@4859.4]
  output [31:0] io_result // @[:@4859.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@4867.4]
  wire [32:0] __io_result; // @[Math.scala 709:24:@4867.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@4874.4]
  wire [32:0] __1_io_result; // @[Math.scala 709:24:@4874.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@4884.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@4884.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@4884.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@4884.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@4884.4]
  wire [32:0] a_upcast_number; // @[Math.scala 712:22:@4872.4 Math.scala 713:14:@4873.4]
  wire [32:0] b_upcast_number; // @[Math.scala 712:22:@4879.4 Math.scala 713:14:@4880.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@4881.4]
  __2 _ ( // @[Math.scala 709:24:@4867.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 709:24:@4874.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_4 fix2fixBox ( // @[Math.scala 141:30:@4884.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@4872.4 Math.scala 713:14:@4873.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@4879.4 Math.scala 713:14:@4880.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@4881.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@4892.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@4870.4]
  assign __1_io_b = 32'h5; // @[Math.scala 710:17:@4877.4]
  assign fix2fixBox_clock = clock; // @[:@4885.4]
  assign fix2fixBox_reset = reset; // @[:@4886.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@4887.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@4890.4]
endmodule
module x116_inr_Foreach_kernelx116_inr_Foreach_concrete1( // @[:@4958.2]
  input         clock, // @[:@4959.4]
  input         reset, // @[:@4960.4]
  output        io_in_x97_a_0_rPort_0_en_0, // @[:@4961.4]
  input  [31:0] io_in_x97_a_0_rPort_0_output_0, // @[:@4961.4]
  input         io_in_x97_a_0_empty, // @[:@4961.4]
  input         io_in_x97_a_0_accessActivesOut_1, // @[:@4961.4]
  output        io_in_x97_a_0_accessActivesIn_1, // @[:@4961.4]
  output [31:0] io_in_x107_b_0_wPort_0_data_0, // @[:@4961.4]
  output        io_in_x107_b_0_wPort_0_en_0, // @[:@4961.4]
  input         io_in_x107_b_0_full, // @[:@4961.4]
  input         io_in_x107_b_0_accessActivesOut_0, // @[:@4961.4]
  output        io_in_x107_b_0_accessActivesIn_0, // @[:@4961.4]
  output [63:0] io_in_instrctrs_4_cycs, // @[:@4961.4]
  output [63:0] io_in_instrctrs_4_iters, // @[:@4961.4]
  output [63:0] io_in_instrctrs_4_stalls, // @[:@4961.4]
  output [63:0] io_in_instrctrs_4_idles, // @[:@4961.4]
  input         io_sigsIn_done, // @[:@4961.4]
  input         io_sigsIn_backpressure, // @[:@4961.4]
  input         io_sigsIn_datapathEn, // @[:@4961.4]
  input         io_sigsIn_baseEn, // @[:@4961.4]
  input         io_sigsIn_break, // @[:@4961.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@4961.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@4961.4]
  input         io_rr // @[:@4961.4]
);
  wire  cycles_clock; // @[sm_x116_inr_Foreach.scala 62:26:@5043.4]
  wire  cycles_reset; // @[sm_x116_inr_Foreach.scala 62:26:@5043.4]
  wire  cycles_io_enable; // @[sm_x116_inr_Foreach.scala 62:26:@5043.4]
  wire [63:0] cycles_io_count; // @[sm_x116_inr_Foreach.scala 62:26:@5043.4]
  wire  iters_clock; // @[sm_x116_inr_Foreach.scala 63:25:@5046.4]
  wire  iters_reset; // @[sm_x116_inr_Foreach.scala 63:25:@5046.4]
  wire  iters_io_enable; // @[sm_x116_inr_Foreach.scala 63:25:@5046.4]
  wire [63:0] iters_io_count; // @[sm_x116_inr_Foreach.scala 63:25:@5046.4]
  wire  stalls_clock; // @[sm_x116_inr_Foreach.scala 66:26:@5055.4]
  wire  stalls_reset; // @[sm_x116_inr_Foreach.scala 66:26:@5055.4]
  wire  stalls_io_enable; // @[sm_x116_inr_Foreach.scala 66:26:@5055.4]
  wire [63:0] stalls_io_count; // @[sm_x116_inr_Foreach.scala 66:26:@5055.4]
  wire  idles_clock; // @[sm_x116_inr_Foreach.scala 67:25:@5058.4]
  wire  idles_reset; // @[sm_x116_inr_Foreach.scala 67:25:@5058.4]
  wire  idles_io_enable; // @[sm_x116_inr_Foreach.scala 67:25:@5058.4]
  wire [63:0] idles_io_count; // @[sm_x116_inr_Foreach.scala 67:25:@5058.4]
  wire [31:0] __io_b; // @[Math.scala 709:24:@5081.4]
  wire [31:0] __io_result; // @[Math.scala 709:24:@5081.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@5104.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@5104.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@5104.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@5104.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@5104.4]
  wire  x114_sum_1_clock; // @[Math.scala 150:24:@5122.4]
  wire  x114_sum_1_reset; // @[Math.scala 150:24:@5122.4]
  wire [31:0] x114_sum_1_io_a; // @[Math.scala 150:24:@5122.4]
  wire  x114_sum_1_io_flow; // @[Math.scala 150:24:@5122.4]
  wire [31:0] x114_sum_1_io_result; // @[Math.scala 150:24:@5122.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@5132.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@5132.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@5132.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@5132.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@5132.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@5143.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@5143.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@5143.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@5143.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@5143.4]
  wire  _T_464; // @[package.scala 100:49:@5050.4]
  reg  _T_467; // @[package.scala 48:56:@5051.4]
  reg [31:0] _RAND_0;
  wire  _T_469; // @[sm_x116_inr_Foreach.scala 68:49:@5061.4]
  wire  _T_470; // @[sm_x116_inr_Foreach.scala 68:66:@5062.4]
  wire  _T_471; // @[sm_x116_inr_Foreach.scala 68:64:@5063.4]
  wire  _T_472; // @[sm_x116_inr_Foreach.scala 68:46:@5064.4]
  wire  _T_474; // @[sm_x116_inr_Foreach.scala 69:48:@5067.4]
  wire  _T_475; // @[sm_x116_inr_Foreach.scala 69:65:@5068.4]
  wire  _T_476; // @[sm_x116_inr_Foreach.scala 69:63:@5069.4]
  wire  _T_477; // @[sm_x116_inr_Foreach.scala 69:45:@5070.4]
  wire  b111; // @[sm_x116_inr_Foreach.scala 72:18:@5089.4]
  wire  _T_492; // @[sm_x116_inr_Foreach.scala 77:143:@5091.4]
  wire  _T_496; // @[implicits.scala 55:10:@5094.4]
  wire  _T_497; // @[sm_x116_inr_Foreach.scala 77:160:@5095.4]
  wire  _T_530; // @[package.scala 96:25:@5148.4 package.scala 96:25:@5149.4]
  wire  _T_532; // @[implicits.scala 55:10:@5150.4]
  wire  _T_533; // @[sm_x116_inr_Foreach.scala 93:137:@5151.4]
  wire  _T_535; // @[sm_x116_inr_Foreach.scala 93:224:@5153.4]
  wire  _T_536; // @[sm_x116_inr_Foreach.scala 93:243:@5154.4]
  wire  x169_b111_D3; // @[package.scala 96:25:@5137.4 package.scala 96:25:@5138.4]
  InstrumentationCounter cycles ( // @[sm_x116_inr_Foreach.scala 62:26:@5043.4]
    .clock(cycles_clock),
    .reset(cycles_reset),
    .io_enable(cycles_io_enable),
    .io_count(cycles_io_count)
  );
  InstrumentationCounter iters ( // @[sm_x116_inr_Foreach.scala 63:25:@5046.4]
    .clock(iters_clock),
    .reset(iters_reset),
    .io_enable(iters_io_enable),
    .io_count(iters_io_count)
  );
  InstrumentationCounter stalls ( // @[sm_x116_inr_Foreach.scala 66:26:@5055.4]
    .clock(stalls_clock),
    .reset(stalls_reset),
    .io_enable(stalls_io_enable),
    .io_count(stalls_io_count)
  );
  InstrumentationCounter idles ( // @[sm_x116_inr_Foreach.scala 67:25:@5058.4]
    .clock(idles_clock),
    .reset(idles_reset),
    .io_enable(idles_io_enable),
    .io_count(idles_io_count)
  );
  _ _ ( // @[Math.scala 709:24:@5081.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  RetimeWrapper_44 RetimeWrapper ( // @[package.scala 93:22:@5104.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x114_sum x114_sum_1 ( // @[Math.scala 150:24:@5122.4]
    .clock(x114_sum_1_clock),
    .reset(x114_sum_1_reset),
    .io_a(x114_sum_1_io_a),
    .io_flow(x114_sum_1_io_flow),
    .io_result(x114_sum_1_io_result)
  );
  RetimeWrapper_40 RetimeWrapper_1 ( // @[package.scala 93:22:@5132.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_40 RetimeWrapper_2 ( // @[package.scala 93:22:@5143.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  assign _T_464 = io_sigsIn_done == 1'h0; // @[package.scala 100:49:@5050.4]
  assign _T_469 = ~ io_in_x107_b_0_full; // @[sm_x116_inr_Foreach.scala 68:49:@5061.4]
  assign _T_470 = ~ io_in_x107_b_0_accessActivesOut_0; // @[sm_x116_inr_Foreach.scala 68:66:@5062.4]
  assign _T_471 = _T_469 | _T_470; // @[sm_x116_inr_Foreach.scala 68:64:@5063.4]
  assign _T_472 = ~ _T_471; // @[sm_x116_inr_Foreach.scala 68:46:@5064.4]
  assign _T_474 = ~ io_in_x97_a_0_empty; // @[sm_x116_inr_Foreach.scala 69:48:@5067.4]
  assign _T_475 = ~ io_in_x97_a_0_accessActivesOut_1; // @[sm_x116_inr_Foreach.scala 69:65:@5068.4]
  assign _T_476 = _T_474 | _T_475; // @[sm_x116_inr_Foreach.scala 69:63:@5069.4]
  assign _T_477 = ~ _T_476; // @[sm_x116_inr_Foreach.scala 69:45:@5070.4]
  assign b111 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x116_inr_Foreach.scala 72:18:@5089.4]
  assign _T_492 = ~ io_sigsIn_break; // @[sm_x116_inr_Foreach.scala 77:143:@5091.4]
  assign _T_496 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 55:10:@5094.4]
  assign _T_497 = _T_492 & _T_496; // @[sm_x116_inr_Foreach.scala 77:160:@5095.4]
  assign _T_530 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@5148.4 package.scala 96:25:@5149.4]
  assign _T_532 = io_rr ? _T_530 : 1'h0; // @[implicits.scala 55:10:@5150.4]
  assign _T_533 = _T_492 & _T_532; // @[sm_x116_inr_Foreach.scala 93:137:@5151.4]
  assign _T_535 = _T_533 & _T_492; // @[sm_x116_inr_Foreach.scala 93:224:@5153.4]
  assign _T_536 = _T_535 & io_sigsIn_backpressure; // @[sm_x116_inr_Foreach.scala 93:243:@5154.4]
  assign x169_b111_D3 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@5137.4 package.scala 96:25:@5138.4]
  assign io_in_x97_a_0_rPort_0_en_0 = _T_497 & b111; // @[MemInterfaceType.scala 110:79:@5099.4]
  assign io_in_x97_a_0_accessActivesIn_1 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[MemInterfaceType.scala 148:24:@5102.4]
  assign io_in_x107_b_0_wPort_0_data_0 = x114_sum_1_io_result; // @[MemInterfaceType.scala 90:56:@5157.4]
  assign io_in_x107_b_0_wPort_0_en_0 = _T_536 & x169_b111_D3; // @[MemInterfaceType.scala 93:57:@5159.4]
  assign io_in_x107_b_0_accessActivesIn_0 = RetimeWrapper_1_io_out; // @[MemInterfaceType.scala 148:24:@5161.4]
  assign io_in_instrctrs_4_cycs = cycles_io_count; // @[Ledger.scala 282:21:@5073.4]
  assign io_in_instrctrs_4_iters = iters_io_count; // @[Ledger.scala 283:22:@5074.4]
  assign io_in_instrctrs_4_stalls = stalls_io_count; // @[Ledger.scala 284:23:@5075.4]
  assign io_in_instrctrs_4_idles = idles_io_count; // @[Ledger.scala 285:22:@5076.4]
  assign cycles_clock = clock; // @[:@5044.4]
  assign cycles_reset = reset; // @[:@5045.4]
  assign cycles_io_enable = io_sigsIn_baseEn; // @[sm_x116_inr_Foreach.scala 64:24:@5049.4]
  assign iters_clock = clock; // @[:@5047.4]
  assign iters_reset = reset; // @[:@5048.4]
  assign iters_io_enable = io_sigsIn_done & _T_467; // @[sm_x116_inr_Foreach.scala 65:23:@5054.4]
  assign stalls_clock = clock; // @[:@5056.4]
  assign stalls_reset = reset; // @[:@5057.4]
  assign stalls_io_enable = io_sigsIn_baseEn & _T_472; // @[sm_x116_inr_Foreach.scala 68:24:@5066.4]
  assign idles_clock = clock; // @[:@5059.4]
  assign idles_reset = reset; // @[:@5060.4]
  assign idles_io_enable = io_sigsIn_baseEn & _T_477; // @[sm_x116_inr_Foreach.scala 69:23:@5072.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 710:17:@5084.4]
  assign RetimeWrapper_clock = clock; // @[:@5105.4]
  assign RetimeWrapper_reset = reset; // @[:@5106.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@5108.4]
  assign RetimeWrapper_io_in = io_in_x97_a_0_rPort_0_output_0; // @[package.scala 94:16:@5107.4]
  assign x114_sum_1_clock = clock; // @[:@5123.4]
  assign x114_sum_1_reset = reset; // @[:@5124.4]
  assign x114_sum_1_io_a = RetimeWrapper_io_out; // @[Math.scala 151:17:@5125.4]
  assign x114_sum_1_io_flow = _T_469 | _T_470; // @[Math.scala 153:20:@5127.4]
  assign RetimeWrapper_1_clock = clock; // @[:@5133.4]
  assign RetimeWrapper_1_reset = reset; // @[:@5134.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@5136.4]
  assign RetimeWrapper_1_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@5135.4]
  assign RetimeWrapper_2_clock = clock; // @[:@5144.4]
  assign RetimeWrapper_2_reset = reset; // @[:@5145.4]
  assign RetimeWrapper_2_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@5147.4]
  assign RetimeWrapper_2_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@5146.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_467 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_467 <= 1'h0;
    end else begin
      _T_467 <= _T_464;
    end
  end
endmodule
module x130_inr_Foreach_kernelx130_inr_Foreach_concrete1( // @[:@6424.2]
  input         clock, // @[:@6425.4]
  input         reset, // @[:@6426.4]
  output        io_in_x95_TVALID, // @[:@6427.4]
  input         io_in_x95_TREADY, // @[:@6427.4]
  output [63:0] io_in_x95_TDATA, // @[:@6427.4]
  output [7:0]  io_in_x95_TSTRB, // @[:@6427.4]
  output [7:0]  io_in_x95_TKEEP, // @[:@6427.4]
  output        io_in_x95_TLAST, // @[:@6427.4]
  output [7:0]  io_in_x95_TID, // @[:@6427.4]
  output [7:0]  io_in_x95_TDEST, // @[:@6427.4]
  output [31:0] io_in_x95_TUSER, // @[:@6427.4]
  output        io_in_x107_b_0_rPort_0_en_0, // @[:@6427.4]
  input  [31:0] io_in_x107_b_0_rPort_0_output_0, // @[:@6427.4]
  input         io_in_x107_b_0_empty, // @[:@6427.4]
  input         io_in_x107_b_0_accessActivesOut_1, // @[:@6427.4]
  output        io_in_x107_b_0_accessActivesIn_1, // @[:@6427.4]
  output [63:0] io_in_instrctrs_6_cycs, // @[:@6427.4]
  output [63:0] io_in_instrctrs_6_iters, // @[:@6427.4]
  output [63:0] io_in_instrctrs_6_stalls, // @[:@6427.4]
  output [63:0] io_in_instrctrs_6_idles, // @[:@6427.4]
  input         io_sigsIn_done, // @[:@6427.4]
  input         io_sigsIn_backpressure, // @[:@6427.4]
  input         io_sigsIn_datapathEn, // @[:@6427.4]
  input         io_sigsIn_baseEn, // @[:@6427.4]
  input         io_sigsIn_break, // @[:@6427.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@6427.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@6427.4]
  input         io_rr // @[:@6427.4]
);
  wire  cycles_clock; // @[sm_x130_inr_Foreach.scala 63:26:@6487.4]
  wire  cycles_reset; // @[sm_x130_inr_Foreach.scala 63:26:@6487.4]
  wire  cycles_io_enable; // @[sm_x130_inr_Foreach.scala 63:26:@6487.4]
  wire [63:0] cycles_io_count; // @[sm_x130_inr_Foreach.scala 63:26:@6487.4]
  wire  iters_clock; // @[sm_x130_inr_Foreach.scala 64:25:@6490.4]
  wire  iters_reset; // @[sm_x130_inr_Foreach.scala 64:25:@6490.4]
  wire  iters_io_enable; // @[sm_x130_inr_Foreach.scala 64:25:@6490.4]
  wire [63:0] iters_io_count; // @[sm_x130_inr_Foreach.scala 64:25:@6490.4]
  wire  stalls_clock; // @[sm_x130_inr_Foreach.scala 67:26:@6499.4]
  wire  stalls_reset; // @[sm_x130_inr_Foreach.scala 67:26:@6499.4]
  wire  stalls_io_enable; // @[sm_x130_inr_Foreach.scala 67:26:@6499.4]
  wire [63:0] stalls_io_count; // @[sm_x130_inr_Foreach.scala 67:26:@6499.4]
  wire  idles_clock; // @[sm_x130_inr_Foreach.scala 68:25:@6502.4]
  wire  idles_reset; // @[sm_x130_inr_Foreach.scala 68:25:@6502.4]
  wire  idles_io_enable; // @[sm_x130_inr_Foreach.scala 68:25:@6502.4]
  wire [63:0] idles_io_count; // @[sm_x130_inr_Foreach.scala 68:25:@6502.4]
  wire [31:0] __io_b; // @[Math.scala 709:24:@6522.4]
  wire [31:0] __io_result; // @[Math.scala 709:24:@6522.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@6559.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@6559.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@6559.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@6559.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@6559.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@6675.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@6675.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@6675.4]
  wire [31:0] RetimeWrapper_1_io_in; // @[package.scala 93:22:@6675.4]
  wire [31:0] RetimeWrapper_1_io_out; // @[package.scala 93:22:@6675.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@6684.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@6684.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@6684.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@6684.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@6684.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@6709.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@6709.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@6709.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@6709.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@6709.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@6718.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@6718.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@6718.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@6718.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@6718.4]
  wire  _T_332; // @[package.scala 100:49:@6494.4]
  reg  _T_335; // @[package.scala 48:56:@6495.4]
  reg [31:0] _RAND_0;
  wire  _T_337; // @[sm_x130_inr_Foreach.scala 69:46:@6505.4]
  wire  _T_339; // @[sm_x130_inr_Foreach.scala 70:48:@6508.4]
  wire  _T_340; // @[sm_x130_inr_Foreach.scala 70:66:@6509.4]
  wire  _T_341; // @[sm_x130_inr_Foreach.scala 70:64:@6510.4]
  wire  _T_342; // @[sm_x130_inr_Foreach.scala 70:45:@6511.4]
  wire  b120; // @[sm_x130_inr_Foreach.scala 73:18:@6530.4]
  wire [31:0] b119_number; // @[Math.scala 712:22:@6527.4 Math.scala 713:14:@6528.4]
  wire [31:0] _T_357; // @[Math.scala 499:37:@6536.4]
  wire  x121; // @[Math.scala 499:44:@6538.4]
  wire  _T_376; // @[sm_x130_inr_Foreach.scala 84:148:@6548.4]
  wire  _T_380; // @[implicits.scala 55:10:@6551.4]
  wire  _T_381; // @[sm_x130_inr_Foreach.scala 84:165:@6552.4]
  wire [31:0] x170_x123_deq_x107_D2_0_number; // @[package.scala 96:25:@6564.4 package.scala 96:25:@6565.4]
  wire  x126_0; // @[FixedPoint.scala 19:42:@6577.4]
  wire  x126_1; // @[FixedPoint.scala 19:42:@6579.4]
  wire  x126_2; // @[FixedPoint.scala 19:42:@6581.4]
  wire  x126_3; // @[FixedPoint.scala 19:42:@6583.4]
  wire  x126_4; // @[FixedPoint.scala 19:42:@6585.4]
  wire  x126_5; // @[FixedPoint.scala 19:42:@6587.4]
  wire  x126_6; // @[FixedPoint.scala 19:42:@6589.4]
  wire  x126_7; // @[FixedPoint.scala 19:42:@6591.4]
  wire  x126_8; // @[FixedPoint.scala 19:42:@6593.4]
  wire  x126_9; // @[FixedPoint.scala 19:42:@6595.4]
  wire  x126_10; // @[FixedPoint.scala 19:42:@6597.4]
  wire  x126_11; // @[FixedPoint.scala 19:42:@6599.4]
  wire  x126_12; // @[FixedPoint.scala 19:42:@6601.4]
  wire  x126_13; // @[FixedPoint.scala 19:42:@6603.4]
  wire  x126_14; // @[FixedPoint.scala 19:42:@6605.4]
  wire  x126_15; // @[FixedPoint.scala 19:42:@6607.4]
  wire  x126_16; // @[FixedPoint.scala 19:42:@6609.4]
  wire  x126_17; // @[FixedPoint.scala 19:42:@6611.4]
  wire  x126_18; // @[FixedPoint.scala 19:42:@6613.4]
  wire  x126_19; // @[FixedPoint.scala 19:42:@6615.4]
  wire  x126_20; // @[FixedPoint.scala 19:42:@6617.4]
  wire  x126_21; // @[FixedPoint.scala 19:42:@6619.4]
  wire  x126_22; // @[FixedPoint.scala 19:42:@6621.4]
  wire  x126_23; // @[FixedPoint.scala 19:42:@6623.4]
  wire  x126_24; // @[FixedPoint.scala 19:42:@6625.4]
  wire  x126_25; // @[FixedPoint.scala 19:42:@6627.4]
  wire  x126_26; // @[FixedPoint.scala 19:42:@6629.4]
  wire  x126_27; // @[FixedPoint.scala 19:42:@6631.4]
  wire  x126_28; // @[FixedPoint.scala 19:42:@6633.4]
  wire  x126_29; // @[FixedPoint.scala 19:42:@6635.4]
  wire  x126_30; // @[FixedPoint.scala 19:42:@6637.4]
  wire  x126_31; // @[FixedPoint.scala 19:42:@6639.4]
  wire [7:0] _T_476; // @[Cat.scala 30:58:@6648.4]
  wire [15:0] _T_484; // @[Cat.scala 30:58:@6656.4]
  wire [7:0] _T_491; // @[Cat.scala 30:58:@6663.4]
  wire [31:0] _T_500; // @[Cat.scala 30:58:@6672.4]
  wire [63:0] x127_number; // @[sm_x130_inr_Foreach.scala 94:22:@6641.4 sm_x130_inr_Foreach.scala 95:14:@6673.4]
  wire  x172_x125_D2; // @[package.scala 96:25:@6689.4 package.scala 96:25:@6690.4]
  wire [31:0] x171_x122_D2_number; // @[package.scala 96:25:@6680.4 package.scala 96:25:@6681.4]
  wire [128:0] x128_tuple; // @[Cat.scala 30:58:@6706.4]
  wire  _T_535; // @[package.scala 96:25:@6723.4 package.scala 96:25:@6724.4]
  wire  _T_537; // @[implicits.scala 55:10:@6725.4]
  wire  x173_b120_D2; // @[package.scala 96:25:@6714.4 package.scala 96:25:@6715.4]
  wire  _T_538; // @[sm_x130_inr_Foreach.scala 104:110:@6726.4]
  InstrumentationCounter cycles ( // @[sm_x130_inr_Foreach.scala 63:26:@6487.4]
    .clock(cycles_clock),
    .reset(cycles_reset),
    .io_enable(cycles_io_enable),
    .io_count(cycles_io_count)
  );
  InstrumentationCounter iters ( // @[sm_x130_inr_Foreach.scala 64:25:@6490.4]
    .clock(iters_clock),
    .reset(iters_reset),
    .io_enable(iters_io_enable),
    .io_count(iters_io_count)
  );
  InstrumentationCounter stalls ( // @[sm_x130_inr_Foreach.scala 67:26:@6499.4]
    .clock(stalls_clock),
    .reset(stalls_reset),
    .io_enable(stalls_io_enable),
    .io_count(stalls_io_count)
  );
  InstrumentationCounter idles ( // @[sm_x130_inr_Foreach.scala 68:25:@6502.4]
    .clock(idles_clock),
    .reset(idles_reset),
    .io_enable(idles_io_enable),
    .io_count(idles_io_count)
  );
  _ _ ( // @[Math.scala 709:24:@6522.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  RetimeWrapper_44 RetimeWrapper ( // @[package.scala 93:22:@6559.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_1 ( // @[package.scala 93:22:@6675.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_2 ( // @[package.scala 93:22:@6684.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_3 ( // @[package.scala 93:22:@6709.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_4 ( // @[package.scala 93:22:@6718.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_332 = io_sigsIn_done == 1'h0; // @[package.scala 100:49:@6494.4]
  assign _T_337 = ~ io_in_x95_TREADY; // @[sm_x130_inr_Foreach.scala 69:46:@6505.4]
  assign _T_339 = ~ io_in_x107_b_0_empty; // @[sm_x130_inr_Foreach.scala 70:48:@6508.4]
  assign _T_340 = ~ io_in_x107_b_0_accessActivesOut_1; // @[sm_x130_inr_Foreach.scala 70:66:@6509.4]
  assign _T_341 = _T_339 | _T_340; // @[sm_x130_inr_Foreach.scala 70:64:@6510.4]
  assign _T_342 = ~ _T_341; // @[sm_x130_inr_Foreach.scala 70:45:@6511.4]
  assign b120 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x130_inr_Foreach.scala 73:18:@6530.4]
  assign b119_number = __io_result; // @[Math.scala 712:22:@6527.4 Math.scala 713:14:@6528.4]
  assign _T_357 = $signed(b119_number); // @[Math.scala 499:37:@6536.4]
  assign x121 = $signed(_T_357) == $signed(32'sh0); // @[Math.scala 499:44:@6538.4]
  assign _T_376 = ~ io_sigsIn_break; // @[sm_x130_inr_Foreach.scala 84:148:@6548.4]
  assign _T_380 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 55:10:@6551.4]
  assign _T_381 = _T_376 & _T_380; // @[sm_x130_inr_Foreach.scala 84:165:@6552.4]
  assign x170_x123_deq_x107_D2_0_number = RetimeWrapper_io_out; // @[package.scala 96:25:@6564.4 package.scala 96:25:@6565.4]
  assign x126_0 = x170_x123_deq_x107_D2_0_number[0]; // @[FixedPoint.scala 19:42:@6577.4]
  assign x126_1 = x170_x123_deq_x107_D2_0_number[1]; // @[FixedPoint.scala 19:42:@6579.4]
  assign x126_2 = x170_x123_deq_x107_D2_0_number[2]; // @[FixedPoint.scala 19:42:@6581.4]
  assign x126_3 = x170_x123_deq_x107_D2_0_number[3]; // @[FixedPoint.scala 19:42:@6583.4]
  assign x126_4 = x170_x123_deq_x107_D2_0_number[4]; // @[FixedPoint.scala 19:42:@6585.4]
  assign x126_5 = x170_x123_deq_x107_D2_0_number[5]; // @[FixedPoint.scala 19:42:@6587.4]
  assign x126_6 = x170_x123_deq_x107_D2_0_number[6]; // @[FixedPoint.scala 19:42:@6589.4]
  assign x126_7 = x170_x123_deq_x107_D2_0_number[7]; // @[FixedPoint.scala 19:42:@6591.4]
  assign x126_8 = x170_x123_deq_x107_D2_0_number[8]; // @[FixedPoint.scala 19:42:@6593.4]
  assign x126_9 = x170_x123_deq_x107_D2_0_number[9]; // @[FixedPoint.scala 19:42:@6595.4]
  assign x126_10 = x170_x123_deq_x107_D2_0_number[10]; // @[FixedPoint.scala 19:42:@6597.4]
  assign x126_11 = x170_x123_deq_x107_D2_0_number[11]; // @[FixedPoint.scala 19:42:@6599.4]
  assign x126_12 = x170_x123_deq_x107_D2_0_number[12]; // @[FixedPoint.scala 19:42:@6601.4]
  assign x126_13 = x170_x123_deq_x107_D2_0_number[13]; // @[FixedPoint.scala 19:42:@6603.4]
  assign x126_14 = x170_x123_deq_x107_D2_0_number[14]; // @[FixedPoint.scala 19:42:@6605.4]
  assign x126_15 = x170_x123_deq_x107_D2_0_number[15]; // @[FixedPoint.scala 19:42:@6607.4]
  assign x126_16 = x170_x123_deq_x107_D2_0_number[16]; // @[FixedPoint.scala 19:42:@6609.4]
  assign x126_17 = x170_x123_deq_x107_D2_0_number[17]; // @[FixedPoint.scala 19:42:@6611.4]
  assign x126_18 = x170_x123_deq_x107_D2_0_number[18]; // @[FixedPoint.scala 19:42:@6613.4]
  assign x126_19 = x170_x123_deq_x107_D2_0_number[19]; // @[FixedPoint.scala 19:42:@6615.4]
  assign x126_20 = x170_x123_deq_x107_D2_0_number[20]; // @[FixedPoint.scala 19:42:@6617.4]
  assign x126_21 = x170_x123_deq_x107_D2_0_number[21]; // @[FixedPoint.scala 19:42:@6619.4]
  assign x126_22 = x170_x123_deq_x107_D2_0_number[22]; // @[FixedPoint.scala 19:42:@6621.4]
  assign x126_23 = x170_x123_deq_x107_D2_0_number[23]; // @[FixedPoint.scala 19:42:@6623.4]
  assign x126_24 = x170_x123_deq_x107_D2_0_number[24]; // @[FixedPoint.scala 19:42:@6625.4]
  assign x126_25 = x170_x123_deq_x107_D2_0_number[25]; // @[FixedPoint.scala 19:42:@6627.4]
  assign x126_26 = x170_x123_deq_x107_D2_0_number[26]; // @[FixedPoint.scala 19:42:@6629.4]
  assign x126_27 = x170_x123_deq_x107_D2_0_number[27]; // @[FixedPoint.scala 19:42:@6631.4]
  assign x126_28 = x170_x123_deq_x107_D2_0_number[28]; // @[FixedPoint.scala 19:42:@6633.4]
  assign x126_29 = x170_x123_deq_x107_D2_0_number[29]; // @[FixedPoint.scala 19:42:@6635.4]
  assign x126_30 = x170_x123_deq_x107_D2_0_number[30]; // @[FixedPoint.scala 19:42:@6637.4]
  assign x126_31 = x170_x123_deq_x107_D2_0_number[31]; // @[FixedPoint.scala 19:42:@6639.4]
  assign _T_476 = {x126_7,x126_6,x126_5,x126_4,x126_3,x126_2,x126_1,x126_0}; // @[Cat.scala 30:58:@6648.4]
  assign _T_484 = {x126_15,x126_14,x126_13,x126_12,x126_11,x126_10,x126_9,x126_8,_T_476}; // @[Cat.scala 30:58:@6656.4]
  assign _T_491 = {x126_23,x126_22,x126_21,x126_20,x126_19,x126_18,x126_17,x126_16}; // @[Cat.scala 30:58:@6663.4]
  assign _T_500 = {x126_31,x126_30,x126_29,x126_28,x126_27,x126_26,x126_25,x126_24,_T_491,_T_484}; // @[Cat.scala 30:58:@6672.4]
  assign x127_number = {{32'd0}, _T_500}; // @[sm_x130_inr_Foreach.scala 94:22:@6641.4 sm_x130_inr_Foreach.scala 95:14:@6673.4]
  assign x172_x125_D2 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@6689.4 package.scala 96:25:@6690.4]
  assign x171_x122_D2_number = RetimeWrapper_1_io_out; // @[package.scala 96:25:@6680.4 package.scala 96:25:@6681.4]
  assign x128_tuple = {x171_x122_D2_number,8'h1,8'h0,x172_x125_D2,16'h0,x127_number}; // @[Cat.scala 30:58:@6706.4]
  assign _T_535 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@6723.4 package.scala 96:25:@6724.4]
  assign _T_537 = io_rr ? _T_535 : 1'h0; // @[implicits.scala 55:10:@6725.4]
  assign x173_b120_D2 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@6714.4 package.scala 96:25:@6715.4]
  assign _T_538 = _T_537 & x173_b120_D2; // @[sm_x130_inr_Foreach.scala 104:110:@6726.4]
  assign io_in_x95_TVALID = _T_538 & io_sigsIn_backpressure; // @[sm_x130_inr_Foreach.scala 104:17:@6728.4]
  assign io_in_x95_TDATA = x128_tuple[63:0]; // @[sm_x130_inr_Foreach.scala 105:19:@6730.4]
  assign io_in_x95_TSTRB = x128_tuple[71:64]; // @[sm_x130_inr_Foreach.scala 106:19:@6732.4]
  assign io_in_x95_TKEEP = x128_tuple[79:72]; // @[sm_x130_inr_Foreach.scala 107:19:@6734.4]
  assign io_in_x95_TLAST = x128_tuple[80]; // @[sm_x130_inr_Foreach.scala 110:17:@6740.4]
  assign io_in_x95_TID = x128_tuple[88:81]; // @[sm_x130_inr_Foreach.scala 108:17:@6736.4]
  assign io_in_x95_TDEST = x128_tuple[96:89]; // @[sm_x130_inr_Foreach.scala 109:19:@6738.4]
  assign io_in_x95_TUSER = x128_tuple[128:97]; // @[sm_x130_inr_Foreach.scala 111:17:@6742.4]
  assign io_in_x107_b_0_rPort_0_en_0 = _T_381 & b120; // @[MemInterfaceType.scala 110:79:@6555.4]
  assign io_in_x107_b_0_accessActivesIn_1 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[MemInterfaceType.scala 148:24:@6557.4]
  assign io_in_instrctrs_6_cycs = cycles_io_count; // @[Ledger.scala 282:21:@6514.4]
  assign io_in_instrctrs_6_iters = iters_io_count; // @[Ledger.scala 283:22:@6515.4]
  assign io_in_instrctrs_6_stalls = stalls_io_count; // @[Ledger.scala 284:23:@6516.4]
  assign io_in_instrctrs_6_idles = idles_io_count; // @[Ledger.scala 285:22:@6517.4]
  assign cycles_clock = clock; // @[:@6488.4]
  assign cycles_reset = reset; // @[:@6489.4]
  assign cycles_io_enable = io_sigsIn_baseEn; // @[sm_x130_inr_Foreach.scala 65:24:@6493.4]
  assign iters_clock = clock; // @[:@6491.4]
  assign iters_reset = reset; // @[:@6492.4]
  assign iters_io_enable = io_sigsIn_done & _T_335; // @[sm_x130_inr_Foreach.scala 66:23:@6498.4]
  assign stalls_clock = clock; // @[:@6500.4]
  assign stalls_reset = reset; // @[:@6501.4]
  assign stalls_io_enable = io_sigsIn_baseEn & _T_337; // @[sm_x130_inr_Foreach.scala 69:24:@6507.4]
  assign idles_clock = clock; // @[:@6503.4]
  assign idles_reset = reset; // @[:@6504.4]
  assign idles_io_enable = io_sigsIn_baseEn & _T_342; // @[sm_x130_inr_Foreach.scala 70:23:@6513.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 710:17:@6525.4]
  assign RetimeWrapper_clock = clock; // @[:@6560.4]
  assign RetimeWrapper_reset = reset; // @[:@6561.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@6563.4]
  assign RetimeWrapper_io_in = io_in_x107_b_0_rPort_0_output_0; // @[package.scala 94:16:@6562.4]
  assign RetimeWrapper_1_clock = clock; // @[:@6676.4]
  assign RetimeWrapper_1_reset = reset; // @[:@6677.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@6679.4]
  assign RetimeWrapper_1_io_in = x121 ? 32'h2 : 32'h0; // @[package.scala 94:16:@6678.4]
  assign RetimeWrapper_2_clock = clock; // @[:@6685.4]
  assign RetimeWrapper_2_reset = reset; // @[:@6686.4]
  assign RetimeWrapper_2_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@6688.4]
  assign RetimeWrapper_2_io_in = $signed(_T_357) == $signed(32'sh3f); // @[package.scala 94:16:@6687.4]
  assign RetimeWrapper_3_clock = clock; // @[:@6710.4]
  assign RetimeWrapper_3_reset = reset; // @[:@6711.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@6713.4]
  assign RetimeWrapper_3_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@6712.4]
  assign RetimeWrapper_4_clock = clock; // @[:@6719.4]
  assign RetimeWrapper_4_reset = reset; // @[:@6720.4]
  assign RetimeWrapper_4_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@6722.4]
  assign RetimeWrapper_4_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@6721.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_335 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_335 <= 1'h0;
    end else begin
      _T_335 <= _T_332;
    end
  end
endmodule
module x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1( // @[:@6744.2]
  input         clock, // @[:@6745.4]
  input         reset, // @[:@6746.4]
  output        io_in_x95_TVALID, // @[:@6747.4]
  input         io_in_x95_TREADY, // @[:@6747.4]
  output [63:0] io_in_x95_TDATA, // @[:@6747.4]
  output [7:0]  io_in_x95_TSTRB, // @[:@6747.4]
  output [7:0]  io_in_x95_TKEEP, // @[:@6747.4]
  output        io_in_x95_TLAST, // @[:@6747.4]
  output [7:0]  io_in_x95_TID, // @[:@6747.4]
  output [7:0]  io_in_x95_TDEST, // @[:@6747.4]
  output [31:0] io_in_x95_TUSER, // @[:@6747.4]
  output        io_in_x107_b_0_rPort_0_en_0, // @[:@6747.4]
  input  [31:0] io_in_x107_b_0_rPort_0_output_0, // @[:@6747.4]
  input         io_in_x107_b_0_empty, // @[:@6747.4]
  input         io_in_x107_b_0_accessActivesOut_1, // @[:@6747.4]
  output        io_in_x107_b_0_accessActivesIn_1, // @[:@6747.4]
  output [63:0] io_in_instrctrs_5_cycs, // @[:@6747.4]
  output [63:0] io_in_instrctrs_5_iters, // @[:@6747.4]
  output [63:0] io_in_instrctrs_6_cycs, // @[:@6747.4]
  output [63:0] io_in_instrctrs_6_iters, // @[:@6747.4]
  output [63:0] io_in_instrctrs_6_stalls, // @[:@6747.4]
  output [63:0] io_in_instrctrs_6_idles, // @[:@6747.4]
  input         io_sigsIn_done, // @[:@6747.4]
  input         io_sigsIn_baseEn, // @[:@6747.4]
  input         io_sigsIn_smEnableOuts_0, // @[:@6747.4]
  input         io_sigsIn_smChildAcks_0, // @[:@6747.4]
  output        io_sigsOut_smDoneIn_0, // @[:@6747.4]
  output        io_sigsOut_smCtrCopyDone_0, // @[:@6747.4]
  input         io_rr // @[:@6747.4]
);
  wire  cycles_clock; // @[sm_x131_outr_UnitPipe.scala 63:26:@6807.4]
  wire  cycles_reset; // @[sm_x131_outr_UnitPipe.scala 63:26:@6807.4]
  wire  cycles_io_enable; // @[sm_x131_outr_UnitPipe.scala 63:26:@6807.4]
  wire [63:0] cycles_io_count; // @[sm_x131_outr_UnitPipe.scala 63:26:@6807.4]
  wire  iters_clock; // @[sm_x131_outr_UnitPipe.scala 64:25:@6810.4]
  wire  iters_reset; // @[sm_x131_outr_UnitPipe.scala 64:25:@6810.4]
  wire  iters_io_enable; // @[sm_x131_outr_UnitPipe.scala 64:25:@6810.4]
  wire [63:0] iters_io_count; // @[sm_x131_outr_UnitPipe.scala 64:25:@6810.4]
  wire  x118_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@6823.4]
  wire  x118_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@6823.4]
  wire  x118_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@6823.4]
  wire  x118_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@6823.4]
  wire [31:0] x118_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@6823.4]
  wire  x118_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@6823.4]
  wire  x118_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@6823.4]
  wire  x130_inr_Foreach_sm_clock; // @[sm_x130_inr_Foreach.scala 33:18:@6875.4]
  wire  x130_inr_Foreach_sm_reset; // @[sm_x130_inr_Foreach.scala 33:18:@6875.4]
  wire  x130_inr_Foreach_sm_io_enable; // @[sm_x130_inr_Foreach.scala 33:18:@6875.4]
  wire  x130_inr_Foreach_sm_io_done; // @[sm_x130_inr_Foreach.scala 33:18:@6875.4]
  wire  x130_inr_Foreach_sm_io_doneLatch; // @[sm_x130_inr_Foreach.scala 33:18:@6875.4]
  wire  x130_inr_Foreach_sm_io_ctrDone; // @[sm_x130_inr_Foreach.scala 33:18:@6875.4]
  wire  x130_inr_Foreach_sm_io_datapathEn; // @[sm_x130_inr_Foreach.scala 33:18:@6875.4]
  wire  x130_inr_Foreach_sm_io_ctrInc; // @[sm_x130_inr_Foreach.scala 33:18:@6875.4]
  wire  x130_inr_Foreach_sm_io_ctrRst; // @[sm_x130_inr_Foreach.scala 33:18:@6875.4]
  wire  x130_inr_Foreach_sm_io_parentAck; // @[sm_x130_inr_Foreach.scala 33:18:@6875.4]
  wire  x130_inr_Foreach_sm_io_backpressure; // @[sm_x130_inr_Foreach.scala 33:18:@6875.4]
  wire  x130_inr_Foreach_sm_io_break; // @[sm_x130_inr_Foreach.scala 33:18:@6875.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@6903.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@6903.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@6903.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@6903.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@6903.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@6946.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@6946.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@6946.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@6946.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@6946.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@6954.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@6954.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@6954.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@6954.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@6954.4]
  wire  x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_clock; // @[sm_x130_inr_Foreach.scala 113:24:@6986.4]
  wire  x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_reset; // @[sm_x130_inr_Foreach.scala 113:24:@6986.4]
  wire  x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_x95_TVALID; // @[sm_x130_inr_Foreach.scala 113:24:@6986.4]
  wire  x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_x95_TREADY; // @[sm_x130_inr_Foreach.scala 113:24:@6986.4]
  wire [63:0] x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_x95_TDATA; // @[sm_x130_inr_Foreach.scala 113:24:@6986.4]
  wire [7:0] x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_x95_TSTRB; // @[sm_x130_inr_Foreach.scala 113:24:@6986.4]
  wire [7:0] x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_x95_TKEEP; // @[sm_x130_inr_Foreach.scala 113:24:@6986.4]
  wire  x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_x95_TLAST; // @[sm_x130_inr_Foreach.scala 113:24:@6986.4]
  wire [7:0] x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_x95_TID; // @[sm_x130_inr_Foreach.scala 113:24:@6986.4]
  wire [7:0] x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_x95_TDEST; // @[sm_x130_inr_Foreach.scala 113:24:@6986.4]
  wire [31:0] x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_x95_TUSER; // @[sm_x130_inr_Foreach.scala 113:24:@6986.4]
  wire  x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_x107_b_0_rPort_0_en_0; // @[sm_x130_inr_Foreach.scala 113:24:@6986.4]
  wire [31:0] x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_x107_b_0_rPort_0_output_0; // @[sm_x130_inr_Foreach.scala 113:24:@6986.4]
  wire  x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_x107_b_0_empty; // @[sm_x130_inr_Foreach.scala 113:24:@6986.4]
  wire  x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_x107_b_0_accessActivesOut_1; // @[sm_x130_inr_Foreach.scala 113:24:@6986.4]
  wire  x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_x107_b_0_accessActivesIn_1; // @[sm_x130_inr_Foreach.scala 113:24:@6986.4]
  wire [63:0] x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_instrctrs_6_cycs; // @[sm_x130_inr_Foreach.scala 113:24:@6986.4]
  wire [63:0] x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_instrctrs_6_iters; // @[sm_x130_inr_Foreach.scala 113:24:@6986.4]
  wire [63:0] x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_instrctrs_6_stalls; // @[sm_x130_inr_Foreach.scala 113:24:@6986.4]
  wire [63:0] x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_instrctrs_6_idles; // @[sm_x130_inr_Foreach.scala 113:24:@6986.4]
  wire  x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_sigsIn_done; // @[sm_x130_inr_Foreach.scala 113:24:@6986.4]
  wire  x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_sigsIn_backpressure; // @[sm_x130_inr_Foreach.scala 113:24:@6986.4]
  wire  x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x130_inr_Foreach.scala 113:24:@6986.4]
  wire  x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_sigsIn_baseEn; // @[sm_x130_inr_Foreach.scala 113:24:@6986.4]
  wire  x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x130_inr_Foreach.scala 113:24:@6986.4]
  wire [31:0] x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x130_inr_Foreach.scala 113:24:@6986.4]
  wire  x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x130_inr_Foreach.scala 113:24:@6986.4]
  wire  x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_rr; // @[sm_x130_inr_Foreach.scala 113:24:@6986.4]
  wire  _T_332; // @[package.scala 100:49:@6814.4]
  reg  _T_335; // @[package.scala 48:56:@6815.4]
  reg [31:0] _RAND_0;
  wire  _T_399; // @[package.scala 96:25:@6908.4 package.scala 96:25:@6909.4]
  wire  _T_403; // @[sm_x131_outr_UnitPipe.scala 75:44:@6914.4]
  wire  _T_404; // @[sm_x131_outr_UnitPipe.scala 75:62:@6915.4]
  wire  _T_405; // @[sm_x131_outr_UnitPipe.scala 75:60:@6916.4]
  wire  x130_inr_Foreach_sigsIn_forwardpressure; // @[sm_x131_outr_UnitPipe.scala 75:95:@6917.4]
  wire  _T_415; // @[package.scala 96:25:@6951.4 package.scala 96:25:@6952.4]
  wire  _T_421; // @[package.scala 96:25:@6959.4 package.scala 96:25:@6960.4]
  wire  _T_424; // @[SpatialBlocks.scala 110:93:@6962.4]
  wire  x130_inr_Foreach_sigsIn_baseEn; // @[SpatialBlocks.scala 110:90:@6963.4]
  wire  _T_426; // @[SpatialBlocks.scala 128:36:@6971.4]
  wire  _T_427; // @[SpatialBlocks.scala 128:78:@6972.4]
  wire  _T_432; // @[SpatialBlocks.scala 130:61:@6981.4]
  InstrumentationCounter cycles ( // @[sm_x131_outr_UnitPipe.scala 63:26:@6807.4]
    .clock(cycles_clock),
    .reset(cycles_reset),
    .io_enable(cycles_io_enable),
    .io_count(cycles_io_count)
  );
  InstrumentationCounter iters ( // @[sm_x131_outr_UnitPipe.scala 64:25:@6810.4]
    .clock(iters_clock),
    .reset(iters_reset),
    .io_enable(iters_io_enable),
    .io_count(iters_io_count)
  );
  x99_ctrchain x118_ctrchain ( // @[SpatialBlocks.scala 37:22:@6823.4]
    .clock(x118_ctrchain_clock),
    .reset(x118_ctrchain_reset),
    .io_input_reset(x118_ctrchain_io_input_reset),
    .io_input_enable(x118_ctrchain_io_input_enable),
    .io_output_counts_0(x118_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x118_ctrchain_io_output_oobs_0),
    .io_output_done(x118_ctrchain_io_output_done)
  );
  x105_inr_Foreach_sm x130_inr_Foreach_sm ( // @[sm_x130_inr_Foreach.scala 33:18:@6875.4]
    .clock(x130_inr_Foreach_sm_clock),
    .reset(x130_inr_Foreach_sm_reset),
    .io_enable(x130_inr_Foreach_sm_io_enable),
    .io_done(x130_inr_Foreach_sm_io_done),
    .io_doneLatch(x130_inr_Foreach_sm_io_doneLatch),
    .io_ctrDone(x130_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x130_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x130_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x130_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x130_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x130_inr_Foreach_sm_io_backpressure),
    .io_break(x130_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@6903.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@6946.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@6954.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x130_inr_Foreach_kernelx130_inr_Foreach_concrete1 x130_inr_Foreach_kernelx130_inr_Foreach_concrete1 ( // @[sm_x130_inr_Foreach.scala 113:24:@6986.4]
    .clock(x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_clock),
    .reset(x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_reset),
    .io_in_x95_TVALID(x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_x95_TVALID),
    .io_in_x95_TREADY(x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_x95_TREADY),
    .io_in_x95_TDATA(x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_x95_TDATA),
    .io_in_x95_TSTRB(x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_x95_TSTRB),
    .io_in_x95_TKEEP(x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_x95_TKEEP),
    .io_in_x95_TLAST(x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_x95_TLAST),
    .io_in_x95_TID(x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_x95_TID),
    .io_in_x95_TDEST(x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_x95_TDEST),
    .io_in_x95_TUSER(x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_x95_TUSER),
    .io_in_x107_b_0_rPort_0_en_0(x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_x107_b_0_rPort_0_en_0),
    .io_in_x107_b_0_rPort_0_output_0(x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_x107_b_0_rPort_0_output_0),
    .io_in_x107_b_0_empty(x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_x107_b_0_empty),
    .io_in_x107_b_0_accessActivesOut_1(x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_x107_b_0_accessActivesOut_1),
    .io_in_x107_b_0_accessActivesIn_1(x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_x107_b_0_accessActivesIn_1),
    .io_in_instrctrs_6_cycs(x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_instrctrs_6_cycs),
    .io_in_instrctrs_6_iters(x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_instrctrs_6_iters),
    .io_in_instrctrs_6_stalls(x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_instrctrs_6_stalls),
    .io_in_instrctrs_6_idles(x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_instrctrs_6_idles),
    .io_sigsIn_done(x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_sigsIn_done),
    .io_sigsIn_backpressure(x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_baseEn(x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_sigsIn_baseEn),
    .io_sigsIn_break(x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_0(x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_rr(x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_rr)
  );
  assign _T_332 = io_sigsIn_done == 1'h0; // @[package.scala 100:49:@6814.4]
  assign _T_399 = RetimeWrapper_io_out; // @[package.scala 96:25:@6908.4 package.scala 96:25:@6909.4]
  assign _T_403 = ~ io_in_x107_b_0_empty; // @[sm_x131_outr_UnitPipe.scala 75:44:@6914.4]
  assign _T_404 = ~ io_in_x107_b_0_accessActivesOut_1; // @[sm_x131_outr_UnitPipe.scala 75:62:@6915.4]
  assign _T_405 = _T_403 | _T_404; // @[sm_x131_outr_UnitPipe.scala 75:60:@6916.4]
  assign x130_inr_Foreach_sigsIn_forwardpressure = _T_405 | x130_inr_Foreach_sm_io_doneLatch; // @[sm_x131_outr_UnitPipe.scala 75:95:@6917.4]
  assign _T_415 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@6951.4 package.scala 96:25:@6952.4]
  assign _T_421 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@6959.4 package.scala 96:25:@6960.4]
  assign _T_424 = ~ _T_421; // @[SpatialBlocks.scala 110:93:@6962.4]
  assign x130_inr_Foreach_sigsIn_baseEn = _T_415 & _T_424; // @[SpatialBlocks.scala 110:90:@6963.4]
  assign _T_426 = x130_inr_Foreach_sm_io_datapathEn; // @[SpatialBlocks.scala 128:36:@6971.4]
  assign _T_427 = ~ x130_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 128:78:@6972.4]
  assign _T_432 = x130_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 130:61:@6981.4]
  assign io_in_x95_TVALID = x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_x95_TVALID; // @[sm_x130_inr_Foreach.scala 50:22:@7083.4]
  assign io_in_x95_TDATA = x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_x95_TDATA; // @[sm_x130_inr_Foreach.scala 50:22:@7081.4]
  assign io_in_x95_TSTRB = x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_x95_TSTRB; // @[sm_x130_inr_Foreach.scala 50:22:@7080.4]
  assign io_in_x95_TKEEP = x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_x95_TKEEP; // @[sm_x130_inr_Foreach.scala 50:22:@7079.4]
  assign io_in_x95_TLAST = x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_x95_TLAST; // @[sm_x130_inr_Foreach.scala 50:22:@7078.4]
  assign io_in_x95_TID = x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_x95_TID; // @[sm_x130_inr_Foreach.scala 50:22:@7077.4]
  assign io_in_x95_TDEST = x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_x95_TDEST; // @[sm_x130_inr_Foreach.scala 50:22:@7076.4]
  assign io_in_x95_TUSER = x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_x95_TUSER; // @[sm_x130_inr_Foreach.scala 50:22:@7075.4]
  assign io_in_x107_b_0_rPort_0_en_0 = x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_x107_b_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@7093.4]
  assign io_in_x107_b_0_accessActivesIn_1 = x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_x107_b_0_accessActivesIn_1; // @[MemInterfaceType.scala 69:92:@7096.4]
  assign io_in_instrctrs_5_cycs = cycles_io_count; // @[Ledger.scala 282:21:@6819.4]
  assign io_in_instrctrs_5_iters = iters_io_count; // @[Ledger.scala 283:22:@6820.4]
  assign io_in_instrctrs_6_cycs = x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_instrctrs_6_cycs; // @[Ledger.scala 291:78:@7100.4]
  assign io_in_instrctrs_6_iters = x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_instrctrs_6_iters; // @[Ledger.scala 291:78:@7099.4]
  assign io_in_instrctrs_6_stalls = x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_instrctrs_6_stalls; // @[Ledger.scala 291:78:@7098.4]
  assign io_in_instrctrs_6_idles = x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_instrctrs_6_idles; // @[Ledger.scala 291:78:@7097.4]
  assign io_sigsOut_smDoneIn_0 = x130_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 127:53:@6969.4]
  assign io_sigsOut_smCtrCopyDone_0 = x130_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 139:125:@6985.4]
  assign cycles_clock = clock; // @[:@6808.4]
  assign cycles_reset = reset; // @[:@6809.4]
  assign cycles_io_enable = io_sigsIn_baseEn; // @[sm_x131_outr_UnitPipe.scala 65:24:@6813.4]
  assign iters_clock = clock; // @[:@6811.4]
  assign iters_reset = reset; // @[:@6812.4]
  assign iters_io_enable = io_sigsIn_done & _T_335; // @[sm_x131_outr_UnitPipe.scala 66:23:@6818.4]
  assign x118_ctrchain_clock = clock; // @[:@6824.4]
  assign x118_ctrchain_reset = reset; // @[:@6825.4]
  assign x118_ctrchain_io_input_reset = x130_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 130:103:@6984.4]
  assign x118_ctrchain_io_input_enable = _T_432 & x130_inr_Foreach_sigsIn_forwardpressure; // @[SpatialBlocks.scala 104:75:@6939.4 SpatialBlocks.scala 130:45:@6983.4]
  assign x130_inr_Foreach_sm_clock = clock; // @[:@6876.4]
  assign x130_inr_Foreach_sm_reset = reset; // @[:@6877.4]
  assign x130_inr_Foreach_sm_io_enable = x130_inr_Foreach_sigsIn_baseEn & x130_inr_Foreach_sigsIn_forwardpressure; // @[SpatialBlocks.scala 112:18:@6966.4]
  assign x130_inr_Foreach_sm_io_ctrDone = io_rr ? _T_399 : 1'h0; // @[sm_x131_outr_UnitPipe.scala 73:38:@6911.4]
  assign x130_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 114:21:@6968.4]
  assign x130_inr_Foreach_sm_io_backpressure = io_in_x95_TREADY | x130_inr_Foreach_sm_io_doneLatch; // @[SpatialBlocks.scala 105:24:@6940.4]
  assign x130_inr_Foreach_sm_io_break = 1'h0; // @[sm_x131_outr_UnitPipe.scala 77:36:@6920.4]
  assign RetimeWrapper_clock = clock; // @[:@6904.4]
  assign RetimeWrapper_reset = reset; // @[:@6905.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@6907.4]
  assign RetimeWrapper_io_in = x118_ctrchain_io_output_done; // @[package.scala 94:16:@6906.4]
  assign RetimeWrapper_1_clock = clock; // @[:@6947.4]
  assign RetimeWrapper_1_reset = reset; // @[:@6948.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@6950.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@6949.4]
  assign RetimeWrapper_2_clock = clock; // @[:@6955.4]
  assign RetimeWrapper_2_reset = reset; // @[:@6956.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@6958.4]
  assign RetimeWrapper_2_io_in = x130_inr_Foreach_sm_io_done; // @[package.scala 94:16:@6957.4]
  assign x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_clock = clock; // @[:@6987.4]
  assign x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_reset = reset; // @[:@6988.4]
  assign x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_x95_TREADY = io_in_x95_TREADY; // @[sm_x130_inr_Foreach.scala 50:22:@7082.4]
  assign x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_x107_b_0_rPort_0_output_0 = io_in_x107_b_0_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@7091.4]
  assign x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_x107_b_0_empty = io_in_x107_b_0_empty; // @[MemInterfaceType.scala 153:14:@7086.4]
  assign x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_in_x107_b_0_accessActivesOut_1 = io_in_x107_b_0_accessActivesOut_1; // @[MemInterfaceType.scala 156:25:@7090.4]
  assign x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_sigsIn_done = x130_inr_Foreach_sm_io_done; // @[sm_x130_inr_Foreach.scala 118:22:@7119.4]
  assign x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_sigsIn_backpressure = io_in_x95_TREADY | x130_inr_Foreach_sm_io_doneLatch; // @[sm_x130_inr_Foreach.scala 118:22:@7115.4]
  assign x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_426 & _T_427; // @[sm_x130_inr_Foreach.scala 118:22:@7113.4]
  assign x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_sigsIn_baseEn = _T_415 & _T_424; // @[sm_x130_inr_Foreach.scala 118:22:@7112.4]
  assign x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_sigsIn_break = x130_inr_Foreach_sm_io_break; // @[sm_x130_inr_Foreach.scala 118:22:@7111.4]
  assign x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = x118_ctrchain_io_output_counts_0; // @[sm_x130_inr_Foreach.scala 118:22:@7106.4]
  assign x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x118_ctrchain_io_output_oobs_0; // @[sm_x130_inr_Foreach.scala 118:22:@7105.4]
  assign x130_inr_Foreach_kernelx130_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x130_inr_Foreach.scala 117:18:@7101.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_335 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_335 <= 1'h0;
    end else begin
      _T_335 <= _T_332;
    end
  end
endmodule
module x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1( // @[:@7128.2]
  input         clock, // @[:@7129.4]
  input         reset, // @[:@7130.4]
  output        io_in_x95_TVALID, // @[:@7131.4]
  input         io_in_x95_TREADY, // @[:@7131.4]
  output [63:0] io_in_x95_TDATA, // @[:@7131.4]
  output [7:0]  io_in_x95_TSTRB, // @[:@7131.4]
  output [7:0]  io_in_x95_TKEEP, // @[:@7131.4]
  output        io_in_x95_TLAST, // @[:@7131.4]
  output [7:0]  io_in_x95_TID, // @[:@7131.4]
  output [7:0]  io_in_x95_TDEST, // @[:@7131.4]
  output [31:0] io_in_x95_TUSER, // @[:@7131.4]
  input         io_in_x90_TVALID, // @[:@7131.4]
  output        io_in_x90_TREADY, // @[:@7131.4]
  input  [63:0] io_in_x90_TDATA, // @[:@7131.4]
  input  [7:0]  io_in_x90_TID, // @[:@7131.4]
  input  [7:0]  io_in_x90_TDEST, // @[:@7131.4]
  output [63:0] io_in_instrctrs_1_cycs, // @[:@7131.4]
  output [63:0] io_in_instrctrs_1_iters, // @[:@7131.4]
  output [63:0] io_in_instrctrs_2_cycs, // @[:@7131.4]
  output [63:0] io_in_instrctrs_2_iters, // @[:@7131.4]
  output [63:0] io_in_instrctrs_3_cycs, // @[:@7131.4]
  output [63:0] io_in_instrctrs_3_iters, // @[:@7131.4]
  output [63:0] io_in_instrctrs_3_stalls, // @[:@7131.4]
  output [63:0] io_in_instrctrs_3_idles, // @[:@7131.4]
  output [63:0] io_in_instrctrs_4_cycs, // @[:@7131.4]
  output [63:0] io_in_instrctrs_4_iters, // @[:@7131.4]
  output [63:0] io_in_instrctrs_4_stalls, // @[:@7131.4]
  output [63:0] io_in_instrctrs_4_idles, // @[:@7131.4]
  output [63:0] io_in_instrctrs_5_cycs, // @[:@7131.4]
  output [63:0] io_in_instrctrs_5_iters, // @[:@7131.4]
  output [63:0] io_in_instrctrs_6_cycs, // @[:@7131.4]
  output [63:0] io_in_instrctrs_6_iters, // @[:@7131.4]
  output [63:0] io_in_instrctrs_6_stalls, // @[:@7131.4]
  output [63:0] io_in_instrctrs_6_idles, // @[:@7131.4]
  input         io_sigsIn_done, // @[:@7131.4]
  input         io_sigsIn_baseEn, // @[:@7131.4]
  input         io_sigsIn_smEnableOuts_0, // @[:@7131.4]
  input         io_sigsIn_smEnableOuts_1, // @[:@7131.4]
  input         io_sigsIn_smEnableOuts_2, // @[:@7131.4]
  input         io_sigsIn_smChildAcks_0, // @[:@7131.4]
  input         io_sigsIn_smChildAcks_1, // @[:@7131.4]
  input         io_sigsIn_smChildAcks_2, // @[:@7131.4]
  output        io_sigsOut_smDoneIn_0, // @[:@7131.4]
  output        io_sigsOut_smDoneIn_1, // @[:@7131.4]
  output        io_sigsOut_smDoneIn_2, // @[:@7131.4]
  output        io_sigsOut_smCtrCopyDone_0, // @[:@7131.4]
  output        io_sigsOut_smCtrCopyDone_1, // @[:@7131.4]
  output        io_sigsOut_smCtrCopyDone_2, // @[:@7131.4]
  input         io_rr // @[:@7131.4]
);
  wire  cycles_clock; // @[sm_x132_outr_UnitPipe.scala 62:26:@7177.4]
  wire  cycles_reset; // @[sm_x132_outr_UnitPipe.scala 62:26:@7177.4]
  wire  cycles_io_enable; // @[sm_x132_outr_UnitPipe.scala 62:26:@7177.4]
  wire [63:0] cycles_io_count; // @[sm_x132_outr_UnitPipe.scala 62:26:@7177.4]
  wire  iters_clock; // @[sm_x132_outr_UnitPipe.scala 63:25:@7180.4]
  wire  iters_reset; // @[sm_x132_outr_UnitPipe.scala 63:25:@7180.4]
  wire  iters_io_enable; // @[sm_x132_outr_UnitPipe.scala 63:25:@7180.4]
  wire [63:0] iters_io_count; // @[sm_x132_outr_UnitPipe.scala 63:25:@7180.4]
  wire  x97_a_0_clock; // @[m_x97_a_0.scala 27:17:@7193.4]
  wire  x97_a_0_reset; // @[m_x97_a_0.scala 27:17:@7193.4]
  wire  x97_a_0_io_rPort_0_en_0; // @[m_x97_a_0.scala 27:17:@7193.4]
  wire [31:0] x97_a_0_io_rPort_0_output_0; // @[m_x97_a_0.scala 27:17:@7193.4]
  wire [31:0] x97_a_0_io_wPort_0_data_0; // @[m_x97_a_0.scala 27:17:@7193.4]
  wire  x97_a_0_io_wPort_0_en_0; // @[m_x97_a_0.scala 27:17:@7193.4]
  wire  x97_a_0_io_full; // @[m_x97_a_0.scala 27:17:@7193.4]
  wire  x97_a_0_io_empty; // @[m_x97_a_0.scala 27:17:@7193.4]
  wire  x97_a_0_io_accessActivesOut_0; // @[m_x97_a_0.scala 27:17:@7193.4]
  wire  x97_a_0_io_accessActivesOut_1; // @[m_x97_a_0.scala 27:17:@7193.4]
  wire  x97_a_0_io_accessActivesIn_0; // @[m_x97_a_0.scala 27:17:@7193.4]
  wire  x97_a_0_io_accessActivesIn_1; // @[m_x97_a_0.scala 27:17:@7193.4]
  wire  x106_outr_UnitPipe_sm_clock; // @[sm_x106_outr_UnitPipe.scala 33:18:@7254.4]
  wire  x106_outr_UnitPipe_sm_reset; // @[sm_x106_outr_UnitPipe.scala 33:18:@7254.4]
  wire  x106_outr_UnitPipe_sm_io_enable; // @[sm_x106_outr_UnitPipe.scala 33:18:@7254.4]
  wire  x106_outr_UnitPipe_sm_io_done; // @[sm_x106_outr_UnitPipe.scala 33:18:@7254.4]
  wire  x106_outr_UnitPipe_sm_io_parentAck; // @[sm_x106_outr_UnitPipe.scala 33:18:@7254.4]
  wire  x106_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x106_outr_UnitPipe.scala 33:18:@7254.4]
  wire  x106_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x106_outr_UnitPipe.scala 33:18:@7254.4]
  wire  x106_outr_UnitPipe_sm_io_childAck_0; // @[sm_x106_outr_UnitPipe.scala 33:18:@7254.4]
  wire  x106_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x106_outr_UnitPipe.scala 33:18:@7254.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@7306.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@7306.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@7306.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@7306.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@7306.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@7314.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@7314.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@7314.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@7314.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@7314.4]
  wire  x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_clock; // @[sm_x106_outr_UnitPipe.scala 82:24:@7342.4]
  wire  x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_reset; // @[sm_x106_outr_UnitPipe.scala 82:24:@7342.4]
  wire [31:0] x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_in_x97_a_0_wPort_0_data_0; // @[sm_x106_outr_UnitPipe.scala 82:24:@7342.4]
  wire  x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_in_x97_a_0_wPort_0_en_0; // @[sm_x106_outr_UnitPipe.scala 82:24:@7342.4]
  wire  x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_in_x97_a_0_full; // @[sm_x106_outr_UnitPipe.scala 82:24:@7342.4]
  wire  x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_in_x97_a_0_accessActivesOut_0; // @[sm_x106_outr_UnitPipe.scala 82:24:@7342.4]
  wire  x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_in_x97_a_0_accessActivesIn_0; // @[sm_x106_outr_UnitPipe.scala 82:24:@7342.4]
  wire  x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_in_x90_TVALID; // @[sm_x106_outr_UnitPipe.scala 82:24:@7342.4]
  wire  x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_in_x90_TREADY; // @[sm_x106_outr_UnitPipe.scala 82:24:@7342.4]
  wire [63:0] x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_in_x90_TDATA; // @[sm_x106_outr_UnitPipe.scala 82:24:@7342.4]
  wire [7:0] x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_in_x90_TID; // @[sm_x106_outr_UnitPipe.scala 82:24:@7342.4]
  wire [7:0] x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_in_x90_TDEST; // @[sm_x106_outr_UnitPipe.scala 82:24:@7342.4]
  wire [63:0] x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_in_instrctrs_2_cycs; // @[sm_x106_outr_UnitPipe.scala 82:24:@7342.4]
  wire [63:0] x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_in_instrctrs_2_iters; // @[sm_x106_outr_UnitPipe.scala 82:24:@7342.4]
  wire [63:0] x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_in_instrctrs_3_cycs; // @[sm_x106_outr_UnitPipe.scala 82:24:@7342.4]
  wire [63:0] x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_in_instrctrs_3_iters; // @[sm_x106_outr_UnitPipe.scala 82:24:@7342.4]
  wire [63:0] x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_in_instrctrs_3_stalls; // @[sm_x106_outr_UnitPipe.scala 82:24:@7342.4]
  wire [63:0] x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_in_instrctrs_3_idles; // @[sm_x106_outr_UnitPipe.scala 82:24:@7342.4]
  wire  x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_sigsIn_done; // @[sm_x106_outr_UnitPipe.scala 82:24:@7342.4]
  wire  x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_sigsIn_baseEn; // @[sm_x106_outr_UnitPipe.scala 82:24:@7342.4]
  wire  x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x106_outr_UnitPipe.scala 82:24:@7342.4]
  wire  x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x106_outr_UnitPipe.scala 82:24:@7342.4]
  wire  x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x106_outr_UnitPipe.scala 82:24:@7342.4]
  wire  x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x106_outr_UnitPipe.scala 82:24:@7342.4]
  wire  x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_rr; // @[sm_x106_outr_UnitPipe.scala 82:24:@7342.4]
  wire  x107_b_0_clock; // @[m_x107_b_0.scala 27:17:@7489.4]
  wire  x107_b_0_reset; // @[m_x107_b_0.scala 27:17:@7489.4]
  wire  x107_b_0_io_rPort_0_en_0; // @[m_x107_b_0.scala 27:17:@7489.4]
  wire [31:0] x107_b_0_io_rPort_0_output_0; // @[m_x107_b_0.scala 27:17:@7489.4]
  wire [31:0] x107_b_0_io_wPort_0_data_0; // @[m_x107_b_0.scala 27:17:@7489.4]
  wire  x107_b_0_io_wPort_0_en_0; // @[m_x107_b_0.scala 27:17:@7489.4]
  wire  x107_b_0_io_full; // @[m_x107_b_0.scala 27:17:@7489.4]
  wire  x107_b_0_io_empty; // @[m_x107_b_0.scala 27:17:@7489.4]
  wire  x107_b_0_io_accessActivesOut_0; // @[m_x107_b_0.scala 27:17:@7489.4]
  wire  x107_b_0_io_accessActivesOut_1; // @[m_x107_b_0.scala 27:17:@7489.4]
  wire  x107_b_0_io_accessActivesIn_0; // @[m_x107_b_0.scala 27:17:@7489.4]
  wire  x107_b_0_io_accessActivesIn_1; // @[m_x107_b_0.scala 27:17:@7489.4]
  wire  x109_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@7515.4]
  wire  x109_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@7515.4]
  wire  x109_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@7515.4]
  wire  x109_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@7515.4]
  wire [31:0] x109_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@7515.4]
  wire  x109_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@7515.4]
  wire  x109_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@7515.4]
  wire  x116_inr_Foreach_sm_clock; // @[sm_x116_inr_Foreach.scala 32:18:@7567.4]
  wire  x116_inr_Foreach_sm_reset; // @[sm_x116_inr_Foreach.scala 32:18:@7567.4]
  wire  x116_inr_Foreach_sm_io_enable; // @[sm_x116_inr_Foreach.scala 32:18:@7567.4]
  wire  x116_inr_Foreach_sm_io_done; // @[sm_x116_inr_Foreach.scala 32:18:@7567.4]
  wire  x116_inr_Foreach_sm_io_doneLatch; // @[sm_x116_inr_Foreach.scala 32:18:@7567.4]
  wire  x116_inr_Foreach_sm_io_ctrDone; // @[sm_x116_inr_Foreach.scala 32:18:@7567.4]
  wire  x116_inr_Foreach_sm_io_datapathEn; // @[sm_x116_inr_Foreach.scala 32:18:@7567.4]
  wire  x116_inr_Foreach_sm_io_ctrInc; // @[sm_x116_inr_Foreach.scala 32:18:@7567.4]
  wire  x116_inr_Foreach_sm_io_ctrRst; // @[sm_x116_inr_Foreach.scala 32:18:@7567.4]
  wire  x116_inr_Foreach_sm_io_parentAck; // @[sm_x116_inr_Foreach.scala 32:18:@7567.4]
  wire  x116_inr_Foreach_sm_io_backpressure; // @[sm_x116_inr_Foreach.scala 32:18:@7567.4]
  wire  x116_inr_Foreach_sm_io_break; // @[sm_x116_inr_Foreach.scala 32:18:@7567.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@7595.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@7595.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@7595.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@7595.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@7595.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@7641.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@7641.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@7641.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@7641.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@7641.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@7649.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@7649.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@7649.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@7649.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@7649.4]
  wire  x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_clock; // @[sm_x116_inr_Foreach.scala 96:24:@7681.4]
  wire  x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_reset; // @[sm_x116_inr_Foreach.scala 96:24:@7681.4]
  wire  x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_in_x97_a_0_rPort_0_en_0; // @[sm_x116_inr_Foreach.scala 96:24:@7681.4]
  wire [31:0] x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_in_x97_a_0_rPort_0_output_0; // @[sm_x116_inr_Foreach.scala 96:24:@7681.4]
  wire  x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_in_x97_a_0_empty; // @[sm_x116_inr_Foreach.scala 96:24:@7681.4]
  wire  x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_in_x97_a_0_accessActivesOut_1; // @[sm_x116_inr_Foreach.scala 96:24:@7681.4]
  wire  x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_in_x97_a_0_accessActivesIn_1; // @[sm_x116_inr_Foreach.scala 96:24:@7681.4]
  wire [31:0] x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_in_x107_b_0_wPort_0_data_0; // @[sm_x116_inr_Foreach.scala 96:24:@7681.4]
  wire  x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_in_x107_b_0_wPort_0_en_0; // @[sm_x116_inr_Foreach.scala 96:24:@7681.4]
  wire  x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_in_x107_b_0_full; // @[sm_x116_inr_Foreach.scala 96:24:@7681.4]
  wire  x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_in_x107_b_0_accessActivesOut_0; // @[sm_x116_inr_Foreach.scala 96:24:@7681.4]
  wire  x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_in_x107_b_0_accessActivesIn_0; // @[sm_x116_inr_Foreach.scala 96:24:@7681.4]
  wire [63:0] x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_in_instrctrs_4_cycs; // @[sm_x116_inr_Foreach.scala 96:24:@7681.4]
  wire [63:0] x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_in_instrctrs_4_iters; // @[sm_x116_inr_Foreach.scala 96:24:@7681.4]
  wire [63:0] x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_in_instrctrs_4_stalls; // @[sm_x116_inr_Foreach.scala 96:24:@7681.4]
  wire [63:0] x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_in_instrctrs_4_idles; // @[sm_x116_inr_Foreach.scala 96:24:@7681.4]
  wire  x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_sigsIn_done; // @[sm_x116_inr_Foreach.scala 96:24:@7681.4]
  wire  x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_sigsIn_backpressure; // @[sm_x116_inr_Foreach.scala 96:24:@7681.4]
  wire  x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x116_inr_Foreach.scala 96:24:@7681.4]
  wire  x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_sigsIn_baseEn; // @[sm_x116_inr_Foreach.scala 96:24:@7681.4]
  wire  x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x116_inr_Foreach.scala 96:24:@7681.4]
  wire [31:0] x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x116_inr_Foreach.scala 96:24:@7681.4]
  wire  x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x116_inr_Foreach.scala 96:24:@7681.4]
  wire  x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_rr; // @[sm_x116_inr_Foreach.scala 96:24:@7681.4]
  wire  x131_outr_UnitPipe_sm_clock; // @[sm_x131_outr_UnitPipe.scala 33:18:@7876.4]
  wire  x131_outr_UnitPipe_sm_reset; // @[sm_x131_outr_UnitPipe.scala 33:18:@7876.4]
  wire  x131_outr_UnitPipe_sm_io_enable; // @[sm_x131_outr_UnitPipe.scala 33:18:@7876.4]
  wire  x131_outr_UnitPipe_sm_io_done; // @[sm_x131_outr_UnitPipe.scala 33:18:@7876.4]
  wire  x131_outr_UnitPipe_sm_io_parentAck; // @[sm_x131_outr_UnitPipe.scala 33:18:@7876.4]
  wire  x131_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x131_outr_UnitPipe.scala 33:18:@7876.4]
  wire  x131_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x131_outr_UnitPipe.scala 33:18:@7876.4]
  wire  x131_outr_UnitPipe_sm_io_childAck_0; // @[sm_x131_outr_UnitPipe.scala 33:18:@7876.4]
  wire  x131_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x131_outr_UnitPipe.scala 33:18:@7876.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@7928.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@7928.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@7928.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@7928.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@7928.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@7936.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@7936.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@7936.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@7936.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@7936.4]
  wire  x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_clock; // @[sm_x131_outr_UnitPipe.scala 82:24:@7964.4]
  wire  x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_reset; // @[sm_x131_outr_UnitPipe.scala 82:24:@7964.4]
  wire  x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_x95_TVALID; // @[sm_x131_outr_UnitPipe.scala 82:24:@7964.4]
  wire  x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_x95_TREADY; // @[sm_x131_outr_UnitPipe.scala 82:24:@7964.4]
  wire [63:0] x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_x95_TDATA; // @[sm_x131_outr_UnitPipe.scala 82:24:@7964.4]
  wire [7:0] x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_x95_TSTRB; // @[sm_x131_outr_UnitPipe.scala 82:24:@7964.4]
  wire [7:0] x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_x95_TKEEP; // @[sm_x131_outr_UnitPipe.scala 82:24:@7964.4]
  wire  x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_x95_TLAST; // @[sm_x131_outr_UnitPipe.scala 82:24:@7964.4]
  wire [7:0] x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_x95_TID; // @[sm_x131_outr_UnitPipe.scala 82:24:@7964.4]
  wire [7:0] x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_x95_TDEST; // @[sm_x131_outr_UnitPipe.scala 82:24:@7964.4]
  wire [31:0] x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_x95_TUSER; // @[sm_x131_outr_UnitPipe.scala 82:24:@7964.4]
  wire  x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_x107_b_0_rPort_0_en_0; // @[sm_x131_outr_UnitPipe.scala 82:24:@7964.4]
  wire [31:0] x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_x107_b_0_rPort_0_output_0; // @[sm_x131_outr_UnitPipe.scala 82:24:@7964.4]
  wire  x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_x107_b_0_empty; // @[sm_x131_outr_UnitPipe.scala 82:24:@7964.4]
  wire  x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_x107_b_0_accessActivesOut_1; // @[sm_x131_outr_UnitPipe.scala 82:24:@7964.4]
  wire  x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_x107_b_0_accessActivesIn_1; // @[sm_x131_outr_UnitPipe.scala 82:24:@7964.4]
  wire [63:0] x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_instrctrs_5_cycs; // @[sm_x131_outr_UnitPipe.scala 82:24:@7964.4]
  wire [63:0] x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_instrctrs_5_iters; // @[sm_x131_outr_UnitPipe.scala 82:24:@7964.4]
  wire [63:0] x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_instrctrs_6_cycs; // @[sm_x131_outr_UnitPipe.scala 82:24:@7964.4]
  wire [63:0] x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_instrctrs_6_iters; // @[sm_x131_outr_UnitPipe.scala 82:24:@7964.4]
  wire [63:0] x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_instrctrs_6_stalls; // @[sm_x131_outr_UnitPipe.scala 82:24:@7964.4]
  wire [63:0] x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_instrctrs_6_idles; // @[sm_x131_outr_UnitPipe.scala 82:24:@7964.4]
  wire  x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_sigsIn_done; // @[sm_x131_outr_UnitPipe.scala 82:24:@7964.4]
  wire  x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_sigsIn_baseEn; // @[sm_x131_outr_UnitPipe.scala 82:24:@7964.4]
  wire  x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x131_outr_UnitPipe.scala 82:24:@7964.4]
  wire  x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x131_outr_UnitPipe.scala 82:24:@7964.4]
  wire  x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x131_outr_UnitPipe.scala 82:24:@7964.4]
  wire  x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x131_outr_UnitPipe.scala 82:24:@7964.4]
  wire  x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_rr; // @[sm_x131_outr_UnitPipe.scala 82:24:@7964.4]
  wire  _T_204; // @[package.scala 100:49:@7184.4]
  reg  _T_207; // @[package.scala 48:56:@7185.4]
  reg [31:0] _RAND_0;
  wire  _T_281; // @[package.scala 96:25:@7311.4 package.scala 96:25:@7312.4]
  wire  _T_287; // @[package.scala 96:25:@7319.4 package.scala 96:25:@7320.4]
  wire  _T_290; // @[SpatialBlocks.scala 110:93:@7322.4]
  wire  _T_359; // @[package.scala 96:25:@7600.4 package.scala 96:25:@7601.4]
  wire  _T_362; // @[sm_x132_outr_UnitPipe.scala 83:41:@7604.4]
  wire  _T_363; // @[sm_x132_outr_UnitPipe.scala 83:58:@7605.4]
  wire  _T_364; // @[sm_x132_outr_UnitPipe.scala 83:56:@7606.4]
  wire  _T_366; // @[sm_x132_outr_UnitPipe.scala 84:44:@7609.4]
  wire  _T_367; // @[sm_x132_outr_UnitPipe.scala 84:61:@7610.4]
  wire  _T_368; // @[sm_x132_outr_UnitPipe.scala 84:59:@7611.4]
  wire  x116_inr_Foreach_sigsIn_forwardpressure; // @[sm_x132_outr_UnitPipe.scala 84:93:@7612.4]
  wire  _T_378; // @[package.scala 96:25:@7646.4 package.scala 96:25:@7647.4]
  wire  _T_384; // @[package.scala 96:25:@7654.4 package.scala 96:25:@7655.4]
  wire  _T_387; // @[SpatialBlocks.scala 110:93:@7657.4]
  wire  x116_inr_Foreach_sigsIn_baseEn; // @[SpatialBlocks.scala 110:90:@7658.4]
  wire  _T_389; // @[SpatialBlocks.scala 128:36:@7666.4]
  wire  _T_390; // @[SpatialBlocks.scala 128:78:@7667.4]
  wire  _T_395; // @[SpatialBlocks.scala 130:61:@7676.4]
  wire  _T_466; // @[package.scala 96:25:@7933.4 package.scala 96:25:@7934.4]
  wire  _T_472; // @[package.scala 96:25:@7941.4 package.scala 96:25:@7942.4]
  wire  _T_475; // @[SpatialBlocks.scala 110:93:@7944.4]
  InstrumentationCounter cycles ( // @[sm_x132_outr_UnitPipe.scala 62:26:@7177.4]
    .clock(cycles_clock),
    .reset(cycles_reset),
    .io_enable(cycles_io_enable),
    .io_count(cycles_io_count)
  );
  InstrumentationCounter iters ( // @[sm_x132_outr_UnitPipe.scala 63:25:@7180.4]
    .clock(iters_clock),
    .reset(iters_reset),
    .io_enable(iters_io_enable),
    .io_count(iters_io_count)
  );
  x97_a_0 x97_a_0 ( // @[m_x97_a_0.scala 27:17:@7193.4]
    .clock(x97_a_0_clock),
    .reset(x97_a_0_reset),
    .io_rPort_0_en_0(x97_a_0_io_rPort_0_en_0),
    .io_rPort_0_output_0(x97_a_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(x97_a_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x97_a_0_io_wPort_0_en_0),
    .io_full(x97_a_0_io_full),
    .io_empty(x97_a_0_io_empty),
    .io_accessActivesOut_0(x97_a_0_io_accessActivesOut_0),
    .io_accessActivesOut_1(x97_a_0_io_accessActivesOut_1),
    .io_accessActivesIn_0(x97_a_0_io_accessActivesIn_0),
    .io_accessActivesIn_1(x97_a_0_io_accessActivesIn_1)
  );
  x106_outr_UnitPipe_sm x106_outr_UnitPipe_sm ( // @[sm_x106_outr_UnitPipe.scala 33:18:@7254.4]
    .clock(x106_outr_UnitPipe_sm_clock),
    .reset(x106_outr_UnitPipe_sm_reset),
    .io_enable(x106_outr_UnitPipe_sm_io_enable),
    .io_done(x106_outr_UnitPipe_sm_io_done),
    .io_parentAck(x106_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x106_outr_UnitPipe_sm_io_doneIn_0),
    .io_enableOut_0(x106_outr_UnitPipe_sm_io_enableOut_0),
    .io_childAck_0(x106_outr_UnitPipe_sm_io_childAck_0),
    .io_ctrCopyDone_0(x106_outr_UnitPipe_sm_io_ctrCopyDone_0)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@7306.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@7314.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1 x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1 ( // @[sm_x106_outr_UnitPipe.scala 82:24:@7342.4]
    .clock(x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_clock),
    .reset(x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_reset),
    .io_in_x97_a_0_wPort_0_data_0(x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_in_x97_a_0_wPort_0_data_0),
    .io_in_x97_a_0_wPort_0_en_0(x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_in_x97_a_0_wPort_0_en_0),
    .io_in_x97_a_0_full(x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_in_x97_a_0_full),
    .io_in_x97_a_0_accessActivesOut_0(x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_in_x97_a_0_accessActivesOut_0),
    .io_in_x97_a_0_accessActivesIn_0(x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_in_x97_a_0_accessActivesIn_0),
    .io_in_x90_TVALID(x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_in_x90_TVALID),
    .io_in_x90_TREADY(x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_in_x90_TREADY),
    .io_in_x90_TDATA(x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_in_x90_TDATA),
    .io_in_x90_TID(x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_in_x90_TID),
    .io_in_x90_TDEST(x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_in_x90_TDEST),
    .io_in_instrctrs_2_cycs(x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_in_instrctrs_2_cycs),
    .io_in_instrctrs_2_iters(x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_in_instrctrs_2_iters),
    .io_in_instrctrs_3_cycs(x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_in_instrctrs_3_cycs),
    .io_in_instrctrs_3_iters(x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_in_instrctrs_3_iters),
    .io_in_instrctrs_3_stalls(x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_in_instrctrs_3_stalls),
    .io_in_instrctrs_3_idles(x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_in_instrctrs_3_idles),
    .io_sigsIn_done(x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_sigsIn_done),
    .io_sigsIn_baseEn(x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_sigsIn_baseEn),
    .io_sigsIn_smEnableOuts_0(x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smCtrCopyDone_0(x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_rr(x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_rr)
  );
  x97_a_0 x107_b_0 ( // @[m_x107_b_0.scala 27:17:@7489.4]
    .clock(x107_b_0_clock),
    .reset(x107_b_0_reset),
    .io_rPort_0_en_0(x107_b_0_io_rPort_0_en_0),
    .io_rPort_0_output_0(x107_b_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(x107_b_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x107_b_0_io_wPort_0_en_0),
    .io_full(x107_b_0_io_full),
    .io_empty(x107_b_0_io_empty),
    .io_accessActivesOut_0(x107_b_0_io_accessActivesOut_0),
    .io_accessActivesOut_1(x107_b_0_io_accessActivesOut_1),
    .io_accessActivesIn_0(x107_b_0_io_accessActivesIn_0),
    .io_accessActivesIn_1(x107_b_0_io_accessActivesIn_1)
  );
  x99_ctrchain x109_ctrchain ( // @[SpatialBlocks.scala 37:22:@7515.4]
    .clock(x109_ctrchain_clock),
    .reset(x109_ctrchain_reset),
    .io_input_reset(x109_ctrchain_io_input_reset),
    .io_input_enable(x109_ctrchain_io_input_enable),
    .io_output_counts_0(x109_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x109_ctrchain_io_output_oobs_0),
    .io_output_done(x109_ctrchain_io_output_done)
  );
  x116_inr_Foreach_sm x116_inr_Foreach_sm ( // @[sm_x116_inr_Foreach.scala 32:18:@7567.4]
    .clock(x116_inr_Foreach_sm_clock),
    .reset(x116_inr_Foreach_sm_reset),
    .io_enable(x116_inr_Foreach_sm_io_enable),
    .io_done(x116_inr_Foreach_sm_io_done),
    .io_doneLatch(x116_inr_Foreach_sm_io_doneLatch),
    .io_ctrDone(x116_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x116_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x116_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x116_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x116_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x116_inr_Foreach_sm_io_backpressure),
    .io_break(x116_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@7595.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@7641.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@7649.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  x116_inr_Foreach_kernelx116_inr_Foreach_concrete1 x116_inr_Foreach_kernelx116_inr_Foreach_concrete1 ( // @[sm_x116_inr_Foreach.scala 96:24:@7681.4]
    .clock(x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_clock),
    .reset(x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_reset),
    .io_in_x97_a_0_rPort_0_en_0(x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_in_x97_a_0_rPort_0_en_0),
    .io_in_x97_a_0_rPort_0_output_0(x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_in_x97_a_0_rPort_0_output_0),
    .io_in_x97_a_0_empty(x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_in_x97_a_0_empty),
    .io_in_x97_a_0_accessActivesOut_1(x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_in_x97_a_0_accessActivesOut_1),
    .io_in_x97_a_0_accessActivesIn_1(x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_in_x97_a_0_accessActivesIn_1),
    .io_in_x107_b_0_wPort_0_data_0(x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_in_x107_b_0_wPort_0_data_0),
    .io_in_x107_b_0_wPort_0_en_0(x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_in_x107_b_0_wPort_0_en_0),
    .io_in_x107_b_0_full(x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_in_x107_b_0_full),
    .io_in_x107_b_0_accessActivesOut_0(x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_in_x107_b_0_accessActivesOut_0),
    .io_in_x107_b_0_accessActivesIn_0(x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_in_x107_b_0_accessActivesIn_0),
    .io_in_instrctrs_4_cycs(x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_in_instrctrs_4_cycs),
    .io_in_instrctrs_4_iters(x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_in_instrctrs_4_iters),
    .io_in_instrctrs_4_stalls(x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_in_instrctrs_4_stalls),
    .io_in_instrctrs_4_idles(x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_in_instrctrs_4_idles),
    .io_sigsIn_done(x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_sigsIn_done),
    .io_sigsIn_backpressure(x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_baseEn(x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_sigsIn_baseEn),
    .io_sigsIn_break(x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_0(x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_rr(x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_rr)
  );
  x106_outr_UnitPipe_sm x131_outr_UnitPipe_sm ( // @[sm_x131_outr_UnitPipe.scala 33:18:@7876.4]
    .clock(x131_outr_UnitPipe_sm_clock),
    .reset(x131_outr_UnitPipe_sm_reset),
    .io_enable(x131_outr_UnitPipe_sm_io_enable),
    .io_done(x131_outr_UnitPipe_sm_io_done),
    .io_parentAck(x131_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x131_outr_UnitPipe_sm_io_doneIn_0),
    .io_enableOut_0(x131_outr_UnitPipe_sm_io_enableOut_0),
    .io_childAck_0(x131_outr_UnitPipe_sm_io_childAck_0),
    .io_ctrCopyDone_0(x131_outr_UnitPipe_sm_io_ctrCopyDone_0)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@7928.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@7936.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1 x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1 ( // @[sm_x131_outr_UnitPipe.scala 82:24:@7964.4]
    .clock(x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_clock),
    .reset(x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_reset),
    .io_in_x95_TVALID(x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_x95_TVALID),
    .io_in_x95_TREADY(x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_x95_TREADY),
    .io_in_x95_TDATA(x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_x95_TDATA),
    .io_in_x95_TSTRB(x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_x95_TSTRB),
    .io_in_x95_TKEEP(x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_x95_TKEEP),
    .io_in_x95_TLAST(x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_x95_TLAST),
    .io_in_x95_TID(x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_x95_TID),
    .io_in_x95_TDEST(x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_x95_TDEST),
    .io_in_x95_TUSER(x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_x95_TUSER),
    .io_in_x107_b_0_rPort_0_en_0(x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_x107_b_0_rPort_0_en_0),
    .io_in_x107_b_0_rPort_0_output_0(x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_x107_b_0_rPort_0_output_0),
    .io_in_x107_b_0_empty(x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_x107_b_0_empty),
    .io_in_x107_b_0_accessActivesOut_1(x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_x107_b_0_accessActivesOut_1),
    .io_in_x107_b_0_accessActivesIn_1(x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_x107_b_0_accessActivesIn_1),
    .io_in_instrctrs_5_cycs(x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_instrctrs_5_cycs),
    .io_in_instrctrs_5_iters(x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_instrctrs_5_iters),
    .io_in_instrctrs_6_cycs(x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_instrctrs_6_cycs),
    .io_in_instrctrs_6_iters(x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_instrctrs_6_iters),
    .io_in_instrctrs_6_stalls(x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_instrctrs_6_stalls),
    .io_in_instrctrs_6_idles(x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_instrctrs_6_idles),
    .io_sigsIn_done(x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_sigsIn_done),
    .io_sigsIn_baseEn(x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_sigsIn_baseEn),
    .io_sigsIn_smEnableOuts_0(x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smCtrCopyDone_0(x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_rr(x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_rr)
  );
  assign _T_204 = io_sigsIn_done == 1'h0; // @[package.scala 100:49:@7184.4]
  assign _T_281 = RetimeWrapper_io_out; // @[package.scala 96:25:@7311.4 package.scala 96:25:@7312.4]
  assign _T_287 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@7319.4 package.scala 96:25:@7320.4]
  assign _T_290 = ~ _T_287; // @[SpatialBlocks.scala 110:93:@7322.4]
  assign _T_359 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@7600.4 package.scala 96:25:@7601.4]
  assign _T_362 = ~ x107_b_0_io_full; // @[sm_x132_outr_UnitPipe.scala 83:41:@7604.4]
  assign _T_363 = ~ x107_b_0_io_accessActivesOut_0; // @[sm_x132_outr_UnitPipe.scala 83:58:@7605.4]
  assign _T_364 = _T_362 | _T_363; // @[sm_x132_outr_UnitPipe.scala 83:56:@7606.4]
  assign _T_366 = ~ x97_a_0_io_empty; // @[sm_x132_outr_UnitPipe.scala 84:44:@7609.4]
  assign _T_367 = ~ x97_a_0_io_accessActivesOut_1; // @[sm_x132_outr_UnitPipe.scala 84:61:@7610.4]
  assign _T_368 = _T_366 | _T_367; // @[sm_x132_outr_UnitPipe.scala 84:59:@7611.4]
  assign x116_inr_Foreach_sigsIn_forwardpressure = _T_368 | x116_inr_Foreach_sm_io_doneLatch; // @[sm_x132_outr_UnitPipe.scala 84:93:@7612.4]
  assign _T_378 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@7646.4 package.scala 96:25:@7647.4]
  assign _T_384 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@7654.4 package.scala 96:25:@7655.4]
  assign _T_387 = ~ _T_384; // @[SpatialBlocks.scala 110:93:@7657.4]
  assign x116_inr_Foreach_sigsIn_baseEn = _T_378 & _T_387; // @[SpatialBlocks.scala 110:90:@7658.4]
  assign _T_389 = x116_inr_Foreach_sm_io_datapathEn; // @[SpatialBlocks.scala 128:36:@7666.4]
  assign _T_390 = ~ x116_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 128:78:@7667.4]
  assign _T_395 = x116_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 130:61:@7676.4]
  assign _T_466 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@7933.4 package.scala 96:25:@7934.4]
  assign _T_472 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@7941.4 package.scala 96:25:@7942.4]
  assign _T_475 = ~ _T_472; // @[SpatialBlocks.scala 110:93:@7944.4]
  assign io_in_x95_TVALID = x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_x95_TVALID; // @[sm_x131_outr_UnitPipe.scala 50:22:@8061.4]
  assign io_in_x95_TDATA = x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_x95_TDATA; // @[sm_x131_outr_UnitPipe.scala 50:22:@8059.4]
  assign io_in_x95_TSTRB = x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_x95_TSTRB; // @[sm_x131_outr_UnitPipe.scala 50:22:@8058.4]
  assign io_in_x95_TKEEP = x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_x95_TKEEP; // @[sm_x131_outr_UnitPipe.scala 50:22:@8057.4]
  assign io_in_x95_TLAST = x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_x95_TLAST; // @[sm_x131_outr_UnitPipe.scala 50:22:@8056.4]
  assign io_in_x95_TID = x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_x95_TID; // @[sm_x131_outr_UnitPipe.scala 50:22:@8055.4]
  assign io_in_x95_TDEST = x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_x95_TDEST; // @[sm_x131_outr_UnitPipe.scala 50:22:@8054.4]
  assign io_in_x95_TUSER = x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_x95_TUSER; // @[sm_x131_outr_UnitPipe.scala 50:22:@8053.4]
  assign io_in_x90_TREADY = x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_in_x90_TREADY; // @[sm_x106_outr_UnitPipe.scala 51:22:@7453.4]
  assign io_in_instrctrs_1_cycs = cycles_io_count; // @[Ledger.scala 282:21:@7189.4]
  assign io_in_instrctrs_1_iters = iters_io_count; // @[Ledger.scala 283:22:@7190.4]
  assign io_in_instrctrs_2_cycs = x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_in_instrctrs_2_cycs; // @[Ledger.scala 291:78:@7458.4]
  assign io_in_instrctrs_2_iters = x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_in_instrctrs_2_iters; // @[Ledger.scala 291:78:@7457.4]
  assign io_in_instrctrs_3_cycs = x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_in_instrctrs_3_cycs; // @[Ledger.scala 291:78:@7462.4]
  assign io_in_instrctrs_3_iters = x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_in_instrctrs_3_iters; // @[Ledger.scala 291:78:@7461.4]
  assign io_in_instrctrs_3_stalls = x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_in_instrctrs_3_stalls; // @[Ledger.scala 291:78:@7460.4]
  assign io_in_instrctrs_3_idles = x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_in_instrctrs_3_idles; // @[Ledger.scala 291:78:@7459.4]
  assign io_in_instrctrs_4_cycs = x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_in_instrctrs_4_cycs; // @[Ledger.scala 291:78:@7814.4]
  assign io_in_instrctrs_4_iters = x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_in_instrctrs_4_iters; // @[Ledger.scala 291:78:@7813.4]
  assign io_in_instrctrs_4_stalls = x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_in_instrctrs_4_stalls; // @[Ledger.scala 291:78:@7812.4]
  assign io_in_instrctrs_4_idles = x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_in_instrctrs_4_idles; // @[Ledger.scala 291:78:@7811.4]
  assign io_in_instrctrs_5_cycs = x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_instrctrs_5_cycs; // @[Ledger.scala 291:78:@8078.4]
  assign io_in_instrctrs_5_iters = x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_instrctrs_5_iters; // @[Ledger.scala 291:78:@8077.4]
  assign io_in_instrctrs_6_cycs = x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_instrctrs_6_cycs; // @[Ledger.scala 291:78:@8082.4]
  assign io_in_instrctrs_6_iters = x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_instrctrs_6_iters; // @[Ledger.scala 291:78:@8081.4]
  assign io_in_instrctrs_6_stalls = x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_instrctrs_6_stalls; // @[Ledger.scala 291:78:@8080.4]
  assign io_in_instrctrs_6_idles = x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_instrctrs_6_idles; // @[Ledger.scala 291:78:@8079.4]
  assign io_sigsOut_smDoneIn_0 = x106_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 127:53:@7329.4]
  assign io_sigsOut_smDoneIn_1 = x116_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 127:53:@7664.4]
  assign io_sigsOut_smDoneIn_2 = x131_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 127:53:@7951.4]
  assign io_sigsOut_smCtrCopyDone_0 = x106_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 139:125:@7341.4]
  assign io_sigsOut_smCtrCopyDone_1 = x116_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 139:125:@7680.4]
  assign io_sigsOut_smCtrCopyDone_2 = x131_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 139:125:@7963.4]
  assign cycles_clock = clock; // @[:@7178.4]
  assign cycles_reset = reset; // @[:@7179.4]
  assign cycles_io_enable = io_sigsIn_baseEn; // @[sm_x132_outr_UnitPipe.scala 64:24:@7183.4]
  assign iters_clock = clock; // @[:@7181.4]
  assign iters_reset = reset; // @[:@7182.4]
  assign iters_io_enable = io_sigsIn_done & _T_207; // @[sm_x132_outr_UnitPipe.scala 65:23:@7188.4]
  assign x97_a_0_clock = clock; // @[:@7194.4]
  assign x97_a_0_reset = reset; // @[:@7195.4]
  assign x97_a_0_io_rPort_0_en_0 = x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_in_x97_a_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@7792.4]
  assign x97_a_0_io_wPort_0_data_0 = x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_in_x97_a_0_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@7442.4]
  assign x97_a_0_io_wPort_0_en_0 = x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_in_x97_a_0_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@7438.4]
  assign x97_a_0_io_accessActivesIn_0 = x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_in_x97_a_0_accessActivesIn_0; // @[MemInterfaceType.scala 69:92:@7445.4]
  assign x97_a_0_io_accessActivesIn_1 = x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_in_x97_a_0_accessActivesIn_1; // @[MemInterfaceType.scala 69:92:@7795.4]
  assign x106_outr_UnitPipe_sm_clock = clock; // @[:@7255.4]
  assign x106_outr_UnitPipe_sm_reset = reset; // @[:@7256.4]
  assign x106_outr_UnitPipe_sm_io_enable = _T_281 & _T_290; // @[SpatialBlocks.scala 112:18:@7326.4]
  assign x106_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 114:21:@7328.4]
  assign x106_outr_UnitPipe_sm_io_doneIn_0 = x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 102:67:@7298.4]
  assign x106_outr_UnitPipe_sm_io_ctrCopyDone_0 = x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 132:80:@7340.4]
  assign RetimeWrapper_clock = clock; // @[:@7307.4]
  assign RetimeWrapper_reset = reset; // @[:@7308.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@7310.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@7309.4]
  assign RetimeWrapper_1_clock = clock; // @[:@7315.4]
  assign RetimeWrapper_1_reset = reset; // @[:@7316.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@7318.4]
  assign RetimeWrapper_1_io_in = x106_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@7317.4]
  assign x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_clock = clock; // @[:@7343.4]
  assign x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_reset = reset; // @[:@7344.4]
  assign x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_in_x97_a_0_full = x97_a_0_io_full; // @[MemInterfaceType.scala 151:13:@7431.4]
  assign x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_in_x97_a_0_accessActivesOut_0 = x97_a_0_io_accessActivesOut_0; // @[MemInterfaceType.scala 156:25:@7436.4]
  assign x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_in_x90_TVALID = io_in_x90_TVALID; // @[sm_x106_outr_UnitPipe.scala 51:22:@7454.4]
  assign x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_in_x90_TDATA = io_in_x90_TDATA; // @[sm_x106_outr_UnitPipe.scala 51:22:@7452.4]
  assign x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_in_x90_TID = io_in_x90_TID; // @[sm_x106_outr_UnitPipe.scala 51:22:@7448.4]
  assign x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_in_x90_TDEST = io_in_x90_TDEST; // @[sm_x106_outr_UnitPipe.scala 51:22:@7447.4]
  assign x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_sigsIn_done = x106_outr_UnitPipe_sm_io_done; // @[sm_x106_outr_UnitPipe.scala 87:22:@7481.4]
  assign x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_sigsIn_baseEn = _T_281 & _T_290; // @[sm_x106_outr_UnitPipe.scala 87:22:@7474.4]
  assign x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x106_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x106_outr_UnitPipe.scala 87:22:@7471.4]
  assign x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x106_outr_UnitPipe_sm_io_childAck_0; // @[sm_x106_outr_UnitPipe.scala 87:22:@7469.4]
  assign x106_outr_UnitPipe_kernelx106_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x106_outr_UnitPipe.scala 86:18:@7463.4]
  assign x107_b_0_clock = clock; // @[:@7490.4]
  assign x107_b_0_reset = reset; // @[:@7491.4]
  assign x107_b_0_io_rPort_0_en_0 = x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_x107_b_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@8071.4]
  assign x107_b_0_io_wPort_0_data_0 = x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_in_x107_b_0_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@7807.4]
  assign x107_b_0_io_wPort_0_en_0 = x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_in_x107_b_0_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@7803.4]
  assign x107_b_0_io_accessActivesIn_0 = x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_in_x107_b_0_accessActivesIn_0; // @[MemInterfaceType.scala 69:92:@7810.4]
  assign x107_b_0_io_accessActivesIn_1 = x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_x107_b_0_accessActivesIn_1; // @[MemInterfaceType.scala 69:92:@8074.4]
  assign x109_ctrchain_clock = clock; // @[:@7516.4]
  assign x109_ctrchain_reset = reset; // @[:@7517.4]
  assign x109_ctrchain_io_input_reset = x116_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 130:103:@7679.4]
  assign x109_ctrchain_io_input_enable = _T_395 & x116_inr_Foreach_sigsIn_forwardpressure; // @[SpatialBlocks.scala 104:75:@7634.4 SpatialBlocks.scala 130:45:@7678.4]
  assign x116_inr_Foreach_sm_clock = clock; // @[:@7568.4]
  assign x116_inr_Foreach_sm_reset = reset; // @[:@7569.4]
  assign x116_inr_Foreach_sm_io_enable = x116_inr_Foreach_sigsIn_baseEn & x116_inr_Foreach_sigsIn_forwardpressure; // @[SpatialBlocks.scala 112:18:@7661.4]
  assign x116_inr_Foreach_sm_io_ctrDone = io_rr ? _T_359 : 1'h0; // @[sm_x132_outr_UnitPipe.scala 82:38:@7603.4]
  assign x116_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 114:21:@7663.4]
  assign x116_inr_Foreach_sm_io_backpressure = _T_364 | x116_inr_Foreach_sm_io_doneLatch; // @[SpatialBlocks.scala 105:24:@7635.4]
  assign x116_inr_Foreach_sm_io_break = 1'h0; // @[sm_x132_outr_UnitPipe.scala 86:36:@7615.4]
  assign RetimeWrapper_2_clock = clock; // @[:@7596.4]
  assign RetimeWrapper_2_reset = reset; // @[:@7597.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@7599.4]
  assign RetimeWrapper_2_io_in = x109_ctrchain_io_output_done; // @[package.scala 94:16:@7598.4]
  assign RetimeWrapper_3_clock = clock; // @[:@7642.4]
  assign RetimeWrapper_3_reset = reset; // @[:@7643.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@7645.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@7644.4]
  assign RetimeWrapper_4_clock = clock; // @[:@7650.4]
  assign RetimeWrapper_4_reset = reset; // @[:@7651.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@7653.4]
  assign RetimeWrapper_4_io_in = x116_inr_Foreach_sm_io_done; // @[package.scala 94:16:@7652.4]
  assign x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_clock = clock; // @[:@7682.4]
  assign x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_reset = reset; // @[:@7683.4]
  assign x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_in_x97_a_0_rPort_0_output_0 = x97_a_0_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@7790.4]
  assign x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_in_x97_a_0_empty = x97_a_0_io_empty; // @[MemInterfaceType.scala 153:14:@7785.4]
  assign x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_in_x97_a_0_accessActivesOut_1 = x97_a_0_io_accessActivesOut_1; // @[MemInterfaceType.scala 156:25:@7789.4]
  assign x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_in_x107_b_0_full = x107_b_0_io_full; // @[MemInterfaceType.scala 151:13:@7796.4]
  assign x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_in_x107_b_0_accessActivesOut_0 = x107_b_0_io_accessActivesOut_0; // @[MemInterfaceType.scala 156:25:@7801.4]
  assign x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_sigsIn_done = x116_inr_Foreach_sm_io_done; // @[sm_x116_inr_Foreach.scala 101:22:@7833.4]
  assign x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_sigsIn_backpressure = _T_364 | x116_inr_Foreach_sm_io_doneLatch; // @[sm_x116_inr_Foreach.scala 101:22:@7829.4]
  assign x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_389 & _T_390; // @[sm_x116_inr_Foreach.scala 101:22:@7827.4]
  assign x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_sigsIn_baseEn = _T_378 & _T_387; // @[sm_x116_inr_Foreach.scala 101:22:@7826.4]
  assign x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_sigsIn_break = x116_inr_Foreach_sm_io_break; // @[sm_x116_inr_Foreach.scala 101:22:@7825.4]
  assign x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = x109_ctrchain_io_output_counts_0; // @[sm_x116_inr_Foreach.scala 101:22:@7820.4]
  assign x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x109_ctrchain_io_output_oobs_0; // @[sm_x116_inr_Foreach.scala 101:22:@7819.4]
  assign x116_inr_Foreach_kernelx116_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x116_inr_Foreach.scala 100:18:@7815.4]
  assign x131_outr_UnitPipe_sm_clock = clock; // @[:@7877.4]
  assign x131_outr_UnitPipe_sm_reset = reset; // @[:@7878.4]
  assign x131_outr_UnitPipe_sm_io_enable = _T_466 & _T_475; // @[SpatialBlocks.scala 112:18:@7948.4]
  assign x131_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_2; // @[SpatialBlocks.scala 114:21:@7950.4]
  assign x131_outr_UnitPipe_sm_io_doneIn_0 = x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 102:67:@7920.4]
  assign x131_outr_UnitPipe_sm_io_ctrCopyDone_0 = x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 132:80:@7962.4]
  assign RetimeWrapper_5_clock = clock; // @[:@7929.4]
  assign RetimeWrapper_5_reset = reset; // @[:@7930.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@7932.4]
  assign RetimeWrapper_5_io_in = io_sigsIn_smEnableOuts_2; // @[package.scala 94:16:@7931.4]
  assign RetimeWrapper_6_clock = clock; // @[:@7937.4]
  assign RetimeWrapper_6_reset = reset; // @[:@7938.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@7940.4]
  assign RetimeWrapper_6_io_in = x131_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@7939.4]
  assign x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_clock = clock; // @[:@7965.4]
  assign x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_reset = reset; // @[:@7966.4]
  assign x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_x95_TREADY = io_in_x95_TREADY; // @[sm_x131_outr_UnitPipe.scala 50:22:@8060.4]
  assign x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_x107_b_0_rPort_0_output_0 = x107_b_0_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@8069.4]
  assign x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_x107_b_0_empty = x107_b_0_io_empty; // @[MemInterfaceType.scala 153:14:@8064.4]
  assign x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_in_x107_b_0_accessActivesOut_1 = x107_b_0_io_accessActivesOut_1; // @[MemInterfaceType.scala 156:25:@8068.4]
  assign x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_sigsIn_done = x131_outr_UnitPipe_sm_io_done; // @[sm_x131_outr_UnitPipe.scala 87:22:@8101.4]
  assign x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_sigsIn_baseEn = _T_466 & _T_475; // @[sm_x131_outr_UnitPipe.scala 87:22:@8094.4]
  assign x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x131_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x131_outr_UnitPipe.scala 87:22:@8091.4]
  assign x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x131_outr_UnitPipe_sm_io_childAck_0; // @[sm_x131_outr_UnitPipe.scala 87:22:@8089.4]
  assign x131_outr_UnitPipe_kernelx131_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x131_outr_UnitPipe.scala 86:18:@8083.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_207 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_207 <= 1'h0;
    end else begin
      _T_207 <= _T_204;
    end
  end
endmodule
module RootController_kernelRootController_concrete1( // @[:@8110.2]
  input         clock, // @[:@8111.4]
  input         reset, // @[:@8112.4]
  output        io_in_x95_TVALID, // @[:@8113.4]
  input         io_in_x95_TREADY, // @[:@8113.4]
  output [63:0] io_in_x95_TDATA, // @[:@8113.4]
  output [7:0]  io_in_x95_TSTRB, // @[:@8113.4]
  output [7:0]  io_in_x95_TKEEP, // @[:@8113.4]
  output        io_in_x95_TLAST, // @[:@8113.4]
  output [7:0]  io_in_x95_TID, // @[:@8113.4]
  output [7:0]  io_in_x95_TDEST, // @[:@8113.4]
  output [31:0] io_in_x95_TUSER, // @[:@8113.4]
  input         io_in_x90_TVALID, // @[:@8113.4]
  output        io_in_x90_TREADY, // @[:@8113.4]
  input  [63:0] io_in_x90_TDATA, // @[:@8113.4]
  input  [7:0]  io_in_x90_TID, // @[:@8113.4]
  input  [7:0]  io_in_x90_TDEST, // @[:@8113.4]
  output [63:0] io_in_instrctrs_0_cycs, // @[:@8113.4]
  output [63:0] io_in_instrctrs_0_iters, // @[:@8113.4]
  output [63:0] io_in_instrctrs_1_cycs, // @[:@8113.4]
  output [63:0] io_in_instrctrs_1_iters, // @[:@8113.4]
  output [63:0] io_in_instrctrs_2_cycs, // @[:@8113.4]
  output [63:0] io_in_instrctrs_2_iters, // @[:@8113.4]
  output [63:0] io_in_instrctrs_3_cycs, // @[:@8113.4]
  output [63:0] io_in_instrctrs_3_iters, // @[:@8113.4]
  output [63:0] io_in_instrctrs_3_stalls, // @[:@8113.4]
  output [63:0] io_in_instrctrs_3_idles, // @[:@8113.4]
  output [63:0] io_in_instrctrs_4_cycs, // @[:@8113.4]
  output [63:0] io_in_instrctrs_4_iters, // @[:@8113.4]
  output [63:0] io_in_instrctrs_4_stalls, // @[:@8113.4]
  output [63:0] io_in_instrctrs_4_idles, // @[:@8113.4]
  output [63:0] io_in_instrctrs_5_cycs, // @[:@8113.4]
  output [63:0] io_in_instrctrs_5_iters, // @[:@8113.4]
  output [63:0] io_in_instrctrs_6_cycs, // @[:@8113.4]
  output [63:0] io_in_instrctrs_6_iters, // @[:@8113.4]
  output [63:0] io_in_instrctrs_6_stalls, // @[:@8113.4]
  output [63:0] io_in_instrctrs_6_idles, // @[:@8113.4]
  input         io_sigsIn_done, // @[:@8113.4]
  input         io_sigsIn_baseEn, // @[:@8113.4]
  input         io_sigsIn_smEnableOuts_0, // @[:@8113.4]
  input         io_sigsIn_smChildAcks_0, // @[:@8113.4]
  output        io_sigsOut_smDoneIn_0, // @[:@8113.4]
  input         io_rr // @[:@8113.4]
);
  wire  cycles_clock; // @[sm_RootController.scala 62:26:@8151.4]
  wire  cycles_reset; // @[sm_RootController.scala 62:26:@8151.4]
  wire  cycles_io_enable; // @[sm_RootController.scala 62:26:@8151.4]
  wire [63:0] cycles_io_count; // @[sm_RootController.scala 62:26:@8151.4]
  wire  iters_clock; // @[sm_RootController.scala 63:25:@8154.4]
  wire  iters_reset; // @[sm_RootController.scala 63:25:@8154.4]
  wire  iters_io_enable; // @[sm_RootController.scala 63:25:@8154.4]
  wire [63:0] iters_io_count; // @[sm_RootController.scala 63:25:@8154.4]
  wire  x132_outr_UnitPipe_sm_clock; // @[sm_x132_outr_UnitPipe.scala 32:18:@8226.4]
  wire  x132_outr_UnitPipe_sm_reset; // @[sm_x132_outr_UnitPipe.scala 32:18:@8226.4]
  wire  x132_outr_UnitPipe_sm_io_enable; // @[sm_x132_outr_UnitPipe.scala 32:18:@8226.4]
  wire  x132_outr_UnitPipe_sm_io_done; // @[sm_x132_outr_UnitPipe.scala 32:18:@8226.4]
  wire  x132_outr_UnitPipe_sm_io_parentAck; // @[sm_x132_outr_UnitPipe.scala 32:18:@8226.4]
  wire  x132_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x132_outr_UnitPipe.scala 32:18:@8226.4]
  wire  x132_outr_UnitPipe_sm_io_doneIn_1; // @[sm_x132_outr_UnitPipe.scala 32:18:@8226.4]
  wire  x132_outr_UnitPipe_sm_io_doneIn_2; // @[sm_x132_outr_UnitPipe.scala 32:18:@8226.4]
  wire  x132_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x132_outr_UnitPipe.scala 32:18:@8226.4]
  wire  x132_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x132_outr_UnitPipe.scala 32:18:@8226.4]
  wire  x132_outr_UnitPipe_sm_io_enableOut_2; // @[sm_x132_outr_UnitPipe.scala 32:18:@8226.4]
  wire  x132_outr_UnitPipe_sm_io_childAck_0; // @[sm_x132_outr_UnitPipe.scala 32:18:@8226.4]
  wire  x132_outr_UnitPipe_sm_io_childAck_1; // @[sm_x132_outr_UnitPipe.scala 32:18:@8226.4]
  wire  x132_outr_UnitPipe_sm_io_childAck_2; // @[sm_x132_outr_UnitPipe.scala 32:18:@8226.4]
  wire  x132_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x132_outr_UnitPipe.scala 32:18:@8226.4]
  wire  x132_outr_UnitPipe_sm_io_ctrCopyDone_1; // @[sm_x132_outr_UnitPipe.scala 32:18:@8226.4]
  wire  x132_outr_UnitPipe_sm_io_ctrCopyDone_2; // @[sm_x132_outr_UnitPipe.scala 32:18:@8226.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@8298.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@8298.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@8298.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@8298.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@8298.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@8306.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@8306.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@8306.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@8306.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@8306.4]
  wire  x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_clock; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire  x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_reset; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire  x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_x95_TVALID; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire  x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_x95_TREADY; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire [63:0] x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_x95_TDATA; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire [7:0] x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_x95_TSTRB; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire [7:0] x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_x95_TKEEP; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire  x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_x95_TLAST; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire [7:0] x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_x95_TID; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire [7:0] x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_x95_TDEST; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire [31:0] x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_x95_TUSER; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire  x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_x90_TVALID; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire  x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_x90_TREADY; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire [63:0] x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_x90_TDATA; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire [7:0] x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_x90_TID; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire [7:0] x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_x90_TDEST; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire [63:0] x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_1_cycs; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire [63:0] x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_1_iters; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire [63:0] x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_2_cycs; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire [63:0] x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_2_iters; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire [63:0] x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_3_cycs; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire [63:0] x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_3_iters; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire [63:0] x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_3_stalls; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire [63:0] x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_3_idles; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire [63:0] x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_4_cycs; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire [63:0] x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_4_iters; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire [63:0] x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_4_stalls; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire [63:0] x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_4_idles; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire [63:0] x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_5_cycs; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire [63:0] x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_5_iters; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire [63:0] x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_6_cycs; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire [63:0] x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_6_iters; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire [63:0] x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_6_stalls; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire [63:0] x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_6_idles; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire  x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_sigsIn_done; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire  x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_sigsIn_baseEn; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire  x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire  x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire  x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire  x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire  x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire  x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire  x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire  x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire  x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire  x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire  x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire  x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire  x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_rr; // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
  wire  _T_180; // @[package.scala 100:49:@8158.4]
  reg  _T_183; // @[package.scala 48:56:@8159.4]
  reg [31:0] _RAND_0;
  wire  _T_268; // @[package.scala 96:25:@8303.4 package.scala 96:25:@8304.4]
  wire  _T_274; // @[package.scala 96:25:@8311.4 package.scala 96:25:@8312.4]
  wire  _T_277; // @[SpatialBlocks.scala 110:93:@8314.4]
  InstrumentationCounter cycles ( // @[sm_RootController.scala 62:26:@8151.4]
    .clock(cycles_clock),
    .reset(cycles_reset),
    .io_enable(cycles_io_enable),
    .io_count(cycles_io_count)
  );
  InstrumentationCounter iters ( // @[sm_RootController.scala 63:25:@8154.4]
    .clock(iters_clock),
    .reset(iters_reset),
    .io_enable(iters_io_enable),
    .io_count(iters_io_count)
  );
  x132_outr_UnitPipe_sm x132_outr_UnitPipe_sm ( // @[sm_x132_outr_UnitPipe.scala 32:18:@8226.4]
    .clock(x132_outr_UnitPipe_sm_clock),
    .reset(x132_outr_UnitPipe_sm_reset),
    .io_enable(x132_outr_UnitPipe_sm_io_enable),
    .io_done(x132_outr_UnitPipe_sm_io_done),
    .io_parentAck(x132_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x132_outr_UnitPipe_sm_io_doneIn_0),
    .io_doneIn_1(x132_outr_UnitPipe_sm_io_doneIn_1),
    .io_doneIn_2(x132_outr_UnitPipe_sm_io_doneIn_2),
    .io_enableOut_0(x132_outr_UnitPipe_sm_io_enableOut_0),
    .io_enableOut_1(x132_outr_UnitPipe_sm_io_enableOut_1),
    .io_enableOut_2(x132_outr_UnitPipe_sm_io_enableOut_2),
    .io_childAck_0(x132_outr_UnitPipe_sm_io_childAck_0),
    .io_childAck_1(x132_outr_UnitPipe_sm_io_childAck_1),
    .io_childAck_2(x132_outr_UnitPipe_sm_io_childAck_2),
    .io_ctrCopyDone_0(x132_outr_UnitPipe_sm_io_ctrCopyDone_0),
    .io_ctrCopyDone_1(x132_outr_UnitPipe_sm_io_ctrCopyDone_1),
    .io_ctrCopyDone_2(x132_outr_UnitPipe_sm_io_ctrCopyDone_2)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@8298.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@8306.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1 x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1 ( // @[sm_x132_outr_UnitPipe.scala 99:24:@8335.4]
    .clock(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_clock),
    .reset(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_reset),
    .io_in_x95_TVALID(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_x95_TVALID),
    .io_in_x95_TREADY(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_x95_TREADY),
    .io_in_x95_TDATA(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_x95_TDATA),
    .io_in_x95_TSTRB(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_x95_TSTRB),
    .io_in_x95_TKEEP(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_x95_TKEEP),
    .io_in_x95_TLAST(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_x95_TLAST),
    .io_in_x95_TID(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_x95_TID),
    .io_in_x95_TDEST(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_x95_TDEST),
    .io_in_x95_TUSER(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_x95_TUSER),
    .io_in_x90_TVALID(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_x90_TVALID),
    .io_in_x90_TREADY(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_x90_TREADY),
    .io_in_x90_TDATA(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_x90_TDATA),
    .io_in_x90_TID(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_x90_TID),
    .io_in_x90_TDEST(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_x90_TDEST),
    .io_in_instrctrs_1_cycs(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_1_cycs),
    .io_in_instrctrs_1_iters(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_1_iters),
    .io_in_instrctrs_2_cycs(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_2_cycs),
    .io_in_instrctrs_2_iters(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_2_iters),
    .io_in_instrctrs_3_cycs(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_3_cycs),
    .io_in_instrctrs_3_iters(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_3_iters),
    .io_in_instrctrs_3_stalls(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_3_stalls),
    .io_in_instrctrs_3_idles(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_3_idles),
    .io_in_instrctrs_4_cycs(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_4_cycs),
    .io_in_instrctrs_4_iters(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_4_iters),
    .io_in_instrctrs_4_stalls(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_4_stalls),
    .io_in_instrctrs_4_idles(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_4_idles),
    .io_in_instrctrs_5_cycs(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_5_cycs),
    .io_in_instrctrs_5_iters(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_5_iters),
    .io_in_instrctrs_6_cycs(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_6_cycs),
    .io_in_instrctrs_6_iters(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_6_iters),
    .io_in_instrctrs_6_stalls(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_6_stalls),
    .io_in_instrctrs_6_idles(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_6_idles),
    .io_sigsIn_done(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_sigsIn_done),
    .io_sigsIn_baseEn(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_sigsIn_baseEn),
    .io_sigsIn_smEnableOuts_0(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smEnableOuts_2(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2),
    .io_sigsIn_smChildAcks_0(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsIn_smChildAcks_2(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2),
    .io_sigsOut_smDoneIn_0(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1),
    .io_sigsOut_smDoneIn_2(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2),
    .io_sigsOut_smCtrCopyDone_0(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_sigsOut_smCtrCopyDone_1(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1),
    .io_sigsOut_smCtrCopyDone_2(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2),
    .io_rr(x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_rr)
  );
  assign _T_180 = io_sigsIn_done == 1'h0; // @[package.scala 100:49:@8158.4]
  assign _T_268 = RetimeWrapper_io_out; // @[package.scala 96:25:@8303.4 package.scala 96:25:@8304.4]
  assign _T_274 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@8311.4 package.scala 96:25:@8312.4]
  assign _T_277 = ~ _T_274; // @[SpatialBlocks.scala 110:93:@8314.4]
  assign io_in_x95_TVALID = x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_x95_TVALID; // @[sm_x132_outr_UnitPipe.scala 49:22:@8443.4]
  assign io_in_x95_TDATA = x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_x95_TDATA; // @[sm_x132_outr_UnitPipe.scala 49:22:@8441.4]
  assign io_in_x95_TSTRB = x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_x95_TSTRB; // @[sm_x132_outr_UnitPipe.scala 49:22:@8440.4]
  assign io_in_x95_TKEEP = x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_x95_TKEEP; // @[sm_x132_outr_UnitPipe.scala 49:22:@8439.4]
  assign io_in_x95_TLAST = x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_x95_TLAST; // @[sm_x132_outr_UnitPipe.scala 49:22:@8438.4]
  assign io_in_x95_TID = x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_x95_TID; // @[sm_x132_outr_UnitPipe.scala 49:22:@8437.4]
  assign io_in_x95_TDEST = x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_x95_TDEST; // @[sm_x132_outr_UnitPipe.scala 49:22:@8436.4]
  assign io_in_x95_TUSER = x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_x95_TUSER; // @[sm_x132_outr_UnitPipe.scala 49:22:@8435.4]
  assign io_in_x90_TREADY = x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_x90_TREADY; // @[sm_x132_outr_UnitPipe.scala 50:22:@8451.4]
  assign io_in_instrctrs_0_cycs = cycles_io_count; // @[Ledger.scala 282:21:@8163.4]
  assign io_in_instrctrs_0_iters = iters_io_count; // @[Ledger.scala 283:22:@8164.4]
  assign io_in_instrctrs_1_cycs = x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_1_cycs; // @[Ledger.scala 291:78:@8456.4]
  assign io_in_instrctrs_1_iters = x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_1_iters; // @[Ledger.scala 291:78:@8455.4]
  assign io_in_instrctrs_2_cycs = x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_2_cycs; // @[Ledger.scala 291:78:@8460.4]
  assign io_in_instrctrs_2_iters = x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_2_iters; // @[Ledger.scala 291:78:@8459.4]
  assign io_in_instrctrs_3_cycs = x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_3_cycs; // @[Ledger.scala 291:78:@8464.4]
  assign io_in_instrctrs_3_iters = x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_3_iters; // @[Ledger.scala 291:78:@8463.4]
  assign io_in_instrctrs_3_stalls = x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_3_stalls; // @[Ledger.scala 291:78:@8462.4]
  assign io_in_instrctrs_3_idles = x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_3_idles; // @[Ledger.scala 291:78:@8461.4]
  assign io_in_instrctrs_4_cycs = x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_4_cycs; // @[Ledger.scala 291:78:@8468.4]
  assign io_in_instrctrs_4_iters = x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_4_iters; // @[Ledger.scala 291:78:@8467.4]
  assign io_in_instrctrs_4_stalls = x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_4_stalls; // @[Ledger.scala 291:78:@8466.4]
  assign io_in_instrctrs_4_idles = x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_4_idles; // @[Ledger.scala 291:78:@8465.4]
  assign io_in_instrctrs_5_cycs = x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_5_cycs; // @[Ledger.scala 291:78:@8472.4]
  assign io_in_instrctrs_5_iters = x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_5_iters; // @[Ledger.scala 291:78:@8471.4]
  assign io_in_instrctrs_6_cycs = x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_6_cycs; // @[Ledger.scala 291:78:@8476.4]
  assign io_in_instrctrs_6_iters = x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_6_iters; // @[Ledger.scala 291:78:@8475.4]
  assign io_in_instrctrs_6_stalls = x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_6_stalls; // @[Ledger.scala 291:78:@8474.4]
  assign io_in_instrctrs_6_idles = x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_instrctrs_6_idles; // @[Ledger.scala 291:78:@8473.4]
  assign io_sigsOut_smDoneIn_0 = x132_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 127:53:@8321.4]
  assign cycles_clock = clock; // @[:@8152.4]
  assign cycles_reset = reset; // @[:@8153.4]
  assign cycles_io_enable = io_sigsIn_baseEn; // @[sm_RootController.scala 64:24:@8157.4]
  assign iters_clock = clock; // @[:@8155.4]
  assign iters_reset = reset; // @[:@8156.4]
  assign iters_io_enable = io_sigsIn_done & _T_183; // @[sm_RootController.scala 65:23:@8162.4]
  assign x132_outr_UnitPipe_sm_clock = clock; // @[:@8227.4]
  assign x132_outr_UnitPipe_sm_reset = reset; // @[:@8228.4]
  assign x132_outr_UnitPipe_sm_io_enable = _T_268 & _T_277; // @[SpatialBlocks.scala 112:18:@8318.4]
  assign x132_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 114:21:@8320.4]
  assign x132_outr_UnitPipe_sm_io_doneIn_0 = x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 102:67:@8286.4]
  assign x132_outr_UnitPipe_sm_io_doneIn_1 = x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 102:67:@8287.4]
  assign x132_outr_UnitPipe_sm_io_doneIn_2 = x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2; // @[SpatialBlocks.scala 102:67:@8288.4]
  assign x132_outr_UnitPipe_sm_io_ctrCopyDone_0 = x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 132:80:@8332.4]
  assign x132_outr_UnitPipe_sm_io_ctrCopyDone_1 = x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[SpatialBlocks.scala 132:80:@8333.4]
  assign x132_outr_UnitPipe_sm_io_ctrCopyDone_2 = x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2; // @[SpatialBlocks.scala 132:80:@8334.4]
  assign RetimeWrapper_clock = clock; // @[:@8299.4]
  assign RetimeWrapper_reset = reset; // @[:@8300.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@8302.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@8301.4]
  assign RetimeWrapper_1_clock = clock; // @[:@8307.4]
  assign RetimeWrapper_1_reset = reset; // @[:@8308.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@8310.4]
  assign RetimeWrapper_1_io_in = x132_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@8309.4]
  assign x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_clock = clock; // @[:@8336.4]
  assign x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_reset = reset; // @[:@8337.4]
  assign x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_x95_TREADY = io_in_x95_TREADY; // @[sm_x132_outr_UnitPipe.scala 49:22:@8442.4]
  assign x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_x90_TVALID = io_in_x90_TVALID; // @[sm_x132_outr_UnitPipe.scala 50:22:@8452.4]
  assign x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_x90_TDATA = io_in_x90_TDATA; // @[sm_x132_outr_UnitPipe.scala 50:22:@8450.4]
  assign x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_x90_TID = io_in_x90_TID; // @[sm_x132_outr_UnitPipe.scala 50:22:@8446.4]
  assign x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_in_x90_TDEST = io_in_x90_TDEST; // @[sm_x132_outr_UnitPipe.scala 50:22:@8445.4]
  assign x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_sigsIn_done = x132_outr_UnitPipe_sm_io_done; // @[sm_x132_outr_UnitPipe.scala 104:22:@8511.4]
  assign x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_sigsIn_baseEn = _T_268 & _T_277; // @[sm_x132_outr_UnitPipe.scala 104:22:@8504.4]
  assign x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x132_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x132_outr_UnitPipe.scala 104:22:@8499.4]
  assign x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1 = x132_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x132_outr_UnitPipe.scala 104:22:@8500.4]
  assign x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2 = x132_outr_UnitPipe_sm_io_enableOut_2; // @[sm_x132_outr_UnitPipe.scala 104:22:@8501.4]
  assign x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x132_outr_UnitPipe_sm_io_childAck_0; // @[sm_x132_outr_UnitPipe.scala 104:22:@8493.4]
  assign x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1 = x132_outr_UnitPipe_sm_io_childAck_1; // @[sm_x132_outr_UnitPipe.scala 104:22:@8494.4]
  assign x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2 = x132_outr_UnitPipe_sm_io_childAck_2; // @[sm_x132_outr_UnitPipe.scala 104:22:@8495.4]
  assign x132_outr_UnitPipe_kernelx132_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x132_outr_UnitPipe.scala 103:18:@8477.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_183 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_183 <= 1'h0;
    end else begin
      _T_183 <= _T_180;
    end
  end
endmodule
module AccelUnit( // @[:@8528.2]
  input         clock, // @[:@8529.4]
  input         reset, // @[:@8530.4]
  input         io_enable, // @[:@8531.4]
  output        io_done, // @[:@8531.4]
  input         io_reset, // @[:@8531.4]
  input         io_memStreams_loads_0_cmd_ready, // @[:@8531.4]
  output        io_memStreams_loads_0_cmd_valid, // @[:@8531.4]
  output [63:0] io_memStreams_loads_0_cmd_bits_addr, // @[:@8531.4]
  output [31:0] io_memStreams_loads_0_cmd_bits_size, // @[:@8531.4]
  output        io_memStreams_loads_0_data_ready, // @[:@8531.4]
  input         io_memStreams_loads_0_data_valid, // @[:@8531.4]
  input  [31:0] io_memStreams_loads_0_data_bits_rdata_0, // @[:@8531.4]
  input  [31:0] io_memStreams_loads_0_data_bits_rdata_1, // @[:@8531.4]
  input  [31:0] io_memStreams_loads_0_data_bits_rdata_2, // @[:@8531.4]
  input  [31:0] io_memStreams_loads_0_data_bits_rdata_3, // @[:@8531.4]
  input  [31:0] io_memStreams_loads_0_data_bits_rdata_4, // @[:@8531.4]
  input  [31:0] io_memStreams_loads_0_data_bits_rdata_5, // @[:@8531.4]
  input  [31:0] io_memStreams_loads_0_data_bits_rdata_6, // @[:@8531.4]
  input  [31:0] io_memStreams_loads_0_data_bits_rdata_7, // @[:@8531.4]
  input  [31:0] io_memStreams_loads_0_data_bits_rdata_8, // @[:@8531.4]
  input  [31:0] io_memStreams_loads_0_data_bits_rdata_9, // @[:@8531.4]
  input  [31:0] io_memStreams_loads_0_data_bits_rdata_10, // @[:@8531.4]
  input  [31:0] io_memStreams_loads_0_data_bits_rdata_11, // @[:@8531.4]
  input  [31:0] io_memStreams_loads_0_data_bits_rdata_12, // @[:@8531.4]
  input  [31:0] io_memStreams_loads_0_data_bits_rdata_13, // @[:@8531.4]
  input  [31:0] io_memStreams_loads_0_data_bits_rdata_14, // @[:@8531.4]
  input  [31:0] io_memStreams_loads_0_data_bits_rdata_15, // @[:@8531.4]
  input         io_memStreams_stores_0_cmd_ready, // @[:@8531.4]
  output        io_memStreams_stores_0_cmd_valid, // @[:@8531.4]
  output [63:0] io_memStreams_stores_0_cmd_bits_addr, // @[:@8531.4]
  output [31:0] io_memStreams_stores_0_cmd_bits_size, // @[:@8531.4]
  input         io_memStreams_stores_0_data_ready, // @[:@8531.4]
  output        io_memStreams_stores_0_data_valid, // @[:@8531.4]
  output [31:0] io_memStreams_stores_0_data_bits_wdata_0, // @[:@8531.4]
  output [31:0] io_memStreams_stores_0_data_bits_wdata_1, // @[:@8531.4]
  output [31:0] io_memStreams_stores_0_data_bits_wdata_2, // @[:@8531.4]
  output [31:0] io_memStreams_stores_0_data_bits_wdata_3, // @[:@8531.4]
  output [31:0] io_memStreams_stores_0_data_bits_wdata_4, // @[:@8531.4]
  output [31:0] io_memStreams_stores_0_data_bits_wdata_5, // @[:@8531.4]
  output [31:0] io_memStreams_stores_0_data_bits_wdata_6, // @[:@8531.4]
  output [31:0] io_memStreams_stores_0_data_bits_wdata_7, // @[:@8531.4]
  output [31:0] io_memStreams_stores_0_data_bits_wdata_8, // @[:@8531.4]
  output [31:0] io_memStreams_stores_0_data_bits_wdata_9, // @[:@8531.4]
  output [31:0] io_memStreams_stores_0_data_bits_wdata_10, // @[:@8531.4]
  output [31:0] io_memStreams_stores_0_data_bits_wdata_11, // @[:@8531.4]
  output [31:0] io_memStreams_stores_0_data_bits_wdata_12, // @[:@8531.4]
  output [31:0] io_memStreams_stores_0_data_bits_wdata_13, // @[:@8531.4]
  output [31:0] io_memStreams_stores_0_data_bits_wdata_14, // @[:@8531.4]
  output [31:0] io_memStreams_stores_0_data_bits_wdata_15, // @[:@8531.4]
  output [15:0] io_memStreams_stores_0_data_bits_wstrb, // @[:@8531.4]
  output        io_memStreams_stores_0_wresp_ready, // @[:@8531.4]
  input         io_memStreams_stores_0_wresp_valid, // @[:@8531.4]
  input         io_memStreams_stores_0_wresp_bits, // @[:@8531.4]
  input         io_memStreams_gathers_0_cmd_ready, // @[:@8531.4]
  output        io_memStreams_gathers_0_cmd_valid, // @[:@8531.4]
  output [63:0] io_memStreams_gathers_0_cmd_bits_addr_0, // @[:@8531.4]
  output [63:0] io_memStreams_gathers_0_cmd_bits_addr_1, // @[:@8531.4]
  output [63:0] io_memStreams_gathers_0_cmd_bits_addr_2, // @[:@8531.4]
  output [63:0] io_memStreams_gathers_0_cmd_bits_addr_3, // @[:@8531.4]
  output [63:0] io_memStreams_gathers_0_cmd_bits_addr_4, // @[:@8531.4]
  output [63:0] io_memStreams_gathers_0_cmd_bits_addr_5, // @[:@8531.4]
  output [63:0] io_memStreams_gathers_0_cmd_bits_addr_6, // @[:@8531.4]
  output [63:0] io_memStreams_gathers_0_cmd_bits_addr_7, // @[:@8531.4]
  output [63:0] io_memStreams_gathers_0_cmd_bits_addr_8, // @[:@8531.4]
  output [63:0] io_memStreams_gathers_0_cmd_bits_addr_9, // @[:@8531.4]
  output [63:0] io_memStreams_gathers_0_cmd_bits_addr_10, // @[:@8531.4]
  output [63:0] io_memStreams_gathers_0_cmd_bits_addr_11, // @[:@8531.4]
  output [63:0] io_memStreams_gathers_0_cmd_bits_addr_12, // @[:@8531.4]
  output [63:0] io_memStreams_gathers_0_cmd_bits_addr_13, // @[:@8531.4]
  output [63:0] io_memStreams_gathers_0_cmd_bits_addr_14, // @[:@8531.4]
  output [63:0] io_memStreams_gathers_0_cmd_bits_addr_15, // @[:@8531.4]
  output        io_memStreams_gathers_0_data_ready, // @[:@8531.4]
  input         io_memStreams_gathers_0_data_valid, // @[:@8531.4]
  input  [31:0] io_memStreams_gathers_0_data_bits_0, // @[:@8531.4]
  input  [31:0] io_memStreams_gathers_0_data_bits_1, // @[:@8531.4]
  input  [31:0] io_memStreams_gathers_0_data_bits_2, // @[:@8531.4]
  input  [31:0] io_memStreams_gathers_0_data_bits_3, // @[:@8531.4]
  input  [31:0] io_memStreams_gathers_0_data_bits_4, // @[:@8531.4]
  input  [31:0] io_memStreams_gathers_0_data_bits_5, // @[:@8531.4]
  input  [31:0] io_memStreams_gathers_0_data_bits_6, // @[:@8531.4]
  input  [31:0] io_memStreams_gathers_0_data_bits_7, // @[:@8531.4]
  input  [31:0] io_memStreams_gathers_0_data_bits_8, // @[:@8531.4]
  input  [31:0] io_memStreams_gathers_0_data_bits_9, // @[:@8531.4]
  input  [31:0] io_memStreams_gathers_0_data_bits_10, // @[:@8531.4]
  input  [31:0] io_memStreams_gathers_0_data_bits_11, // @[:@8531.4]
  input  [31:0] io_memStreams_gathers_0_data_bits_12, // @[:@8531.4]
  input  [31:0] io_memStreams_gathers_0_data_bits_13, // @[:@8531.4]
  input  [31:0] io_memStreams_gathers_0_data_bits_14, // @[:@8531.4]
  input  [31:0] io_memStreams_gathers_0_data_bits_15, // @[:@8531.4]
  input         io_memStreams_scatters_0_cmd_ready, // @[:@8531.4]
  output        io_memStreams_scatters_0_cmd_valid, // @[:@8531.4]
  output [63:0] io_memStreams_scatters_0_cmd_bits_addr_addr_0, // @[:@8531.4]
  output [63:0] io_memStreams_scatters_0_cmd_bits_addr_addr_1, // @[:@8531.4]
  output [63:0] io_memStreams_scatters_0_cmd_bits_addr_addr_2, // @[:@8531.4]
  output [63:0] io_memStreams_scatters_0_cmd_bits_addr_addr_3, // @[:@8531.4]
  output [63:0] io_memStreams_scatters_0_cmd_bits_addr_addr_4, // @[:@8531.4]
  output [63:0] io_memStreams_scatters_0_cmd_bits_addr_addr_5, // @[:@8531.4]
  output [63:0] io_memStreams_scatters_0_cmd_bits_addr_addr_6, // @[:@8531.4]
  output [63:0] io_memStreams_scatters_0_cmd_bits_addr_addr_7, // @[:@8531.4]
  output [63:0] io_memStreams_scatters_0_cmd_bits_addr_addr_8, // @[:@8531.4]
  output [63:0] io_memStreams_scatters_0_cmd_bits_addr_addr_9, // @[:@8531.4]
  output [63:0] io_memStreams_scatters_0_cmd_bits_addr_addr_10, // @[:@8531.4]
  output [63:0] io_memStreams_scatters_0_cmd_bits_addr_addr_11, // @[:@8531.4]
  output [63:0] io_memStreams_scatters_0_cmd_bits_addr_addr_12, // @[:@8531.4]
  output [63:0] io_memStreams_scatters_0_cmd_bits_addr_addr_13, // @[:@8531.4]
  output [63:0] io_memStreams_scatters_0_cmd_bits_addr_addr_14, // @[:@8531.4]
  output [63:0] io_memStreams_scatters_0_cmd_bits_addr_addr_15, // @[:@8531.4]
  output [31:0] io_memStreams_scatters_0_cmd_bits_wdata_0, // @[:@8531.4]
  output [31:0] io_memStreams_scatters_0_cmd_bits_wdata_1, // @[:@8531.4]
  output [31:0] io_memStreams_scatters_0_cmd_bits_wdata_2, // @[:@8531.4]
  output [31:0] io_memStreams_scatters_0_cmd_bits_wdata_3, // @[:@8531.4]
  output [31:0] io_memStreams_scatters_0_cmd_bits_wdata_4, // @[:@8531.4]
  output [31:0] io_memStreams_scatters_0_cmd_bits_wdata_5, // @[:@8531.4]
  output [31:0] io_memStreams_scatters_0_cmd_bits_wdata_6, // @[:@8531.4]
  output [31:0] io_memStreams_scatters_0_cmd_bits_wdata_7, // @[:@8531.4]
  output [31:0] io_memStreams_scatters_0_cmd_bits_wdata_8, // @[:@8531.4]
  output [31:0] io_memStreams_scatters_0_cmd_bits_wdata_9, // @[:@8531.4]
  output [31:0] io_memStreams_scatters_0_cmd_bits_wdata_10, // @[:@8531.4]
  output [31:0] io_memStreams_scatters_0_cmd_bits_wdata_11, // @[:@8531.4]
  output [31:0] io_memStreams_scatters_0_cmd_bits_wdata_12, // @[:@8531.4]
  output [31:0] io_memStreams_scatters_0_cmd_bits_wdata_13, // @[:@8531.4]
  output [31:0] io_memStreams_scatters_0_cmd_bits_wdata_14, // @[:@8531.4]
  output [31:0] io_memStreams_scatters_0_cmd_bits_wdata_15, // @[:@8531.4]
  output        io_memStreams_scatters_0_wresp_ready, // @[:@8531.4]
  input         io_memStreams_scatters_0_wresp_valid, // @[:@8531.4]
  input         io_memStreams_scatters_0_wresp_bits, // @[:@8531.4]
  input         io_axiStreamsIn_0_TVALID, // @[:@8531.4]
  output        io_axiStreamsIn_0_TREADY, // @[:@8531.4]
  input  [63:0] io_axiStreamsIn_0_TDATA, // @[:@8531.4]
  input  [7:0]  io_axiStreamsIn_0_TSTRB, // @[:@8531.4]
  input  [7:0]  io_axiStreamsIn_0_TKEEP, // @[:@8531.4]
  input         io_axiStreamsIn_0_TLAST, // @[:@8531.4]
  input  [7:0]  io_axiStreamsIn_0_TID, // @[:@8531.4]
  input  [7:0]  io_axiStreamsIn_0_TDEST, // @[:@8531.4]
  input  [31:0] io_axiStreamsIn_0_TUSER, // @[:@8531.4]
  output        io_axiStreamsOut_0_TVALID, // @[:@8531.4]
  input         io_axiStreamsOut_0_TREADY, // @[:@8531.4]
  output [63:0] io_axiStreamsOut_0_TDATA, // @[:@8531.4]
  output [7:0]  io_axiStreamsOut_0_TSTRB, // @[:@8531.4]
  output [7:0]  io_axiStreamsOut_0_TKEEP, // @[:@8531.4]
  output        io_axiStreamsOut_0_TLAST, // @[:@8531.4]
  output [7:0]  io_axiStreamsOut_0_TID, // @[:@8531.4]
  output [7:0]  io_axiStreamsOut_0_TDEST, // @[:@8531.4]
  output [31:0] io_axiStreamsOut_0_TUSER, // @[:@8531.4]
  output        io_heap_0_req_valid, // @[:@8531.4]
  output        io_heap_0_req_bits_allocDealloc, // @[:@8531.4]
  output [63:0] io_heap_0_req_bits_sizeAddr, // @[:@8531.4]
  input         io_heap_0_resp_valid, // @[:@8531.4]
  input         io_heap_0_resp_bits_allocDealloc, // @[:@8531.4]
  input  [63:0] io_heap_0_resp_bits_sizeAddr, // @[:@8531.4]
  input  [63:0] io_argIns_0, // @[:@8531.4]
  input         io_argOuts_0_port_ready, // @[:@8531.4]
  output        io_argOuts_0_port_valid, // @[:@8531.4]
  output [63:0] io_argOuts_0_port_bits, // @[:@8531.4]
  input  [63:0] io_argOuts_0_echo, // @[:@8531.4]
  input         io_argOuts_1_port_ready, // @[:@8531.4]
  output        io_argOuts_1_port_valid, // @[:@8531.4]
  output [63:0] io_argOuts_1_port_bits, // @[:@8531.4]
  input  [63:0] io_argOuts_1_echo, // @[:@8531.4]
  input         io_argOuts_2_port_ready, // @[:@8531.4]
  output        io_argOuts_2_port_valid, // @[:@8531.4]
  output [63:0] io_argOuts_2_port_bits, // @[:@8531.4]
  input  [63:0] io_argOuts_2_echo, // @[:@8531.4]
  input         io_argOuts_3_port_ready, // @[:@8531.4]
  output        io_argOuts_3_port_valid, // @[:@8531.4]
  output [63:0] io_argOuts_3_port_bits, // @[:@8531.4]
  input  [63:0] io_argOuts_3_echo, // @[:@8531.4]
  input         io_argOuts_4_port_ready, // @[:@8531.4]
  output        io_argOuts_4_port_valid, // @[:@8531.4]
  output [63:0] io_argOuts_4_port_bits, // @[:@8531.4]
  input  [63:0] io_argOuts_4_echo, // @[:@8531.4]
  input         io_argOuts_5_port_ready, // @[:@8531.4]
  output        io_argOuts_5_port_valid, // @[:@8531.4]
  output [63:0] io_argOuts_5_port_bits, // @[:@8531.4]
  input  [63:0] io_argOuts_5_echo, // @[:@8531.4]
  input         io_argOuts_6_port_ready, // @[:@8531.4]
  output        io_argOuts_6_port_valid, // @[:@8531.4]
  output [63:0] io_argOuts_6_port_bits, // @[:@8531.4]
  input  [63:0] io_argOuts_6_echo, // @[:@8531.4]
  input         io_argOuts_7_port_ready, // @[:@8531.4]
  output        io_argOuts_7_port_valid, // @[:@8531.4]
  output [63:0] io_argOuts_7_port_bits, // @[:@8531.4]
  input  [63:0] io_argOuts_7_echo, // @[:@8531.4]
  input         io_argOuts_8_port_ready, // @[:@8531.4]
  output        io_argOuts_8_port_valid, // @[:@8531.4]
  output [63:0] io_argOuts_8_port_bits, // @[:@8531.4]
  input  [63:0] io_argOuts_8_echo, // @[:@8531.4]
  input         io_argOuts_9_port_ready, // @[:@8531.4]
  output        io_argOuts_9_port_valid, // @[:@8531.4]
  output [63:0] io_argOuts_9_port_bits, // @[:@8531.4]
  input  [63:0] io_argOuts_9_echo, // @[:@8531.4]
  input         io_argOuts_10_port_ready, // @[:@8531.4]
  output        io_argOuts_10_port_valid, // @[:@8531.4]
  output [63:0] io_argOuts_10_port_bits, // @[:@8531.4]
  input  [63:0] io_argOuts_10_echo, // @[:@8531.4]
  input         io_argOuts_11_port_ready, // @[:@8531.4]
  output        io_argOuts_11_port_valid, // @[:@8531.4]
  output [63:0] io_argOuts_11_port_bits, // @[:@8531.4]
  input  [63:0] io_argOuts_11_echo, // @[:@8531.4]
  input         io_argOuts_12_port_ready, // @[:@8531.4]
  output        io_argOuts_12_port_valid, // @[:@8531.4]
  output [63:0] io_argOuts_12_port_bits, // @[:@8531.4]
  input  [63:0] io_argOuts_12_echo, // @[:@8531.4]
  input         io_argOuts_13_port_ready, // @[:@8531.4]
  output        io_argOuts_13_port_valid, // @[:@8531.4]
  output [63:0] io_argOuts_13_port_bits, // @[:@8531.4]
  input  [63:0] io_argOuts_13_echo, // @[:@8531.4]
  input         io_argOuts_14_port_ready, // @[:@8531.4]
  output        io_argOuts_14_port_valid, // @[:@8531.4]
  output [63:0] io_argOuts_14_port_bits, // @[:@8531.4]
  input  [63:0] io_argOuts_14_echo, // @[:@8531.4]
  input         io_argOuts_15_port_ready, // @[:@8531.4]
  output        io_argOuts_15_port_valid, // @[:@8531.4]
  output [63:0] io_argOuts_15_port_bits, // @[:@8531.4]
  input  [63:0] io_argOuts_15_echo, // @[:@8531.4]
  input         io_argOuts_16_port_ready, // @[:@8531.4]
  output        io_argOuts_16_port_valid, // @[:@8531.4]
  output [63:0] io_argOuts_16_port_bits, // @[:@8531.4]
  input  [63:0] io_argOuts_16_echo, // @[:@8531.4]
  input         io_argOuts_17_port_ready, // @[:@8531.4]
  output        io_argOuts_17_port_valid, // @[:@8531.4]
  output [63:0] io_argOuts_17_port_bits, // @[:@8531.4]
  input  [63:0] io_argOuts_17_echo, // @[:@8531.4]
  input         io_argOuts_18_port_ready, // @[:@8531.4]
  output        io_argOuts_18_port_valid, // @[:@8531.4]
  output [63:0] io_argOuts_18_port_bits, // @[:@8531.4]
  input  [63:0] io_argOuts_18_echo, // @[:@8531.4]
  input         io_argOuts_19_port_ready, // @[:@8531.4]
  output        io_argOuts_19_port_valid, // @[:@8531.4]
  output [63:0] io_argOuts_19_port_bits, // @[:@8531.4]
  input  [63:0] io_argOuts_19_echo // @[:@8531.4]
);
  wire  SingleCounter_clock; // @[Main.scala 29:32:@8765.4]
  wire  SingleCounter_reset; // @[Main.scala 29:32:@8765.4]
  wire  SingleCounter_io_input_reset; // @[Main.scala 29:32:@8765.4]
  wire  SingleCounter_io_output_done; // @[Main.scala 29:32:@8765.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@8783.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@8783.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@8783.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@8783.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@8783.4]
  wire  SRFF_clock; // @[Main.scala 34:28:@8799.4]
  wire  SRFF_reset; // @[Main.scala 34:28:@8799.4]
  wire  SRFF_io_input_set; // @[Main.scala 34:28:@8799.4]
  wire  SRFF_io_input_reset; // @[Main.scala 34:28:@8799.4]
  wire  SRFF_io_input_asyn_reset; // @[Main.scala 34:28:@8799.4]
  wire  SRFF_io_output; // @[Main.scala 34:28:@8799.4]
  wire  RootController_sm_clock; // @[sm_RootController.scala 32:18:@8837.4]
  wire  RootController_sm_reset; // @[sm_RootController.scala 32:18:@8837.4]
  wire  RootController_sm_io_enable; // @[sm_RootController.scala 32:18:@8837.4]
  wire  RootController_sm_io_done; // @[sm_RootController.scala 32:18:@8837.4]
  wire  RootController_sm_io_rst; // @[sm_RootController.scala 32:18:@8837.4]
  wire  RootController_sm_io_ctrDone; // @[sm_RootController.scala 32:18:@8837.4]
  wire  RootController_sm_io_ctrInc; // @[sm_RootController.scala 32:18:@8837.4]
  wire  RootController_sm_io_doneIn_0; // @[sm_RootController.scala 32:18:@8837.4]
  wire  RootController_sm_io_enableOut_0; // @[sm_RootController.scala 32:18:@8837.4]
  wire  RootController_sm_io_childAck_0; // @[sm_RootController.scala 32:18:@8837.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@8869.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@8869.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@8869.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@8869.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@8869.4]
  wire  RootController_kernelRootController_concrete1_clock; // @[sm_RootController.scala 76:24:@8928.4]
  wire  RootController_kernelRootController_concrete1_reset; // @[sm_RootController.scala 76:24:@8928.4]
  wire  RootController_kernelRootController_concrete1_io_in_x95_TVALID; // @[sm_RootController.scala 76:24:@8928.4]
  wire  RootController_kernelRootController_concrete1_io_in_x95_TREADY; // @[sm_RootController.scala 76:24:@8928.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x95_TDATA; // @[sm_RootController.scala 76:24:@8928.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x95_TSTRB; // @[sm_RootController.scala 76:24:@8928.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x95_TKEEP; // @[sm_RootController.scala 76:24:@8928.4]
  wire  RootController_kernelRootController_concrete1_io_in_x95_TLAST; // @[sm_RootController.scala 76:24:@8928.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x95_TID; // @[sm_RootController.scala 76:24:@8928.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x95_TDEST; // @[sm_RootController.scala 76:24:@8928.4]
  wire [31:0] RootController_kernelRootController_concrete1_io_in_x95_TUSER; // @[sm_RootController.scala 76:24:@8928.4]
  wire  RootController_kernelRootController_concrete1_io_in_x90_TVALID; // @[sm_RootController.scala 76:24:@8928.4]
  wire  RootController_kernelRootController_concrete1_io_in_x90_TREADY; // @[sm_RootController.scala 76:24:@8928.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x90_TDATA; // @[sm_RootController.scala 76:24:@8928.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x90_TID; // @[sm_RootController.scala 76:24:@8928.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x90_TDEST; // @[sm_RootController.scala 76:24:@8928.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_0_cycs; // @[sm_RootController.scala 76:24:@8928.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_0_iters; // @[sm_RootController.scala 76:24:@8928.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_1_cycs; // @[sm_RootController.scala 76:24:@8928.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_1_iters; // @[sm_RootController.scala 76:24:@8928.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_2_cycs; // @[sm_RootController.scala 76:24:@8928.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_2_iters; // @[sm_RootController.scala 76:24:@8928.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_3_cycs; // @[sm_RootController.scala 76:24:@8928.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_3_iters; // @[sm_RootController.scala 76:24:@8928.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_3_stalls; // @[sm_RootController.scala 76:24:@8928.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_3_idles; // @[sm_RootController.scala 76:24:@8928.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_4_cycs; // @[sm_RootController.scala 76:24:@8928.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_4_iters; // @[sm_RootController.scala 76:24:@8928.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_4_stalls; // @[sm_RootController.scala 76:24:@8928.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_4_idles; // @[sm_RootController.scala 76:24:@8928.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_5_cycs; // @[sm_RootController.scala 76:24:@8928.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_5_iters; // @[sm_RootController.scala 76:24:@8928.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_6_cycs; // @[sm_RootController.scala 76:24:@8928.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_6_iters; // @[sm_RootController.scala 76:24:@8928.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_6_stalls; // @[sm_RootController.scala 76:24:@8928.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_6_idles; // @[sm_RootController.scala 76:24:@8928.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_done; // @[sm_RootController.scala 76:24:@8928.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_baseEn; // @[sm_RootController.scala 76:24:@8928.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_RootController.scala 76:24:@8928.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0; // @[sm_RootController.scala 76:24:@8928.4]
  wire  RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[sm_RootController.scala 76:24:@8928.4]
  wire  RootController_kernelRootController_concrete1_io_rr; // @[sm_RootController.scala 76:24:@8928.4]
  wire  _T_745; // @[package.scala 96:25:@8788.4 package.scala 96:25:@8789.4]
  wire  _T_824; // @[Main.scala 36:50:@8865.4]
  wire  _T_825; // @[Main.scala 36:59:@8866.4]
  wire  _T_837; // @[package.scala 100:49:@8886.4]
  reg  _T_840; // @[package.scala 48:56:@8887.4]
  reg [31:0] _RAND_0;
  SingleCounter SingleCounter ( // @[Main.scala 29:32:@8765.4]
    .clock(SingleCounter_clock),
    .reset(SingleCounter_reset),
    .io_input_reset(SingleCounter_io_input_reset),
    .io_output_done(SingleCounter_io_output_done)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@8783.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  SRFF SRFF ( // @[Main.scala 34:28:@8799.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  RootController_sm RootController_sm ( // @[sm_RootController.scala 32:18:@8837.4]
    .clock(RootController_sm_clock),
    .reset(RootController_sm_reset),
    .io_enable(RootController_sm_io_enable),
    .io_done(RootController_sm_io_done),
    .io_rst(RootController_sm_io_rst),
    .io_ctrDone(RootController_sm_io_ctrDone),
    .io_ctrInc(RootController_sm_io_ctrInc),
    .io_doneIn_0(RootController_sm_io_doneIn_0),
    .io_enableOut_0(RootController_sm_io_enableOut_0),
    .io_childAck_0(RootController_sm_io_childAck_0)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@8869.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RootController_kernelRootController_concrete1 RootController_kernelRootController_concrete1 ( // @[sm_RootController.scala 76:24:@8928.4]
    .clock(RootController_kernelRootController_concrete1_clock),
    .reset(RootController_kernelRootController_concrete1_reset),
    .io_in_x95_TVALID(RootController_kernelRootController_concrete1_io_in_x95_TVALID),
    .io_in_x95_TREADY(RootController_kernelRootController_concrete1_io_in_x95_TREADY),
    .io_in_x95_TDATA(RootController_kernelRootController_concrete1_io_in_x95_TDATA),
    .io_in_x95_TSTRB(RootController_kernelRootController_concrete1_io_in_x95_TSTRB),
    .io_in_x95_TKEEP(RootController_kernelRootController_concrete1_io_in_x95_TKEEP),
    .io_in_x95_TLAST(RootController_kernelRootController_concrete1_io_in_x95_TLAST),
    .io_in_x95_TID(RootController_kernelRootController_concrete1_io_in_x95_TID),
    .io_in_x95_TDEST(RootController_kernelRootController_concrete1_io_in_x95_TDEST),
    .io_in_x95_TUSER(RootController_kernelRootController_concrete1_io_in_x95_TUSER),
    .io_in_x90_TVALID(RootController_kernelRootController_concrete1_io_in_x90_TVALID),
    .io_in_x90_TREADY(RootController_kernelRootController_concrete1_io_in_x90_TREADY),
    .io_in_x90_TDATA(RootController_kernelRootController_concrete1_io_in_x90_TDATA),
    .io_in_x90_TID(RootController_kernelRootController_concrete1_io_in_x90_TID),
    .io_in_x90_TDEST(RootController_kernelRootController_concrete1_io_in_x90_TDEST),
    .io_in_instrctrs_0_cycs(RootController_kernelRootController_concrete1_io_in_instrctrs_0_cycs),
    .io_in_instrctrs_0_iters(RootController_kernelRootController_concrete1_io_in_instrctrs_0_iters),
    .io_in_instrctrs_1_cycs(RootController_kernelRootController_concrete1_io_in_instrctrs_1_cycs),
    .io_in_instrctrs_1_iters(RootController_kernelRootController_concrete1_io_in_instrctrs_1_iters),
    .io_in_instrctrs_2_cycs(RootController_kernelRootController_concrete1_io_in_instrctrs_2_cycs),
    .io_in_instrctrs_2_iters(RootController_kernelRootController_concrete1_io_in_instrctrs_2_iters),
    .io_in_instrctrs_3_cycs(RootController_kernelRootController_concrete1_io_in_instrctrs_3_cycs),
    .io_in_instrctrs_3_iters(RootController_kernelRootController_concrete1_io_in_instrctrs_3_iters),
    .io_in_instrctrs_3_stalls(RootController_kernelRootController_concrete1_io_in_instrctrs_3_stalls),
    .io_in_instrctrs_3_idles(RootController_kernelRootController_concrete1_io_in_instrctrs_3_idles),
    .io_in_instrctrs_4_cycs(RootController_kernelRootController_concrete1_io_in_instrctrs_4_cycs),
    .io_in_instrctrs_4_iters(RootController_kernelRootController_concrete1_io_in_instrctrs_4_iters),
    .io_in_instrctrs_4_stalls(RootController_kernelRootController_concrete1_io_in_instrctrs_4_stalls),
    .io_in_instrctrs_4_idles(RootController_kernelRootController_concrete1_io_in_instrctrs_4_idles),
    .io_in_instrctrs_5_cycs(RootController_kernelRootController_concrete1_io_in_instrctrs_5_cycs),
    .io_in_instrctrs_5_iters(RootController_kernelRootController_concrete1_io_in_instrctrs_5_iters),
    .io_in_instrctrs_6_cycs(RootController_kernelRootController_concrete1_io_in_instrctrs_6_cycs),
    .io_in_instrctrs_6_iters(RootController_kernelRootController_concrete1_io_in_instrctrs_6_iters),
    .io_in_instrctrs_6_stalls(RootController_kernelRootController_concrete1_io_in_instrctrs_6_stalls),
    .io_in_instrctrs_6_idles(RootController_kernelRootController_concrete1_io_in_instrctrs_6_idles),
    .io_sigsIn_done(RootController_kernelRootController_concrete1_io_sigsIn_done),
    .io_sigsIn_baseEn(RootController_kernelRootController_concrete1_io_sigsIn_baseEn),
    .io_sigsIn_smEnableOuts_0(RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0),
    .io_rr(RootController_kernelRootController_concrete1_io_rr)
  );
  assign _T_745 = RetimeWrapper_io_out; // @[package.scala 96:25:@8788.4 package.scala 96:25:@8789.4]
  assign _T_824 = io_enable & _T_745; // @[Main.scala 36:50:@8865.4]
  assign _T_825 = ~ SRFF_io_output; // @[Main.scala 36:59:@8866.4]
  assign _T_837 = RootController_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@8886.4]
  assign io_done = SRFF_io_output; // @[Main.scala 43:23:@8885.4]
  assign io_memStreams_loads_0_cmd_valid = 1'h0;
  assign io_memStreams_loads_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_loads_0_cmd_bits_size = 32'h0;
  assign io_memStreams_loads_0_data_ready = 1'h0;
  assign io_memStreams_stores_0_cmd_valid = 1'h0;
  assign io_memStreams_stores_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_stores_0_cmd_bits_size = 32'h0;
  assign io_memStreams_stores_0_data_valid = 1'h0;
  assign io_memStreams_stores_0_data_bits_wdata_0 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_1 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_2 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_3 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_4 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_5 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_6 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_7 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_8 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_9 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_10 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_11 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_12 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_13 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_14 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_15 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wstrb = 16'h0;
  assign io_memStreams_stores_0_wresp_ready = 1'h0;
  assign io_memStreams_gathers_0_cmd_valid = 1'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_0 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_1 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_2 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_3 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_4 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_5 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_6 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_7 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_8 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_9 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_10 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_11 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_12 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_13 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_14 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_15 = 64'h0;
  assign io_memStreams_gathers_0_data_ready = 1'h0;
  assign io_memStreams_scatters_0_cmd_valid = 1'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_0 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_1 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_2 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_3 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_4 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_5 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_6 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_7 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_8 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_9 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_10 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_11 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_12 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_13 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_14 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_15 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_0 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_1 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_2 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_3 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_4 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_5 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_6 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_7 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_8 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_9 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_10 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_11 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_12 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_13 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_14 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_15 = 32'h0;
  assign io_memStreams_scatters_0_wresp_ready = 1'h0;
  assign io_axiStreamsIn_0_TREADY = RootController_kernelRootController_concrete1_io_in_x90_TREADY; // @[sm_RootController.scala 50:22:@9020.4]
  assign io_axiStreamsOut_0_TVALID = RootController_kernelRootController_concrete1_io_in_x95_TVALID; // @[sm_RootController.scala 49:22:@9012.4]
  assign io_axiStreamsOut_0_TDATA = RootController_kernelRootController_concrete1_io_in_x95_TDATA; // @[sm_RootController.scala 49:22:@9010.4]
  assign io_axiStreamsOut_0_TSTRB = RootController_kernelRootController_concrete1_io_in_x95_TSTRB; // @[sm_RootController.scala 49:22:@9009.4]
  assign io_axiStreamsOut_0_TKEEP = RootController_kernelRootController_concrete1_io_in_x95_TKEEP; // @[sm_RootController.scala 49:22:@9008.4]
  assign io_axiStreamsOut_0_TLAST = RootController_kernelRootController_concrete1_io_in_x95_TLAST; // @[sm_RootController.scala 49:22:@9007.4]
  assign io_axiStreamsOut_0_TID = RootController_kernelRootController_concrete1_io_in_x95_TID; // @[sm_RootController.scala 49:22:@9006.4]
  assign io_axiStreamsOut_0_TDEST = RootController_kernelRootController_concrete1_io_in_x95_TDEST; // @[sm_RootController.scala 49:22:@9005.4]
  assign io_axiStreamsOut_0_TUSER = RootController_kernelRootController_concrete1_io_in_x95_TUSER; // @[sm_RootController.scala 49:22:@9004.4]
  assign io_heap_0_req_valid = 1'h0;
  assign io_heap_0_req_bits_allocDealloc = 1'h0;
  assign io_heap_0_req_bits_sizeAddr = 64'h0;
  assign io_argOuts_0_port_valid = io_enable; // @[Instrument.scala 27:57:@9078.4]
  assign io_argOuts_0_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_0_cycs; // @[Instrument.scala 26:56:@9077.4]
  assign io_argOuts_1_port_valid = io_enable; // @[Instrument.scala 29:56:@9080.4]
  assign io_argOuts_1_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_0_iters; // @[Instrument.scala 28:55:@9079.4]
  assign io_argOuts_2_port_valid = io_enable; // @[Instrument.scala 31:58:@9082.4]
  assign io_argOuts_2_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_1_cycs; // @[Instrument.scala 30:57:@9081.4]
  assign io_argOuts_3_port_valid = io_enable; // @[Instrument.scala 33:57:@9084.4]
  assign io_argOuts_3_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_1_iters; // @[Instrument.scala 32:56:@9083.4]
  assign io_argOuts_4_port_valid = io_enable; // @[Instrument.scala 35:58:@9086.4]
  assign io_argOuts_4_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_2_cycs; // @[Instrument.scala 34:57:@9085.4]
  assign io_argOuts_5_port_valid = io_enable; // @[Instrument.scala 37:57:@9088.4]
  assign io_argOuts_5_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_2_iters; // @[Instrument.scala 36:56:@9087.4]
  assign io_argOuts_6_port_valid = io_enable; // @[Instrument.scala 39:58:@9090.4]
  assign io_argOuts_6_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_3_cycs; // @[Instrument.scala 38:57:@9089.4]
  assign io_argOuts_7_port_valid = io_enable; // @[Instrument.scala 41:57:@9092.4]
  assign io_argOuts_7_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_3_iters; // @[Instrument.scala 40:56:@9091.4]
  assign io_argOuts_8_port_valid = io_enable; // @[Instrument.scala 43:59:@9094.4]
  assign io_argOuts_8_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_3_stalls; // @[Instrument.scala 42:58:@9093.4]
  assign io_argOuts_9_port_valid = io_enable; // @[Instrument.scala 45:56:@9096.4]
  assign io_argOuts_9_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_3_idles; // @[Instrument.scala 44:55:@9095.4]
  assign io_argOuts_10_port_valid = io_enable; // @[Instrument.scala 47:58:@9098.4]
  assign io_argOuts_10_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_4_cycs; // @[Instrument.scala 46:57:@9097.4]
  assign io_argOuts_11_port_valid = io_enable; // @[Instrument.scala 49:57:@9100.4]
  assign io_argOuts_11_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_4_iters; // @[Instrument.scala 48:56:@9099.4]
  assign io_argOuts_12_port_valid = io_enable; // @[Instrument.scala 51:59:@9102.4]
  assign io_argOuts_12_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_4_stalls; // @[Instrument.scala 50:58:@9101.4]
  assign io_argOuts_13_port_valid = io_enable; // @[Instrument.scala 53:56:@9104.4]
  assign io_argOuts_13_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_4_idles; // @[Instrument.scala 52:55:@9103.4]
  assign io_argOuts_14_port_valid = io_enable; // @[Instrument.scala 55:58:@9106.4]
  assign io_argOuts_14_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_5_cycs; // @[Instrument.scala 54:57:@9105.4]
  assign io_argOuts_15_port_valid = io_enable; // @[Instrument.scala 57:57:@9108.4]
  assign io_argOuts_15_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_5_iters; // @[Instrument.scala 56:56:@9107.4]
  assign io_argOuts_16_port_valid = io_enable; // @[Instrument.scala 59:58:@9110.4]
  assign io_argOuts_16_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_6_cycs; // @[Instrument.scala 58:57:@9109.4]
  assign io_argOuts_17_port_valid = io_enable; // @[Instrument.scala 61:57:@9112.4]
  assign io_argOuts_17_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_6_iters; // @[Instrument.scala 60:56:@9111.4]
  assign io_argOuts_18_port_valid = io_enable; // @[Instrument.scala 63:59:@9114.4]
  assign io_argOuts_18_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_6_stalls; // @[Instrument.scala 62:58:@9113.4]
  assign io_argOuts_19_port_valid = io_enable; // @[Instrument.scala 65:56:@9116.4]
  assign io_argOuts_19_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_6_idles; // @[Instrument.scala 64:55:@9115.4]
  assign SingleCounter_clock = clock; // @[:@8766.4]
  assign SingleCounter_reset = reset; // @[:@8767.4]
  assign SingleCounter_io_input_reset = reset; // @[Main.scala 30:79:@8781.4]
  assign RetimeWrapper_clock = clock; // @[:@8784.4]
  assign RetimeWrapper_reset = reset; // @[:@8785.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@8787.4]
  assign RetimeWrapper_io_in = SingleCounter_io_output_done; // @[package.scala 94:16:@8786.4]
  assign SRFF_clock = clock; // @[:@8800.4]
  assign SRFF_reset = reset; // @[:@8801.4]
  assign SRFF_io_input_set = RootController_sm_io_done; // @[Main.scala 52:29:@9076.4]
  assign SRFF_io_input_reset = RetimeWrapper_1_io_out; // @[Main.scala 41:31:@8883.4]
  assign SRFF_io_input_asyn_reset = RetimeWrapper_1_io_out; // @[Main.scala 42:36:@8884.4]
  assign RootController_sm_clock = clock; // @[:@8838.4]
  assign RootController_sm_reset = reset; // @[:@8839.4]
  assign RootController_sm_io_enable = _T_824 & _T_825; // @[Main.scala 40:33:@8882.4 SpatialBlocks.scala 112:18:@8916.4]
  assign RootController_sm_io_rst = RetimeWrapper_1_io_out; // @[SpatialBlocks.scala 106:15:@8910.4]
  assign RootController_sm_io_ctrDone = RootController_sm_io_ctrInc & _T_840; // @[Main.scala 44:34:@8890.4]
  assign RootController_sm_io_doneIn_0 = RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 102:67:@8907.4]
  assign RetimeWrapper_1_clock = clock; // @[:@8870.4]
  assign RetimeWrapper_1_reset = reset; // @[:@8871.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@8873.4]
  assign RetimeWrapper_1_io_in = reset | io_reset; // @[package.scala 94:16:@8872.4]
  assign RootController_kernelRootController_concrete1_clock = clock; // @[:@8929.4]
  assign RootController_kernelRootController_concrete1_reset = reset; // @[:@8930.4]
  assign RootController_kernelRootController_concrete1_io_in_x95_TREADY = io_axiStreamsOut_0_TREADY; // @[sm_RootController.scala 49:22:@9011.4]
  assign RootController_kernelRootController_concrete1_io_in_x90_TVALID = io_axiStreamsIn_0_TVALID; // @[sm_RootController.scala 50:22:@9021.4]
  assign RootController_kernelRootController_concrete1_io_in_x90_TDATA = io_axiStreamsIn_0_TDATA; // @[sm_RootController.scala 50:22:@9019.4]
  assign RootController_kernelRootController_concrete1_io_in_x90_TID = io_axiStreamsIn_0_TID; // @[sm_RootController.scala 50:22:@9015.4]
  assign RootController_kernelRootController_concrete1_io_in_x90_TDEST = io_axiStreamsIn_0_TDEST; // @[sm_RootController.scala 50:22:@9014.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_done = RootController_sm_io_done; // @[sm_RootController.scala 81:22:@9068.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_baseEn = _T_824 & _T_825; // @[sm_RootController.scala 81:22:@9061.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0 = RootController_sm_io_enableOut_0; // @[sm_RootController.scala 81:22:@9058.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0 = RootController_sm_io_childAck_0; // @[sm_RootController.scala 81:22:@9056.4]
  assign RootController_kernelRootController_concrete1_io_rr = RetimeWrapper_io_out; // @[sm_RootController.scala 80:18:@9050.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_840 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_840 <= 1'h0;
    end else begin
      _T_840 <= _T_837;
    end
  end
endmodule
module DRAMHeap( // @[:@10023.2]
  input         io_accel_0_req_valid, // @[:@10026.4]
  input         io_accel_0_req_bits_allocDealloc, // @[:@10026.4]
  input  [63:0] io_accel_0_req_bits_sizeAddr, // @[:@10026.4]
  output        io_accel_0_resp_valid, // @[:@10026.4]
  output        io_accel_0_resp_bits_allocDealloc, // @[:@10026.4]
  output [63:0] io_accel_0_resp_bits_sizeAddr, // @[:@10026.4]
  output        io_host_0_req_valid, // @[:@10026.4]
  output        io_host_0_req_bits_allocDealloc, // @[:@10026.4]
  output [63:0] io_host_0_req_bits_sizeAddr, // @[:@10026.4]
  input         io_host_0_resp_valid, // @[:@10026.4]
  input         io_host_0_resp_bits_allocDealloc, // @[:@10026.4]
  input  [63:0] io_host_0_resp_bits_sizeAddr // @[:@10026.4]
);
  assign io_accel_0_resp_valid = io_host_0_resp_valid; // @[DRAMHeap.scala 24:18:@10033.4]
  assign io_accel_0_resp_bits_allocDealloc = io_host_0_resp_bits_allocDealloc; // @[DRAMHeap.scala 25:17:@10035.4]
  assign io_accel_0_resp_bits_sizeAddr = io_host_0_resp_bits_sizeAddr; // @[DRAMHeap.scala 25:17:@10034.4]
  assign io_host_0_req_valid = io_accel_0_req_valid; // @[DRAMHeap.scala 21:18:@10030.4]
  assign io_host_0_req_bits_allocDealloc = io_accel_0_req_bits_allocDealloc; // @[DRAMHeap.scala 21:18:@10029.4]
  assign io_host_0_req_bits_sizeAddr = io_accel_0_req_bits_sizeAddr; // @[DRAMHeap.scala 21:18:@10028.4]
endmodule
module RetimeWrapper_68( // @[:@10049.2]
  input         clock, // @[:@10050.4]
  input         reset, // @[:@10051.4]
  input         io_flow, // @[:@10052.4]
  input  [63:0] io_in, // @[:@10052.4]
  output [63:0] io_out // @[:@10052.4]
);
  wire [63:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@10054.4]
  wire [63:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@10054.4]
  wire [63:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@10054.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@10054.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@10054.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@10054.4]
  RetimeShiftRegister #(.WIDTH(64), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@10054.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@10067.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@10066.4]
  assign sr_init = 64'h0; // @[RetimeShiftRegister.scala 19:16:@10065.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@10064.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@10063.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@10061.4]
endmodule
module FringeFF( // @[:@10069.2]
  input         clock, // @[:@10070.4]
  input         reset, // @[:@10071.4]
  input  [63:0] io_in, // @[:@10072.4]
  input         io_reset, // @[:@10072.4]
  output [63:0] io_out, // @[:@10072.4]
  input         io_enable // @[:@10072.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@10075.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@10075.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@10075.4]
  wire [63:0] RetimeWrapper_io_in; // @[package.scala 93:22:@10075.4]
  wire [63:0] RetimeWrapper_io_out; // @[package.scala 93:22:@10075.4]
  wire [63:0] _T_18; // @[package.scala 96:25:@10080.4 package.scala 96:25:@10081.4]
  wire [63:0] _GEN_0; // @[FringeFF.scala 21:27:@10086.6]
  RetimeWrapper_68 RetimeWrapper ( // @[package.scala 93:22:@10075.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@10080.4 package.scala 96:25:@10081.4]
  assign _GEN_0 = io_reset ? 64'h0 : _T_18; // @[FringeFF.scala 21:27:@10086.6]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@10092.4]
  assign RetimeWrapper_clock = clock; // @[:@10076.4]
  assign RetimeWrapper_reset = reset; // @[:@10077.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@10079.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _GEN_0; // @[package.scala 94:16:@10078.4]
endmodule
module MuxN( // @[:@39791.2]
  input  [63:0] io_ins_0, // @[:@39794.4]
  input  [63:0] io_ins_1, // @[:@39794.4]
  input  [63:0] io_ins_2, // @[:@39794.4]
  input  [63:0] io_ins_3, // @[:@39794.4]
  input  [63:0] io_ins_4, // @[:@39794.4]
  input  [63:0] io_ins_5, // @[:@39794.4]
  input  [63:0] io_ins_6, // @[:@39794.4]
  input  [63:0] io_ins_7, // @[:@39794.4]
  input  [63:0] io_ins_8, // @[:@39794.4]
  input  [63:0] io_ins_9, // @[:@39794.4]
  input  [63:0] io_ins_10, // @[:@39794.4]
  input  [63:0] io_ins_11, // @[:@39794.4]
  input  [63:0] io_ins_12, // @[:@39794.4]
  input  [63:0] io_ins_13, // @[:@39794.4]
  input  [63:0] io_ins_14, // @[:@39794.4]
  input  [63:0] io_ins_15, // @[:@39794.4]
  input  [63:0] io_ins_16, // @[:@39794.4]
  input  [63:0] io_ins_17, // @[:@39794.4]
  input  [63:0] io_ins_18, // @[:@39794.4]
  input  [63:0] io_ins_19, // @[:@39794.4]
  input  [63:0] io_ins_20, // @[:@39794.4]
  input  [63:0] io_ins_21, // @[:@39794.4]
  input  [63:0] io_ins_22, // @[:@39794.4]
  input  [63:0] io_ins_23, // @[:@39794.4]
  input  [63:0] io_ins_24, // @[:@39794.4]
  input  [63:0] io_ins_25, // @[:@39794.4]
  input  [63:0] io_ins_26, // @[:@39794.4]
  input  [63:0] io_ins_27, // @[:@39794.4]
  input  [63:0] io_ins_28, // @[:@39794.4]
  input  [63:0] io_ins_29, // @[:@39794.4]
  input  [63:0] io_ins_30, // @[:@39794.4]
  input  [63:0] io_ins_31, // @[:@39794.4]
  input  [63:0] io_ins_32, // @[:@39794.4]
  input  [63:0] io_ins_33, // @[:@39794.4]
  input  [63:0] io_ins_34, // @[:@39794.4]
  input  [63:0] io_ins_35, // @[:@39794.4]
  input  [63:0] io_ins_36, // @[:@39794.4]
  input  [63:0] io_ins_37, // @[:@39794.4]
  input  [63:0] io_ins_38, // @[:@39794.4]
  input  [63:0] io_ins_39, // @[:@39794.4]
  input  [63:0] io_ins_40, // @[:@39794.4]
  input  [63:0] io_ins_41, // @[:@39794.4]
  input  [63:0] io_ins_42, // @[:@39794.4]
  input  [63:0] io_ins_43, // @[:@39794.4]
  input  [63:0] io_ins_44, // @[:@39794.4]
  input  [63:0] io_ins_45, // @[:@39794.4]
  input  [63:0] io_ins_46, // @[:@39794.4]
  input  [63:0] io_ins_47, // @[:@39794.4]
  input  [63:0] io_ins_48, // @[:@39794.4]
  input  [63:0] io_ins_49, // @[:@39794.4]
  input  [63:0] io_ins_50, // @[:@39794.4]
  input  [63:0] io_ins_51, // @[:@39794.4]
  input  [63:0] io_ins_52, // @[:@39794.4]
  input  [63:0] io_ins_53, // @[:@39794.4]
  input  [63:0] io_ins_54, // @[:@39794.4]
  input  [63:0] io_ins_55, // @[:@39794.4]
  input  [63:0] io_ins_56, // @[:@39794.4]
  input  [63:0] io_ins_57, // @[:@39794.4]
  input  [63:0] io_ins_58, // @[:@39794.4]
  input  [63:0] io_ins_59, // @[:@39794.4]
  input  [63:0] io_ins_60, // @[:@39794.4]
  input  [63:0] io_ins_61, // @[:@39794.4]
  input  [63:0] io_ins_62, // @[:@39794.4]
  input  [63:0] io_ins_63, // @[:@39794.4]
  input  [63:0] io_ins_64, // @[:@39794.4]
  input  [63:0] io_ins_65, // @[:@39794.4]
  input  [63:0] io_ins_66, // @[:@39794.4]
  input  [63:0] io_ins_67, // @[:@39794.4]
  input  [63:0] io_ins_68, // @[:@39794.4]
  input  [63:0] io_ins_69, // @[:@39794.4]
  input  [63:0] io_ins_70, // @[:@39794.4]
  input  [63:0] io_ins_71, // @[:@39794.4]
  input  [63:0] io_ins_72, // @[:@39794.4]
  input  [63:0] io_ins_73, // @[:@39794.4]
  input  [63:0] io_ins_74, // @[:@39794.4]
  input  [63:0] io_ins_75, // @[:@39794.4]
  input  [63:0] io_ins_76, // @[:@39794.4]
  input  [63:0] io_ins_77, // @[:@39794.4]
  input  [63:0] io_ins_78, // @[:@39794.4]
  input  [63:0] io_ins_79, // @[:@39794.4]
  input  [63:0] io_ins_80, // @[:@39794.4]
  input  [63:0] io_ins_81, // @[:@39794.4]
  input  [63:0] io_ins_82, // @[:@39794.4]
  input  [63:0] io_ins_83, // @[:@39794.4]
  input  [63:0] io_ins_84, // @[:@39794.4]
  input  [63:0] io_ins_85, // @[:@39794.4]
  input  [63:0] io_ins_86, // @[:@39794.4]
  input  [63:0] io_ins_87, // @[:@39794.4]
  input  [63:0] io_ins_88, // @[:@39794.4]
  input  [63:0] io_ins_89, // @[:@39794.4]
  input  [63:0] io_ins_90, // @[:@39794.4]
  input  [63:0] io_ins_91, // @[:@39794.4]
  input  [63:0] io_ins_92, // @[:@39794.4]
  input  [63:0] io_ins_93, // @[:@39794.4]
  input  [63:0] io_ins_94, // @[:@39794.4]
  input  [63:0] io_ins_95, // @[:@39794.4]
  input  [63:0] io_ins_96, // @[:@39794.4]
  input  [63:0] io_ins_97, // @[:@39794.4]
  input  [63:0] io_ins_98, // @[:@39794.4]
  input  [63:0] io_ins_99, // @[:@39794.4]
  input  [63:0] io_ins_100, // @[:@39794.4]
  input  [63:0] io_ins_101, // @[:@39794.4]
  input  [63:0] io_ins_102, // @[:@39794.4]
  input  [63:0] io_ins_103, // @[:@39794.4]
  input  [63:0] io_ins_104, // @[:@39794.4]
  input  [63:0] io_ins_105, // @[:@39794.4]
  input  [63:0] io_ins_106, // @[:@39794.4]
  input  [63:0] io_ins_107, // @[:@39794.4]
  input  [63:0] io_ins_108, // @[:@39794.4]
  input  [63:0] io_ins_109, // @[:@39794.4]
  input  [63:0] io_ins_110, // @[:@39794.4]
  input  [63:0] io_ins_111, // @[:@39794.4]
  input  [63:0] io_ins_112, // @[:@39794.4]
  input  [63:0] io_ins_113, // @[:@39794.4]
  input  [63:0] io_ins_114, // @[:@39794.4]
  input  [63:0] io_ins_115, // @[:@39794.4]
  input  [63:0] io_ins_116, // @[:@39794.4]
  input  [63:0] io_ins_117, // @[:@39794.4]
  input  [63:0] io_ins_118, // @[:@39794.4]
  input  [63:0] io_ins_119, // @[:@39794.4]
  input  [63:0] io_ins_120, // @[:@39794.4]
  input  [63:0] io_ins_121, // @[:@39794.4]
  input  [63:0] io_ins_122, // @[:@39794.4]
  input  [63:0] io_ins_123, // @[:@39794.4]
  input  [63:0] io_ins_124, // @[:@39794.4]
  input  [63:0] io_ins_125, // @[:@39794.4]
  input  [63:0] io_ins_126, // @[:@39794.4]
  input  [63:0] io_ins_127, // @[:@39794.4]
  input  [63:0] io_ins_128, // @[:@39794.4]
  input  [63:0] io_ins_129, // @[:@39794.4]
  input  [63:0] io_ins_130, // @[:@39794.4]
  input  [63:0] io_ins_131, // @[:@39794.4]
  input  [63:0] io_ins_132, // @[:@39794.4]
  input  [63:0] io_ins_133, // @[:@39794.4]
  input  [63:0] io_ins_134, // @[:@39794.4]
  input  [63:0] io_ins_135, // @[:@39794.4]
  input  [63:0] io_ins_136, // @[:@39794.4]
  input  [63:0] io_ins_137, // @[:@39794.4]
  input  [63:0] io_ins_138, // @[:@39794.4]
  input  [63:0] io_ins_139, // @[:@39794.4]
  input  [63:0] io_ins_140, // @[:@39794.4]
  input  [63:0] io_ins_141, // @[:@39794.4]
  input  [63:0] io_ins_142, // @[:@39794.4]
  input  [63:0] io_ins_143, // @[:@39794.4]
  input  [63:0] io_ins_144, // @[:@39794.4]
  input  [63:0] io_ins_145, // @[:@39794.4]
  input  [63:0] io_ins_146, // @[:@39794.4]
  input  [63:0] io_ins_147, // @[:@39794.4]
  input  [63:0] io_ins_148, // @[:@39794.4]
  input  [63:0] io_ins_149, // @[:@39794.4]
  input  [63:0] io_ins_150, // @[:@39794.4]
  input  [63:0] io_ins_151, // @[:@39794.4]
  input  [63:0] io_ins_152, // @[:@39794.4]
  input  [63:0] io_ins_153, // @[:@39794.4]
  input  [63:0] io_ins_154, // @[:@39794.4]
  input  [63:0] io_ins_155, // @[:@39794.4]
  input  [63:0] io_ins_156, // @[:@39794.4]
  input  [63:0] io_ins_157, // @[:@39794.4]
  input  [63:0] io_ins_158, // @[:@39794.4]
  input  [63:0] io_ins_159, // @[:@39794.4]
  input  [63:0] io_ins_160, // @[:@39794.4]
  input  [63:0] io_ins_161, // @[:@39794.4]
  input  [63:0] io_ins_162, // @[:@39794.4]
  input  [63:0] io_ins_163, // @[:@39794.4]
  input  [63:0] io_ins_164, // @[:@39794.4]
  input  [63:0] io_ins_165, // @[:@39794.4]
  input  [63:0] io_ins_166, // @[:@39794.4]
  input  [63:0] io_ins_167, // @[:@39794.4]
  input  [63:0] io_ins_168, // @[:@39794.4]
  input  [63:0] io_ins_169, // @[:@39794.4]
  input  [63:0] io_ins_170, // @[:@39794.4]
  input  [63:0] io_ins_171, // @[:@39794.4]
  input  [63:0] io_ins_172, // @[:@39794.4]
  input  [63:0] io_ins_173, // @[:@39794.4]
  input  [63:0] io_ins_174, // @[:@39794.4]
  input  [63:0] io_ins_175, // @[:@39794.4]
  input  [63:0] io_ins_176, // @[:@39794.4]
  input  [63:0] io_ins_177, // @[:@39794.4]
  input  [63:0] io_ins_178, // @[:@39794.4]
  input  [63:0] io_ins_179, // @[:@39794.4]
  input  [63:0] io_ins_180, // @[:@39794.4]
  input  [63:0] io_ins_181, // @[:@39794.4]
  input  [63:0] io_ins_182, // @[:@39794.4]
  input  [63:0] io_ins_183, // @[:@39794.4]
  input  [63:0] io_ins_184, // @[:@39794.4]
  input  [63:0] io_ins_185, // @[:@39794.4]
  input  [63:0] io_ins_186, // @[:@39794.4]
  input  [63:0] io_ins_187, // @[:@39794.4]
  input  [63:0] io_ins_188, // @[:@39794.4]
  input  [63:0] io_ins_189, // @[:@39794.4]
  input  [63:0] io_ins_190, // @[:@39794.4]
  input  [63:0] io_ins_191, // @[:@39794.4]
  input  [63:0] io_ins_192, // @[:@39794.4]
  input  [63:0] io_ins_193, // @[:@39794.4]
  input  [63:0] io_ins_194, // @[:@39794.4]
  input  [63:0] io_ins_195, // @[:@39794.4]
  input  [63:0] io_ins_196, // @[:@39794.4]
  input  [63:0] io_ins_197, // @[:@39794.4]
  input  [63:0] io_ins_198, // @[:@39794.4]
  input  [63:0] io_ins_199, // @[:@39794.4]
  input  [63:0] io_ins_200, // @[:@39794.4]
  input  [63:0] io_ins_201, // @[:@39794.4]
  input  [63:0] io_ins_202, // @[:@39794.4]
  input  [63:0] io_ins_203, // @[:@39794.4]
  input  [63:0] io_ins_204, // @[:@39794.4]
  input  [63:0] io_ins_205, // @[:@39794.4]
  input  [63:0] io_ins_206, // @[:@39794.4]
  input  [63:0] io_ins_207, // @[:@39794.4]
  input  [63:0] io_ins_208, // @[:@39794.4]
  input  [63:0] io_ins_209, // @[:@39794.4]
  input  [63:0] io_ins_210, // @[:@39794.4]
  input  [63:0] io_ins_211, // @[:@39794.4]
  input  [63:0] io_ins_212, // @[:@39794.4]
  input  [63:0] io_ins_213, // @[:@39794.4]
  input  [63:0] io_ins_214, // @[:@39794.4]
  input  [63:0] io_ins_215, // @[:@39794.4]
  input  [63:0] io_ins_216, // @[:@39794.4]
  input  [63:0] io_ins_217, // @[:@39794.4]
  input  [63:0] io_ins_218, // @[:@39794.4]
  input  [63:0] io_ins_219, // @[:@39794.4]
  input  [63:0] io_ins_220, // @[:@39794.4]
  input  [63:0] io_ins_221, // @[:@39794.4]
  input  [63:0] io_ins_222, // @[:@39794.4]
  input  [63:0] io_ins_223, // @[:@39794.4]
  input  [63:0] io_ins_224, // @[:@39794.4]
  input  [63:0] io_ins_225, // @[:@39794.4]
  input  [63:0] io_ins_226, // @[:@39794.4]
  input  [63:0] io_ins_227, // @[:@39794.4]
  input  [63:0] io_ins_228, // @[:@39794.4]
  input  [63:0] io_ins_229, // @[:@39794.4]
  input  [63:0] io_ins_230, // @[:@39794.4]
  input  [63:0] io_ins_231, // @[:@39794.4]
  input  [63:0] io_ins_232, // @[:@39794.4]
  input  [63:0] io_ins_233, // @[:@39794.4]
  input  [63:0] io_ins_234, // @[:@39794.4]
  input  [63:0] io_ins_235, // @[:@39794.4]
  input  [63:0] io_ins_236, // @[:@39794.4]
  input  [63:0] io_ins_237, // @[:@39794.4]
  input  [63:0] io_ins_238, // @[:@39794.4]
  input  [63:0] io_ins_239, // @[:@39794.4]
  input  [63:0] io_ins_240, // @[:@39794.4]
  input  [63:0] io_ins_241, // @[:@39794.4]
  input  [63:0] io_ins_242, // @[:@39794.4]
  input  [63:0] io_ins_243, // @[:@39794.4]
  input  [63:0] io_ins_244, // @[:@39794.4]
  input  [63:0] io_ins_245, // @[:@39794.4]
  input  [63:0] io_ins_246, // @[:@39794.4]
  input  [63:0] io_ins_247, // @[:@39794.4]
  input  [63:0] io_ins_248, // @[:@39794.4]
  input  [63:0] io_ins_249, // @[:@39794.4]
  input  [63:0] io_ins_250, // @[:@39794.4]
  input  [63:0] io_ins_251, // @[:@39794.4]
  input  [63:0] io_ins_252, // @[:@39794.4]
  input  [63:0] io_ins_253, // @[:@39794.4]
  input  [63:0] io_ins_254, // @[:@39794.4]
  input  [63:0] io_ins_255, // @[:@39794.4]
  input  [63:0] io_ins_256, // @[:@39794.4]
  input  [63:0] io_ins_257, // @[:@39794.4]
  input  [63:0] io_ins_258, // @[:@39794.4]
  input  [63:0] io_ins_259, // @[:@39794.4]
  input  [63:0] io_ins_260, // @[:@39794.4]
  input  [63:0] io_ins_261, // @[:@39794.4]
  input  [63:0] io_ins_262, // @[:@39794.4]
  input  [63:0] io_ins_263, // @[:@39794.4]
  input  [63:0] io_ins_264, // @[:@39794.4]
  input  [63:0] io_ins_265, // @[:@39794.4]
  input  [63:0] io_ins_266, // @[:@39794.4]
  input  [63:0] io_ins_267, // @[:@39794.4]
  input  [63:0] io_ins_268, // @[:@39794.4]
  input  [63:0] io_ins_269, // @[:@39794.4]
  input  [63:0] io_ins_270, // @[:@39794.4]
  input  [63:0] io_ins_271, // @[:@39794.4]
  input  [63:0] io_ins_272, // @[:@39794.4]
  input  [63:0] io_ins_273, // @[:@39794.4]
  input  [63:0] io_ins_274, // @[:@39794.4]
  input  [63:0] io_ins_275, // @[:@39794.4]
  input  [63:0] io_ins_276, // @[:@39794.4]
  input  [63:0] io_ins_277, // @[:@39794.4]
  input  [63:0] io_ins_278, // @[:@39794.4]
  input  [63:0] io_ins_279, // @[:@39794.4]
  input  [63:0] io_ins_280, // @[:@39794.4]
  input  [63:0] io_ins_281, // @[:@39794.4]
  input  [63:0] io_ins_282, // @[:@39794.4]
  input  [63:0] io_ins_283, // @[:@39794.4]
  input  [63:0] io_ins_284, // @[:@39794.4]
  input  [63:0] io_ins_285, // @[:@39794.4]
  input  [63:0] io_ins_286, // @[:@39794.4]
  input  [63:0] io_ins_287, // @[:@39794.4]
  input  [63:0] io_ins_288, // @[:@39794.4]
  input  [63:0] io_ins_289, // @[:@39794.4]
  input  [63:0] io_ins_290, // @[:@39794.4]
  input  [63:0] io_ins_291, // @[:@39794.4]
  input  [63:0] io_ins_292, // @[:@39794.4]
  input  [63:0] io_ins_293, // @[:@39794.4]
  input  [63:0] io_ins_294, // @[:@39794.4]
  input  [63:0] io_ins_295, // @[:@39794.4]
  input  [63:0] io_ins_296, // @[:@39794.4]
  input  [63:0] io_ins_297, // @[:@39794.4]
  input  [63:0] io_ins_298, // @[:@39794.4]
  input  [63:0] io_ins_299, // @[:@39794.4]
  input  [63:0] io_ins_300, // @[:@39794.4]
  input  [63:0] io_ins_301, // @[:@39794.4]
  input  [63:0] io_ins_302, // @[:@39794.4]
  input  [63:0] io_ins_303, // @[:@39794.4]
  input  [63:0] io_ins_304, // @[:@39794.4]
  input  [63:0] io_ins_305, // @[:@39794.4]
  input  [63:0] io_ins_306, // @[:@39794.4]
  input  [63:0] io_ins_307, // @[:@39794.4]
  input  [63:0] io_ins_308, // @[:@39794.4]
  input  [63:0] io_ins_309, // @[:@39794.4]
  input  [63:0] io_ins_310, // @[:@39794.4]
  input  [63:0] io_ins_311, // @[:@39794.4]
  input  [63:0] io_ins_312, // @[:@39794.4]
  input  [63:0] io_ins_313, // @[:@39794.4]
  input  [63:0] io_ins_314, // @[:@39794.4]
  input  [63:0] io_ins_315, // @[:@39794.4]
  input  [63:0] io_ins_316, // @[:@39794.4]
  input  [63:0] io_ins_317, // @[:@39794.4]
  input  [63:0] io_ins_318, // @[:@39794.4]
  input  [63:0] io_ins_319, // @[:@39794.4]
  input  [63:0] io_ins_320, // @[:@39794.4]
  input  [63:0] io_ins_321, // @[:@39794.4]
  input  [63:0] io_ins_322, // @[:@39794.4]
  input  [63:0] io_ins_323, // @[:@39794.4]
  input  [63:0] io_ins_324, // @[:@39794.4]
  input  [63:0] io_ins_325, // @[:@39794.4]
  input  [63:0] io_ins_326, // @[:@39794.4]
  input  [63:0] io_ins_327, // @[:@39794.4]
  input  [63:0] io_ins_328, // @[:@39794.4]
  input  [63:0] io_ins_329, // @[:@39794.4]
  input  [63:0] io_ins_330, // @[:@39794.4]
  input  [63:0] io_ins_331, // @[:@39794.4]
  input  [63:0] io_ins_332, // @[:@39794.4]
  input  [63:0] io_ins_333, // @[:@39794.4]
  input  [63:0] io_ins_334, // @[:@39794.4]
  input  [63:0] io_ins_335, // @[:@39794.4]
  input  [63:0] io_ins_336, // @[:@39794.4]
  input  [63:0] io_ins_337, // @[:@39794.4]
  input  [63:0] io_ins_338, // @[:@39794.4]
  input  [63:0] io_ins_339, // @[:@39794.4]
  input  [63:0] io_ins_340, // @[:@39794.4]
  input  [63:0] io_ins_341, // @[:@39794.4]
  input  [63:0] io_ins_342, // @[:@39794.4]
  input  [63:0] io_ins_343, // @[:@39794.4]
  input  [63:0] io_ins_344, // @[:@39794.4]
  input  [63:0] io_ins_345, // @[:@39794.4]
  input  [63:0] io_ins_346, // @[:@39794.4]
  input  [63:0] io_ins_347, // @[:@39794.4]
  input  [63:0] io_ins_348, // @[:@39794.4]
  input  [63:0] io_ins_349, // @[:@39794.4]
  input  [63:0] io_ins_350, // @[:@39794.4]
  input  [63:0] io_ins_351, // @[:@39794.4]
  input  [63:0] io_ins_352, // @[:@39794.4]
  input  [63:0] io_ins_353, // @[:@39794.4]
  input  [63:0] io_ins_354, // @[:@39794.4]
  input  [63:0] io_ins_355, // @[:@39794.4]
  input  [63:0] io_ins_356, // @[:@39794.4]
  input  [63:0] io_ins_357, // @[:@39794.4]
  input  [63:0] io_ins_358, // @[:@39794.4]
  input  [63:0] io_ins_359, // @[:@39794.4]
  input  [63:0] io_ins_360, // @[:@39794.4]
  input  [63:0] io_ins_361, // @[:@39794.4]
  input  [63:0] io_ins_362, // @[:@39794.4]
  input  [63:0] io_ins_363, // @[:@39794.4]
  input  [63:0] io_ins_364, // @[:@39794.4]
  input  [63:0] io_ins_365, // @[:@39794.4]
  input  [63:0] io_ins_366, // @[:@39794.4]
  input  [63:0] io_ins_367, // @[:@39794.4]
  input  [63:0] io_ins_368, // @[:@39794.4]
  input  [63:0] io_ins_369, // @[:@39794.4]
  input  [63:0] io_ins_370, // @[:@39794.4]
  input  [63:0] io_ins_371, // @[:@39794.4]
  input  [63:0] io_ins_372, // @[:@39794.4]
  input  [63:0] io_ins_373, // @[:@39794.4]
  input  [63:0] io_ins_374, // @[:@39794.4]
  input  [63:0] io_ins_375, // @[:@39794.4]
  input  [63:0] io_ins_376, // @[:@39794.4]
  input  [63:0] io_ins_377, // @[:@39794.4]
  input  [63:0] io_ins_378, // @[:@39794.4]
  input  [63:0] io_ins_379, // @[:@39794.4]
  input  [63:0] io_ins_380, // @[:@39794.4]
  input  [63:0] io_ins_381, // @[:@39794.4]
  input  [63:0] io_ins_382, // @[:@39794.4]
  input  [63:0] io_ins_383, // @[:@39794.4]
  input  [63:0] io_ins_384, // @[:@39794.4]
  input  [63:0] io_ins_385, // @[:@39794.4]
  input  [63:0] io_ins_386, // @[:@39794.4]
  input  [63:0] io_ins_387, // @[:@39794.4]
  input  [63:0] io_ins_388, // @[:@39794.4]
  input  [63:0] io_ins_389, // @[:@39794.4]
  input  [63:0] io_ins_390, // @[:@39794.4]
  input  [63:0] io_ins_391, // @[:@39794.4]
  input  [63:0] io_ins_392, // @[:@39794.4]
  input  [63:0] io_ins_393, // @[:@39794.4]
  input  [63:0] io_ins_394, // @[:@39794.4]
  input  [63:0] io_ins_395, // @[:@39794.4]
  input  [63:0] io_ins_396, // @[:@39794.4]
  input  [63:0] io_ins_397, // @[:@39794.4]
  input  [63:0] io_ins_398, // @[:@39794.4]
  input  [63:0] io_ins_399, // @[:@39794.4]
  input  [63:0] io_ins_400, // @[:@39794.4]
  input  [63:0] io_ins_401, // @[:@39794.4]
  input  [63:0] io_ins_402, // @[:@39794.4]
  input  [63:0] io_ins_403, // @[:@39794.4]
  input  [63:0] io_ins_404, // @[:@39794.4]
  input  [63:0] io_ins_405, // @[:@39794.4]
  input  [63:0] io_ins_406, // @[:@39794.4]
  input  [63:0] io_ins_407, // @[:@39794.4]
  input  [63:0] io_ins_408, // @[:@39794.4]
  input  [63:0] io_ins_409, // @[:@39794.4]
  input  [63:0] io_ins_410, // @[:@39794.4]
  input  [63:0] io_ins_411, // @[:@39794.4]
  input  [63:0] io_ins_412, // @[:@39794.4]
  input  [63:0] io_ins_413, // @[:@39794.4]
  input  [63:0] io_ins_414, // @[:@39794.4]
  input  [63:0] io_ins_415, // @[:@39794.4]
  input  [63:0] io_ins_416, // @[:@39794.4]
  input  [63:0] io_ins_417, // @[:@39794.4]
  input  [63:0] io_ins_418, // @[:@39794.4]
  input  [63:0] io_ins_419, // @[:@39794.4]
  input  [63:0] io_ins_420, // @[:@39794.4]
  input  [63:0] io_ins_421, // @[:@39794.4]
  input  [63:0] io_ins_422, // @[:@39794.4]
  input  [63:0] io_ins_423, // @[:@39794.4]
  input  [63:0] io_ins_424, // @[:@39794.4]
  input  [63:0] io_ins_425, // @[:@39794.4]
  input  [63:0] io_ins_426, // @[:@39794.4]
  input  [63:0] io_ins_427, // @[:@39794.4]
  input  [63:0] io_ins_428, // @[:@39794.4]
  input  [63:0] io_ins_429, // @[:@39794.4]
  input  [63:0] io_ins_430, // @[:@39794.4]
  input  [63:0] io_ins_431, // @[:@39794.4]
  input  [63:0] io_ins_432, // @[:@39794.4]
  input  [63:0] io_ins_433, // @[:@39794.4]
  input  [63:0] io_ins_434, // @[:@39794.4]
  input  [63:0] io_ins_435, // @[:@39794.4]
  input  [63:0] io_ins_436, // @[:@39794.4]
  input  [63:0] io_ins_437, // @[:@39794.4]
  input  [63:0] io_ins_438, // @[:@39794.4]
  input  [63:0] io_ins_439, // @[:@39794.4]
  input  [63:0] io_ins_440, // @[:@39794.4]
  input  [63:0] io_ins_441, // @[:@39794.4]
  input  [63:0] io_ins_442, // @[:@39794.4]
  input  [63:0] io_ins_443, // @[:@39794.4]
  input  [63:0] io_ins_444, // @[:@39794.4]
  input  [63:0] io_ins_445, // @[:@39794.4]
  input  [63:0] io_ins_446, // @[:@39794.4]
  input  [63:0] io_ins_447, // @[:@39794.4]
  input  [63:0] io_ins_448, // @[:@39794.4]
  input  [63:0] io_ins_449, // @[:@39794.4]
  input  [63:0] io_ins_450, // @[:@39794.4]
  input  [63:0] io_ins_451, // @[:@39794.4]
  input  [63:0] io_ins_452, // @[:@39794.4]
  input  [63:0] io_ins_453, // @[:@39794.4]
  input  [63:0] io_ins_454, // @[:@39794.4]
  input  [63:0] io_ins_455, // @[:@39794.4]
  input  [63:0] io_ins_456, // @[:@39794.4]
  input  [63:0] io_ins_457, // @[:@39794.4]
  input  [63:0] io_ins_458, // @[:@39794.4]
  input  [63:0] io_ins_459, // @[:@39794.4]
  input  [63:0] io_ins_460, // @[:@39794.4]
  input  [63:0] io_ins_461, // @[:@39794.4]
  input  [63:0] io_ins_462, // @[:@39794.4]
  input  [63:0] io_ins_463, // @[:@39794.4]
  input  [63:0] io_ins_464, // @[:@39794.4]
  input  [63:0] io_ins_465, // @[:@39794.4]
  input  [63:0] io_ins_466, // @[:@39794.4]
  input  [63:0] io_ins_467, // @[:@39794.4]
  input  [63:0] io_ins_468, // @[:@39794.4]
  input  [63:0] io_ins_469, // @[:@39794.4]
  input  [63:0] io_ins_470, // @[:@39794.4]
  input  [63:0] io_ins_471, // @[:@39794.4]
  input  [63:0] io_ins_472, // @[:@39794.4]
  input  [63:0] io_ins_473, // @[:@39794.4]
  input  [63:0] io_ins_474, // @[:@39794.4]
  input  [63:0] io_ins_475, // @[:@39794.4]
  input  [63:0] io_ins_476, // @[:@39794.4]
  input  [63:0] io_ins_477, // @[:@39794.4]
  input  [63:0] io_ins_478, // @[:@39794.4]
  input  [63:0] io_ins_479, // @[:@39794.4]
  input  [63:0] io_ins_480, // @[:@39794.4]
  input  [63:0] io_ins_481, // @[:@39794.4]
  input  [63:0] io_ins_482, // @[:@39794.4]
  input  [63:0] io_ins_483, // @[:@39794.4]
  input  [63:0] io_ins_484, // @[:@39794.4]
  input  [63:0] io_ins_485, // @[:@39794.4]
  input  [63:0] io_ins_486, // @[:@39794.4]
  input  [63:0] io_ins_487, // @[:@39794.4]
  input  [63:0] io_ins_488, // @[:@39794.4]
  input  [63:0] io_ins_489, // @[:@39794.4]
  input  [63:0] io_ins_490, // @[:@39794.4]
  input  [63:0] io_ins_491, // @[:@39794.4]
  input  [63:0] io_ins_492, // @[:@39794.4]
  input  [63:0] io_ins_493, // @[:@39794.4]
  input  [63:0] io_ins_494, // @[:@39794.4]
  input  [63:0] io_ins_495, // @[:@39794.4]
  input  [63:0] io_ins_496, // @[:@39794.4]
  input  [63:0] io_ins_497, // @[:@39794.4]
  input  [63:0] io_ins_498, // @[:@39794.4]
  input  [63:0] io_ins_499, // @[:@39794.4]
  input  [63:0] io_ins_500, // @[:@39794.4]
  input  [63:0] io_ins_501, // @[:@39794.4]
  input  [63:0] io_ins_502, // @[:@39794.4]
  input  [63:0] io_ins_503, // @[:@39794.4]
  input  [63:0] io_ins_504, // @[:@39794.4]
  input  [63:0] io_ins_505, // @[:@39794.4]
  input  [63:0] io_ins_506, // @[:@39794.4]
  input  [63:0] io_ins_507, // @[:@39794.4]
  input  [63:0] io_ins_508, // @[:@39794.4]
  input  [63:0] io_ins_509, // @[:@39794.4]
  input  [63:0] io_ins_510, // @[:@39794.4]
  input  [63:0] io_ins_511, // @[:@39794.4]
  input  [63:0] io_ins_512, // @[:@39794.4]
  input  [63:0] io_ins_513, // @[:@39794.4]
  input  [63:0] io_ins_514, // @[:@39794.4]
  input  [63:0] io_ins_515, // @[:@39794.4]
  input  [63:0] io_ins_516, // @[:@39794.4]
  input  [63:0] io_ins_517, // @[:@39794.4]
  input  [63:0] io_ins_518, // @[:@39794.4]
  input  [63:0] io_ins_519, // @[:@39794.4]
  input  [63:0] io_ins_520, // @[:@39794.4]
  input  [63:0] io_ins_521, // @[:@39794.4]
  input  [9:0]  io_sel, // @[:@39794.4]
  output [63:0] io_out // @[:@39794.4]
);
  wire [63:0] _GEN_1; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_2; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_3; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_4; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_5; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_6; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_7; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_8; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_9; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_10; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_11; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_12; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_13; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_14; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_15; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_16; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_17; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_18; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_19; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_20; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_21; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_22; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_23; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_24; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_25; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_26; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_27; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_28; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_29; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_30; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_31; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_32; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_33; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_34; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_35; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_36; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_37; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_38; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_39; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_40; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_41; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_42; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_43; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_44; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_45; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_46; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_47; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_48; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_49; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_50; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_51; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_52; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_53; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_54; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_55; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_56; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_57; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_58; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_59; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_60; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_61; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_62; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_63; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_64; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_65; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_66; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_67; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_68; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_69; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_70; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_71; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_72; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_73; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_74; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_75; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_76; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_77; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_78; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_79; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_80; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_81; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_82; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_83; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_84; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_85; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_86; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_87; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_88; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_89; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_90; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_91; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_92; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_93; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_94; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_95; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_96; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_97; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_98; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_99; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_100; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_101; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_102; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_103; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_104; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_105; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_106; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_107; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_108; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_109; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_110; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_111; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_112; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_113; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_114; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_115; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_116; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_117; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_118; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_119; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_120; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_121; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_122; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_123; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_124; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_125; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_126; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_127; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_128; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_129; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_130; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_131; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_132; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_133; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_134; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_135; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_136; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_137; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_138; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_139; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_140; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_141; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_142; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_143; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_144; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_145; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_146; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_147; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_148; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_149; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_150; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_151; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_152; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_153; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_154; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_155; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_156; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_157; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_158; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_159; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_160; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_161; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_162; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_163; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_164; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_165; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_166; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_167; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_168; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_169; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_170; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_171; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_172; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_173; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_174; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_175; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_176; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_177; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_178; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_179; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_180; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_181; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_182; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_183; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_184; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_185; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_186; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_187; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_188; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_189; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_190; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_191; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_192; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_193; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_194; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_195; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_196; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_197; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_198; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_199; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_200; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_201; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_202; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_203; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_204; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_205; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_206; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_207; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_208; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_209; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_210; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_211; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_212; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_213; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_214; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_215; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_216; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_217; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_218; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_219; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_220; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_221; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_222; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_223; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_224; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_225; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_226; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_227; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_228; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_229; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_230; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_231; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_232; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_233; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_234; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_235; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_236; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_237; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_238; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_239; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_240; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_241; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_242; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_243; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_244; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_245; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_246; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_247; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_248; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_249; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_250; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_251; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_252; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_253; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_254; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_255; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_256; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_257; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_258; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_259; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_260; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_261; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_262; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_263; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_264; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_265; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_266; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_267; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_268; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_269; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_270; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_271; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_272; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_273; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_274; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_275; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_276; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_277; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_278; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_279; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_280; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_281; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_282; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_283; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_284; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_285; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_286; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_287; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_288; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_289; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_290; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_291; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_292; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_293; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_294; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_295; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_296; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_297; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_298; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_299; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_300; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_301; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_302; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_303; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_304; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_305; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_306; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_307; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_308; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_309; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_310; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_311; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_312; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_313; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_314; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_315; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_316; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_317; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_318; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_319; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_320; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_321; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_322; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_323; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_324; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_325; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_326; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_327; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_328; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_329; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_330; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_331; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_332; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_333; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_334; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_335; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_336; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_337; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_338; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_339; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_340; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_341; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_342; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_343; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_344; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_345; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_346; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_347; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_348; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_349; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_350; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_351; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_352; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_353; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_354; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_355; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_356; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_357; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_358; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_359; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_360; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_361; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_362; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_363; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_364; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_365; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_366; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_367; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_368; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_369; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_370; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_371; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_372; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_373; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_374; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_375; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_376; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_377; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_378; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_379; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_380; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_381; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_382; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_383; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_384; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_385; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_386; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_387; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_388; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_389; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_390; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_391; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_392; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_393; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_394; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_395; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_396; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_397; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_398; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_399; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_400; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_401; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_402; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_403; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_404; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_405; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_406; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_407; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_408; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_409; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_410; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_411; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_412; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_413; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_414; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_415; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_416; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_417; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_418; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_419; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_420; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_421; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_422; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_423; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_424; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_425; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_426; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_427; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_428; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_429; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_430; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_431; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_432; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_433; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_434; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_435; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_436; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_437; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_438; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_439; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_440; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_441; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_442; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_443; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_444; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_445; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_446; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_447; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_448; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_449; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_450; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_451; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_452; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_453; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_454; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_455; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_456; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_457; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_458; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_459; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_460; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_461; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_462; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_463; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_464; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_465; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_466; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_467; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_468; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_469; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_470; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_471; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_472; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_473; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_474; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_475; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_476; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_477; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_478; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_479; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_480; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_481; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_482; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_483; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_484; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_485; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_486; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_487; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_488; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_489; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_490; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_491; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_492; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_493; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_494; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_495; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_496; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_497; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_498; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_499; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_500; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_501; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_502; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_503; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_504; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_505; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_506; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_507; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_508; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_509; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_510; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_511; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_512; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_513; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_514; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_515; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_516; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_517; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_518; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_519; // @[MuxN.scala 16:10:@39796.4]
  wire [63:0] _GEN_520; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_1 = 10'h1 == io_sel ? io_ins_1 : io_ins_0; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_2 = 10'h2 == io_sel ? io_ins_2 : _GEN_1; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_3 = 10'h3 == io_sel ? io_ins_3 : _GEN_2; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_4 = 10'h4 == io_sel ? io_ins_4 : _GEN_3; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_5 = 10'h5 == io_sel ? io_ins_5 : _GEN_4; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_6 = 10'h6 == io_sel ? io_ins_6 : _GEN_5; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_7 = 10'h7 == io_sel ? io_ins_7 : _GEN_6; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_8 = 10'h8 == io_sel ? io_ins_8 : _GEN_7; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_9 = 10'h9 == io_sel ? io_ins_9 : _GEN_8; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_10 = 10'ha == io_sel ? io_ins_10 : _GEN_9; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_11 = 10'hb == io_sel ? io_ins_11 : _GEN_10; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_12 = 10'hc == io_sel ? io_ins_12 : _GEN_11; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_13 = 10'hd == io_sel ? io_ins_13 : _GEN_12; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_14 = 10'he == io_sel ? io_ins_14 : _GEN_13; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_15 = 10'hf == io_sel ? io_ins_15 : _GEN_14; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_16 = 10'h10 == io_sel ? io_ins_16 : _GEN_15; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_17 = 10'h11 == io_sel ? io_ins_17 : _GEN_16; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_18 = 10'h12 == io_sel ? io_ins_18 : _GEN_17; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_19 = 10'h13 == io_sel ? io_ins_19 : _GEN_18; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_20 = 10'h14 == io_sel ? io_ins_20 : _GEN_19; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_21 = 10'h15 == io_sel ? io_ins_21 : _GEN_20; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_22 = 10'h16 == io_sel ? io_ins_22 : _GEN_21; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_23 = 10'h17 == io_sel ? io_ins_23 : _GEN_22; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_24 = 10'h18 == io_sel ? io_ins_24 : _GEN_23; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_25 = 10'h19 == io_sel ? io_ins_25 : _GEN_24; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_26 = 10'h1a == io_sel ? io_ins_26 : _GEN_25; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_27 = 10'h1b == io_sel ? io_ins_27 : _GEN_26; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_28 = 10'h1c == io_sel ? io_ins_28 : _GEN_27; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_29 = 10'h1d == io_sel ? io_ins_29 : _GEN_28; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_30 = 10'h1e == io_sel ? io_ins_30 : _GEN_29; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_31 = 10'h1f == io_sel ? io_ins_31 : _GEN_30; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_32 = 10'h20 == io_sel ? io_ins_32 : _GEN_31; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_33 = 10'h21 == io_sel ? io_ins_33 : _GEN_32; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_34 = 10'h22 == io_sel ? io_ins_34 : _GEN_33; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_35 = 10'h23 == io_sel ? io_ins_35 : _GEN_34; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_36 = 10'h24 == io_sel ? io_ins_36 : _GEN_35; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_37 = 10'h25 == io_sel ? io_ins_37 : _GEN_36; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_38 = 10'h26 == io_sel ? io_ins_38 : _GEN_37; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_39 = 10'h27 == io_sel ? io_ins_39 : _GEN_38; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_40 = 10'h28 == io_sel ? io_ins_40 : _GEN_39; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_41 = 10'h29 == io_sel ? io_ins_41 : _GEN_40; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_42 = 10'h2a == io_sel ? io_ins_42 : _GEN_41; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_43 = 10'h2b == io_sel ? io_ins_43 : _GEN_42; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_44 = 10'h2c == io_sel ? io_ins_44 : _GEN_43; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_45 = 10'h2d == io_sel ? io_ins_45 : _GEN_44; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_46 = 10'h2e == io_sel ? io_ins_46 : _GEN_45; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_47 = 10'h2f == io_sel ? io_ins_47 : _GEN_46; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_48 = 10'h30 == io_sel ? io_ins_48 : _GEN_47; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_49 = 10'h31 == io_sel ? io_ins_49 : _GEN_48; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_50 = 10'h32 == io_sel ? io_ins_50 : _GEN_49; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_51 = 10'h33 == io_sel ? io_ins_51 : _GEN_50; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_52 = 10'h34 == io_sel ? io_ins_52 : _GEN_51; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_53 = 10'h35 == io_sel ? io_ins_53 : _GEN_52; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_54 = 10'h36 == io_sel ? io_ins_54 : _GEN_53; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_55 = 10'h37 == io_sel ? io_ins_55 : _GEN_54; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_56 = 10'h38 == io_sel ? io_ins_56 : _GEN_55; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_57 = 10'h39 == io_sel ? io_ins_57 : _GEN_56; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_58 = 10'h3a == io_sel ? io_ins_58 : _GEN_57; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_59 = 10'h3b == io_sel ? io_ins_59 : _GEN_58; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_60 = 10'h3c == io_sel ? io_ins_60 : _GEN_59; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_61 = 10'h3d == io_sel ? io_ins_61 : _GEN_60; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_62 = 10'h3e == io_sel ? io_ins_62 : _GEN_61; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_63 = 10'h3f == io_sel ? io_ins_63 : _GEN_62; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_64 = 10'h40 == io_sel ? io_ins_64 : _GEN_63; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_65 = 10'h41 == io_sel ? io_ins_65 : _GEN_64; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_66 = 10'h42 == io_sel ? io_ins_66 : _GEN_65; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_67 = 10'h43 == io_sel ? io_ins_67 : _GEN_66; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_68 = 10'h44 == io_sel ? io_ins_68 : _GEN_67; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_69 = 10'h45 == io_sel ? io_ins_69 : _GEN_68; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_70 = 10'h46 == io_sel ? io_ins_70 : _GEN_69; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_71 = 10'h47 == io_sel ? io_ins_71 : _GEN_70; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_72 = 10'h48 == io_sel ? io_ins_72 : _GEN_71; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_73 = 10'h49 == io_sel ? io_ins_73 : _GEN_72; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_74 = 10'h4a == io_sel ? io_ins_74 : _GEN_73; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_75 = 10'h4b == io_sel ? io_ins_75 : _GEN_74; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_76 = 10'h4c == io_sel ? io_ins_76 : _GEN_75; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_77 = 10'h4d == io_sel ? io_ins_77 : _GEN_76; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_78 = 10'h4e == io_sel ? io_ins_78 : _GEN_77; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_79 = 10'h4f == io_sel ? io_ins_79 : _GEN_78; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_80 = 10'h50 == io_sel ? io_ins_80 : _GEN_79; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_81 = 10'h51 == io_sel ? io_ins_81 : _GEN_80; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_82 = 10'h52 == io_sel ? io_ins_82 : _GEN_81; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_83 = 10'h53 == io_sel ? io_ins_83 : _GEN_82; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_84 = 10'h54 == io_sel ? io_ins_84 : _GEN_83; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_85 = 10'h55 == io_sel ? io_ins_85 : _GEN_84; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_86 = 10'h56 == io_sel ? io_ins_86 : _GEN_85; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_87 = 10'h57 == io_sel ? io_ins_87 : _GEN_86; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_88 = 10'h58 == io_sel ? io_ins_88 : _GEN_87; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_89 = 10'h59 == io_sel ? io_ins_89 : _GEN_88; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_90 = 10'h5a == io_sel ? io_ins_90 : _GEN_89; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_91 = 10'h5b == io_sel ? io_ins_91 : _GEN_90; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_92 = 10'h5c == io_sel ? io_ins_92 : _GEN_91; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_93 = 10'h5d == io_sel ? io_ins_93 : _GEN_92; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_94 = 10'h5e == io_sel ? io_ins_94 : _GEN_93; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_95 = 10'h5f == io_sel ? io_ins_95 : _GEN_94; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_96 = 10'h60 == io_sel ? io_ins_96 : _GEN_95; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_97 = 10'h61 == io_sel ? io_ins_97 : _GEN_96; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_98 = 10'h62 == io_sel ? io_ins_98 : _GEN_97; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_99 = 10'h63 == io_sel ? io_ins_99 : _GEN_98; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_100 = 10'h64 == io_sel ? io_ins_100 : _GEN_99; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_101 = 10'h65 == io_sel ? io_ins_101 : _GEN_100; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_102 = 10'h66 == io_sel ? io_ins_102 : _GEN_101; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_103 = 10'h67 == io_sel ? io_ins_103 : _GEN_102; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_104 = 10'h68 == io_sel ? io_ins_104 : _GEN_103; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_105 = 10'h69 == io_sel ? io_ins_105 : _GEN_104; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_106 = 10'h6a == io_sel ? io_ins_106 : _GEN_105; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_107 = 10'h6b == io_sel ? io_ins_107 : _GEN_106; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_108 = 10'h6c == io_sel ? io_ins_108 : _GEN_107; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_109 = 10'h6d == io_sel ? io_ins_109 : _GEN_108; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_110 = 10'h6e == io_sel ? io_ins_110 : _GEN_109; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_111 = 10'h6f == io_sel ? io_ins_111 : _GEN_110; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_112 = 10'h70 == io_sel ? io_ins_112 : _GEN_111; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_113 = 10'h71 == io_sel ? io_ins_113 : _GEN_112; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_114 = 10'h72 == io_sel ? io_ins_114 : _GEN_113; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_115 = 10'h73 == io_sel ? io_ins_115 : _GEN_114; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_116 = 10'h74 == io_sel ? io_ins_116 : _GEN_115; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_117 = 10'h75 == io_sel ? io_ins_117 : _GEN_116; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_118 = 10'h76 == io_sel ? io_ins_118 : _GEN_117; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_119 = 10'h77 == io_sel ? io_ins_119 : _GEN_118; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_120 = 10'h78 == io_sel ? io_ins_120 : _GEN_119; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_121 = 10'h79 == io_sel ? io_ins_121 : _GEN_120; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_122 = 10'h7a == io_sel ? io_ins_122 : _GEN_121; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_123 = 10'h7b == io_sel ? io_ins_123 : _GEN_122; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_124 = 10'h7c == io_sel ? io_ins_124 : _GEN_123; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_125 = 10'h7d == io_sel ? io_ins_125 : _GEN_124; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_126 = 10'h7e == io_sel ? io_ins_126 : _GEN_125; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_127 = 10'h7f == io_sel ? io_ins_127 : _GEN_126; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_128 = 10'h80 == io_sel ? io_ins_128 : _GEN_127; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_129 = 10'h81 == io_sel ? io_ins_129 : _GEN_128; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_130 = 10'h82 == io_sel ? io_ins_130 : _GEN_129; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_131 = 10'h83 == io_sel ? io_ins_131 : _GEN_130; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_132 = 10'h84 == io_sel ? io_ins_132 : _GEN_131; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_133 = 10'h85 == io_sel ? io_ins_133 : _GEN_132; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_134 = 10'h86 == io_sel ? io_ins_134 : _GEN_133; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_135 = 10'h87 == io_sel ? io_ins_135 : _GEN_134; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_136 = 10'h88 == io_sel ? io_ins_136 : _GEN_135; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_137 = 10'h89 == io_sel ? io_ins_137 : _GEN_136; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_138 = 10'h8a == io_sel ? io_ins_138 : _GEN_137; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_139 = 10'h8b == io_sel ? io_ins_139 : _GEN_138; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_140 = 10'h8c == io_sel ? io_ins_140 : _GEN_139; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_141 = 10'h8d == io_sel ? io_ins_141 : _GEN_140; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_142 = 10'h8e == io_sel ? io_ins_142 : _GEN_141; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_143 = 10'h8f == io_sel ? io_ins_143 : _GEN_142; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_144 = 10'h90 == io_sel ? io_ins_144 : _GEN_143; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_145 = 10'h91 == io_sel ? io_ins_145 : _GEN_144; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_146 = 10'h92 == io_sel ? io_ins_146 : _GEN_145; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_147 = 10'h93 == io_sel ? io_ins_147 : _GEN_146; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_148 = 10'h94 == io_sel ? io_ins_148 : _GEN_147; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_149 = 10'h95 == io_sel ? io_ins_149 : _GEN_148; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_150 = 10'h96 == io_sel ? io_ins_150 : _GEN_149; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_151 = 10'h97 == io_sel ? io_ins_151 : _GEN_150; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_152 = 10'h98 == io_sel ? io_ins_152 : _GEN_151; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_153 = 10'h99 == io_sel ? io_ins_153 : _GEN_152; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_154 = 10'h9a == io_sel ? io_ins_154 : _GEN_153; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_155 = 10'h9b == io_sel ? io_ins_155 : _GEN_154; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_156 = 10'h9c == io_sel ? io_ins_156 : _GEN_155; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_157 = 10'h9d == io_sel ? io_ins_157 : _GEN_156; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_158 = 10'h9e == io_sel ? io_ins_158 : _GEN_157; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_159 = 10'h9f == io_sel ? io_ins_159 : _GEN_158; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_160 = 10'ha0 == io_sel ? io_ins_160 : _GEN_159; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_161 = 10'ha1 == io_sel ? io_ins_161 : _GEN_160; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_162 = 10'ha2 == io_sel ? io_ins_162 : _GEN_161; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_163 = 10'ha3 == io_sel ? io_ins_163 : _GEN_162; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_164 = 10'ha4 == io_sel ? io_ins_164 : _GEN_163; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_165 = 10'ha5 == io_sel ? io_ins_165 : _GEN_164; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_166 = 10'ha6 == io_sel ? io_ins_166 : _GEN_165; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_167 = 10'ha7 == io_sel ? io_ins_167 : _GEN_166; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_168 = 10'ha8 == io_sel ? io_ins_168 : _GEN_167; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_169 = 10'ha9 == io_sel ? io_ins_169 : _GEN_168; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_170 = 10'haa == io_sel ? io_ins_170 : _GEN_169; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_171 = 10'hab == io_sel ? io_ins_171 : _GEN_170; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_172 = 10'hac == io_sel ? io_ins_172 : _GEN_171; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_173 = 10'had == io_sel ? io_ins_173 : _GEN_172; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_174 = 10'hae == io_sel ? io_ins_174 : _GEN_173; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_175 = 10'haf == io_sel ? io_ins_175 : _GEN_174; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_176 = 10'hb0 == io_sel ? io_ins_176 : _GEN_175; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_177 = 10'hb1 == io_sel ? io_ins_177 : _GEN_176; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_178 = 10'hb2 == io_sel ? io_ins_178 : _GEN_177; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_179 = 10'hb3 == io_sel ? io_ins_179 : _GEN_178; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_180 = 10'hb4 == io_sel ? io_ins_180 : _GEN_179; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_181 = 10'hb5 == io_sel ? io_ins_181 : _GEN_180; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_182 = 10'hb6 == io_sel ? io_ins_182 : _GEN_181; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_183 = 10'hb7 == io_sel ? io_ins_183 : _GEN_182; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_184 = 10'hb8 == io_sel ? io_ins_184 : _GEN_183; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_185 = 10'hb9 == io_sel ? io_ins_185 : _GEN_184; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_186 = 10'hba == io_sel ? io_ins_186 : _GEN_185; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_187 = 10'hbb == io_sel ? io_ins_187 : _GEN_186; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_188 = 10'hbc == io_sel ? io_ins_188 : _GEN_187; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_189 = 10'hbd == io_sel ? io_ins_189 : _GEN_188; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_190 = 10'hbe == io_sel ? io_ins_190 : _GEN_189; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_191 = 10'hbf == io_sel ? io_ins_191 : _GEN_190; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_192 = 10'hc0 == io_sel ? io_ins_192 : _GEN_191; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_193 = 10'hc1 == io_sel ? io_ins_193 : _GEN_192; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_194 = 10'hc2 == io_sel ? io_ins_194 : _GEN_193; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_195 = 10'hc3 == io_sel ? io_ins_195 : _GEN_194; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_196 = 10'hc4 == io_sel ? io_ins_196 : _GEN_195; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_197 = 10'hc5 == io_sel ? io_ins_197 : _GEN_196; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_198 = 10'hc6 == io_sel ? io_ins_198 : _GEN_197; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_199 = 10'hc7 == io_sel ? io_ins_199 : _GEN_198; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_200 = 10'hc8 == io_sel ? io_ins_200 : _GEN_199; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_201 = 10'hc9 == io_sel ? io_ins_201 : _GEN_200; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_202 = 10'hca == io_sel ? io_ins_202 : _GEN_201; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_203 = 10'hcb == io_sel ? io_ins_203 : _GEN_202; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_204 = 10'hcc == io_sel ? io_ins_204 : _GEN_203; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_205 = 10'hcd == io_sel ? io_ins_205 : _GEN_204; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_206 = 10'hce == io_sel ? io_ins_206 : _GEN_205; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_207 = 10'hcf == io_sel ? io_ins_207 : _GEN_206; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_208 = 10'hd0 == io_sel ? io_ins_208 : _GEN_207; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_209 = 10'hd1 == io_sel ? io_ins_209 : _GEN_208; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_210 = 10'hd2 == io_sel ? io_ins_210 : _GEN_209; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_211 = 10'hd3 == io_sel ? io_ins_211 : _GEN_210; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_212 = 10'hd4 == io_sel ? io_ins_212 : _GEN_211; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_213 = 10'hd5 == io_sel ? io_ins_213 : _GEN_212; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_214 = 10'hd6 == io_sel ? io_ins_214 : _GEN_213; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_215 = 10'hd7 == io_sel ? io_ins_215 : _GEN_214; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_216 = 10'hd8 == io_sel ? io_ins_216 : _GEN_215; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_217 = 10'hd9 == io_sel ? io_ins_217 : _GEN_216; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_218 = 10'hda == io_sel ? io_ins_218 : _GEN_217; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_219 = 10'hdb == io_sel ? io_ins_219 : _GEN_218; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_220 = 10'hdc == io_sel ? io_ins_220 : _GEN_219; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_221 = 10'hdd == io_sel ? io_ins_221 : _GEN_220; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_222 = 10'hde == io_sel ? io_ins_222 : _GEN_221; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_223 = 10'hdf == io_sel ? io_ins_223 : _GEN_222; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_224 = 10'he0 == io_sel ? io_ins_224 : _GEN_223; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_225 = 10'he1 == io_sel ? io_ins_225 : _GEN_224; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_226 = 10'he2 == io_sel ? io_ins_226 : _GEN_225; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_227 = 10'he3 == io_sel ? io_ins_227 : _GEN_226; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_228 = 10'he4 == io_sel ? io_ins_228 : _GEN_227; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_229 = 10'he5 == io_sel ? io_ins_229 : _GEN_228; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_230 = 10'he6 == io_sel ? io_ins_230 : _GEN_229; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_231 = 10'he7 == io_sel ? io_ins_231 : _GEN_230; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_232 = 10'he8 == io_sel ? io_ins_232 : _GEN_231; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_233 = 10'he9 == io_sel ? io_ins_233 : _GEN_232; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_234 = 10'hea == io_sel ? io_ins_234 : _GEN_233; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_235 = 10'heb == io_sel ? io_ins_235 : _GEN_234; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_236 = 10'hec == io_sel ? io_ins_236 : _GEN_235; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_237 = 10'hed == io_sel ? io_ins_237 : _GEN_236; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_238 = 10'hee == io_sel ? io_ins_238 : _GEN_237; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_239 = 10'hef == io_sel ? io_ins_239 : _GEN_238; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_240 = 10'hf0 == io_sel ? io_ins_240 : _GEN_239; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_241 = 10'hf1 == io_sel ? io_ins_241 : _GEN_240; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_242 = 10'hf2 == io_sel ? io_ins_242 : _GEN_241; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_243 = 10'hf3 == io_sel ? io_ins_243 : _GEN_242; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_244 = 10'hf4 == io_sel ? io_ins_244 : _GEN_243; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_245 = 10'hf5 == io_sel ? io_ins_245 : _GEN_244; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_246 = 10'hf6 == io_sel ? io_ins_246 : _GEN_245; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_247 = 10'hf7 == io_sel ? io_ins_247 : _GEN_246; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_248 = 10'hf8 == io_sel ? io_ins_248 : _GEN_247; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_249 = 10'hf9 == io_sel ? io_ins_249 : _GEN_248; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_250 = 10'hfa == io_sel ? io_ins_250 : _GEN_249; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_251 = 10'hfb == io_sel ? io_ins_251 : _GEN_250; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_252 = 10'hfc == io_sel ? io_ins_252 : _GEN_251; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_253 = 10'hfd == io_sel ? io_ins_253 : _GEN_252; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_254 = 10'hfe == io_sel ? io_ins_254 : _GEN_253; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_255 = 10'hff == io_sel ? io_ins_255 : _GEN_254; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_256 = 10'h100 == io_sel ? io_ins_256 : _GEN_255; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_257 = 10'h101 == io_sel ? io_ins_257 : _GEN_256; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_258 = 10'h102 == io_sel ? io_ins_258 : _GEN_257; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_259 = 10'h103 == io_sel ? io_ins_259 : _GEN_258; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_260 = 10'h104 == io_sel ? io_ins_260 : _GEN_259; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_261 = 10'h105 == io_sel ? io_ins_261 : _GEN_260; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_262 = 10'h106 == io_sel ? io_ins_262 : _GEN_261; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_263 = 10'h107 == io_sel ? io_ins_263 : _GEN_262; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_264 = 10'h108 == io_sel ? io_ins_264 : _GEN_263; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_265 = 10'h109 == io_sel ? io_ins_265 : _GEN_264; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_266 = 10'h10a == io_sel ? io_ins_266 : _GEN_265; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_267 = 10'h10b == io_sel ? io_ins_267 : _GEN_266; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_268 = 10'h10c == io_sel ? io_ins_268 : _GEN_267; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_269 = 10'h10d == io_sel ? io_ins_269 : _GEN_268; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_270 = 10'h10e == io_sel ? io_ins_270 : _GEN_269; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_271 = 10'h10f == io_sel ? io_ins_271 : _GEN_270; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_272 = 10'h110 == io_sel ? io_ins_272 : _GEN_271; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_273 = 10'h111 == io_sel ? io_ins_273 : _GEN_272; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_274 = 10'h112 == io_sel ? io_ins_274 : _GEN_273; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_275 = 10'h113 == io_sel ? io_ins_275 : _GEN_274; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_276 = 10'h114 == io_sel ? io_ins_276 : _GEN_275; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_277 = 10'h115 == io_sel ? io_ins_277 : _GEN_276; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_278 = 10'h116 == io_sel ? io_ins_278 : _GEN_277; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_279 = 10'h117 == io_sel ? io_ins_279 : _GEN_278; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_280 = 10'h118 == io_sel ? io_ins_280 : _GEN_279; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_281 = 10'h119 == io_sel ? io_ins_281 : _GEN_280; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_282 = 10'h11a == io_sel ? io_ins_282 : _GEN_281; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_283 = 10'h11b == io_sel ? io_ins_283 : _GEN_282; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_284 = 10'h11c == io_sel ? io_ins_284 : _GEN_283; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_285 = 10'h11d == io_sel ? io_ins_285 : _GEN_284; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_286 = 10'h11e == io_sel ? io_ins_286 : _GEN_285; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_287 = 10'h11f == io_sel ? io_ins_287 : _GEN_286; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_288 = 10'h120 == io_sel ? io_ins_288 : _GEN_287; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_289 = 10'h121 == io_sel ? io_ins_289 : _GEN_288; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_290 = 10'h122 == io_sel ? io_ins_290 : _GEN_289; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_291 = 10'h123 == io_sel ? io_ins_291 : _GEN_290; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_292 = 10'h124 == io_sel ? io_ins_292 : _GEN_291; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_293 = 10'h125 == io_sel ? io_ins_293 : _GEN_292; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_294 = 10'h126 == io_sel ? io_ins_294 : _GEN_293; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_295 = 10'h127 == io_sel ? io_ins_295 : _GEN_294; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_296 = 10'h128 == io_sel ? io_ins_296 : _GEN_295; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_297 = 10'h129 == io_sel ? io_ins_297 : _GEN_296; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_298 = 10'h12a == io_sel ? io_ins_298 : _GEN_297; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_299 = 10'h12b == io_sel ? io_ins_299 : _GEN_298; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_300 = 10'h12c == io_sel ? io_ins_300 : _GEN_299; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_301 = 10'h12d == io_sel ? io_ins_301 : _GEN_300; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_302 = 10'h12e == io_sel ? io_ins_302 : _GEN_301; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_303 = 10'h12f == io_sel ? io_ins_303 : _GEN_302; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_304 = 10'h130 == io_sel ? io_ins_304 : _GEN_303; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_305 = 10'h131 == io_sel ? io_ins_305 : _GEN_304; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_306 = 10'h132 == io_sel ? io_ins_306 : _GEN_305; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_307 = 10'h133 == io_sel ? io_ins_307 : _GEN_306; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_308 = 10'h134 == io_sel ? io_ins_308 : _GEN_307; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_309 = 10'h135 == io_sel ? io_ins_309 : _GEN_308; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_310 = 10'h136 == io_sel ? io_ins_310 : _GEN_309; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_311 = 10'h137 == io_sel ? io_ins_311 : _GEN_310; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_312 = 10'h138 == io_sel ? io_ins_312 : _GEN_311; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_313 = 10'h139 == io_sel ? io_ins_313 : _GEN_312; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_314 = 10'h13a == io_sel ? io_ins_314 : _GEN_313; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_315 = 10'h13b == io_sel ? io_ins_315 : _GEN_314; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_316 = 10'h13c == io_sel ? io_ins_316 : _GEN_315; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_317 = 10'h13d == io_sel ? io_ins_317 : _GEN_316; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_318 = 10'h13e == io_sel ? io_ins_318 : _GEN_317; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_319 = 10'h13f == io_sel ? io_ins_319 : _GEN_318; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_320 = 10'h140 == io_sel ? io_ins_320 : _GEN_319; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_321 = 10'h141 == io_sel ? io_ins_321 : _GEN_320; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_322 = 10'h142 == io_sel ? io_ins_322 : _GEN_321; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_323 = 10'h143 == io_sel ? io_ins_323 : _GEN_322; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_324 = 10'h144 == io_sel ? io_ins_324 : _GEN_323; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_325 = 10'h145 == io_sel ? io_ins_325 : _GEN_324; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_326 = 10'h146 == io_sel ? io_ins_326 : _GEN_325; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_327 = 10'h147 == io_sel ? io_ins_327 : _GEN_326; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_328 = 10'h148 == io_sel ? io_ins_328 : _GEN_327; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_329 = 10'h149 == io_sel ? io_ins_329 : _GEN_328; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_330 = 10'h14a == io_sel ? io_ins_330 : _GEN_329; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_331 = 10'h14b == io_sel ? io_ins_331 : _GEN_330; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_332 = 10'h14c == io_sel ? io_ins_332 : _GEN_331; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_333 = 10'h14d == io_sel ? io_ins_333 : _GEN_332; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_334 = 10'h14e == io_sel ? io_ins_334 : _GEN_333; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_335 = 10'h14f == io_sel ? io_ins_335 : _GEN_334; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_336 = 10'h150 == io_sel ? io_ins_336 : _GEN_335; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_337 = 10'h151 == io_sel ? io_ins_337 : _GEN_336; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_338 = 10'h152 == io_sel ? io_ins_338 : _GEN_337; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_339 = 10'h153 == io_sel ? io_ins_339 : _GEN_338; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_340 = 10'h154 == io_sel ? io_ins_340 : _GEN_339; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_341 = 10'h155 == io_sel ? io_ins_341 : _GEN_340; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_342 = 10'h156 == io_sel ? io_ins_342 : _GEN_341; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_343 = 10'h157 == io_sel ? io_ins_343 : _GEN_342; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_344 = 10'h158 == io_sel ? io_ins_344 : _GEN_343; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_345 = 10'h159 == io_sel ? io_ins_345 : _GEN_344; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_346 = 10'h15a == io_sel ? io_ins_346 : _GEN_345; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_347 = 10'h15b == io_sel ? io_ins_347 : _GEN_346; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_348 = 10'h15c == io_sel ? io_ins_348 : _GEN_347; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_349 = 10'h15d == io_sel ? io_ins_349 : _GEN_348; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_350 = 10'h15e == io_sel ? io_ins_350 : _GEN_349; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_351 = 10'h15f == io_sel ? io_ins_351 : _GEN_350; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_352 = 10'h160 == io_sel ? io_ins_352 : _GEN_351; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_353 = 10'h161 == io_sel ? io_ins_353 : _GEN_352; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_354 = 10'h162 == io_sel ? io_ins_354 : _GEN_353; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_355 = 10'h163 == io_sel ? io_ins_355 : _GEN_354; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_356 = 10'h164 == io_sel ? io_ins_356 : _GEN_355; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_357 = 10'h165 == io_sel ? io_ins_357 : _GEN_356; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_358 = 10'h166 == io_sel ? io_ins_358 : _GEN_357; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_359 = 10'h167 == io_sel ? io_ins_359 : _GEN_358; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_360 = 10'h168 == io_sel ? io_ins_360 : _GEN_359; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_361 = 10'h169 == io_sel ? io_ins_361 : _GEN_360; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_362 = 10'h16a == io_sel ? io_ins_362 : _GEN_361; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_363 = 10'h16b == io_sel ? io_ins_363 : _GEN_362; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_364 = 10'h16c == io_sel ? io_ins_364 : _GEN_363; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_365 = 10'h16d == io_sel ? io_ins_365 : _GEN_364; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_366 = 10'h16e == io_sel ? io_ins_366 : _GEN_365; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_367 = 10'h16f == io_sel ? io_ins_367 : _GEN_366; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_368 = 10'h170 == io_sel ? io_ins_368 : _GEN_367; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_369 = 10'h171 == io_sel ? io_ins_369 : _GEN_368; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_370 = 10'h172 == io_sel ? io_ins_370 : _GEN_369; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_371 = 10'h173 == io_sel ? io_ins_371 : _GEN_370; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_372 = 10'h174 == io_sel ? io_ins_372 : _GEN_371; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_373 = 10'h175 == io_sel ? io_ins_373 : _GEN_372; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_374 = 10'h176 == io_sel ? io_ins_374 : _GEN_373; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_375 = 10'h177 == io_sel ? io_ins_375 : _GEN_374; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_376 = 10'h178 == io_sel ? io_ins_376 : _GEN_375; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_377 = 10'h179 == io_sel ? io_ins_377 : _GEN_376; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_378 = 10'h17a == io_sel ? io_ins_378 : _GEN_377; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_379 = 10'h17b == io_sel ? io_ins_379 : _GEN_378; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_380 = 10'h17c == io_sel ? io_ins_380 : _GEN_379; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_381 = 10'h17d == io_sel ? io_ins_381 : _GEN_380; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_382 = 10'h17e == io_sel ? io_ins_382 : _GEN_381; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_383 = 10'h17f == io_sel ? io_ins_383 : _GEN_382; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_384 = 10'h180 == io_sel ? io_ins_384 : _GEN_383; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_385 = 10'h181 == io_sel ? io_ins_385 : _GEN_384; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_386 = 10'h182 == io_sel ? io_ins_386 : _GEN_385; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_387 = 10'h183 == io_sel ? io_ins_387 : _GEN_386; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_388 = 10'h184 == io_sel ? io_ins_388 : _GEN_387; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_389 = 10'h185 == io_sel ? io_ins_389 : _GEN_388; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_390 = 10'h186 == io_sel ? io_ins_390 : _GEN_389; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_391 = 10'h187 == io_sel ? io_ins_391 : _GEN_390; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_392 = 10'h188 == io_sel ? io_ins_392 : _GEN_391; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_393 = 10'h189 == io_sel ? io_ins_393 : _GEN_392; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_394 = 10'h18a == io_sel ? io_ins_394 : _GEN_393; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_395 = 10'h18b == io_sel ? io_ins_395 : _GEN_394; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_396 = 10'h18c == io_sel ? io_ins_396 : _GEN_395; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_397 = 10'h18d == io_sel ? io_ins_397 : _GEN_396; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_398 = 10'h18e == io_sel ? io_ins_398 : _GEN_397; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_399 = 10'h18f == io_sel ? io_ins_399 : _GEN_398; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_400 = 10'h190 == io_sel ? io_ins_400 : _GEN_399; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_401 = 10'h191 == io_sel ? io_ins_401 : _GEN_400; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_402 = 10'h192 == io_sel ? io_ins_402 : _GEN_401; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_403 = 10'h193 == io_sel ? io_ins_403 : _GEN_402; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_404 = 10'h194 == io_sel ? io_ins_404 : _GEN_403; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_405 = 10'h195 == io_sel ? io_ins_405 : _GEN_404; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_406 = 10'h196 == io_sel ? io_ins_406 : _GEN_405; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_407 = 10'h197 == io_sel ? io_ins_407 : _GEN_406; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_408 = 10'h198 == io_sel ? io_ins_408 : _GEN_407; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_409 = 10'h199 == io_sel ? io_ins_409 : _GEN_408; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_410 = 10'h19a == io_sel ? io_ins_410 : _GEN_409; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_411 = 10'h19b == io_sel ? io_ins_411 : _GEN_410; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_412 = 10'h19c == io_sel ? io_ins_412 : _GEN_411; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_413 = 10'h19d == io_sel ? io_ins_413 : _GEN_412; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_414 = 10'h19e == io_sel ? io_ins_414 : _GEN_413; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_415 = 10'h19f == io_sel ? io_ins_415 : _GEN_414; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_416 = 10'h1a0 == io_sel ? io_ins_416 : _GEN_415; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_417 = 10'h1a1 == io_sel ? io_ins_417 : _GEN_416; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_418 = 10'h1a2 == io_sel ? io_ins_418 : _GEN_417; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_419 = 10'h1a3 == io_sel ? io_ins_419 : _GEN_418; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_420 = 10'h1a4 == io_sel ? io_ins_420 : _GEN_419; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_421 = 10'h1a5 == io_sel ? io_ins_421 : _GEN_420; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_422 = 10'h1a6 == io_sel ? io_ins_422 : _GEN_421; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_423 = 10'h1a7 == io_sel ? io_ins_423 : _GEN_422; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_424 = 10'h1a8 == io_sel ? io_ins_424 : _GEN_423; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_425 = 10'h1a9 == io_sel ? io_ins_425 : _GEN_424; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_426 = 10'h1aa == io_sel ? io_ins_426 : _GEN_425; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_427 = 10'h1ab == io_sel ? io_ins_427 : _GEN_426; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_428 = 10'h1ac == io_sel ? io_ins_428 : _GEN_427; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_429 = 10'h1ad == io_sel ? io_ins_429 : _GEN_428; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_430 = 10'h1ae == io_sel ? io_ins_430 : _GEN_429; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_431 = 10'h1af == io_sel ? io_ins_431 : _GEN_430; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_432 = 10'h1b0 == io_sel ? io_ins_432 : _GEN_431; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_433 = 10'h1b1 == io_sel ? io_ins_433 : _GEN_432; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_434 = 10'h1b2 == io_sel ? io_ins_434 : _GEN_433; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_435 = 10'h1b3 == io_sel ? io_ins_435 : _GEN_434; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_436 = 10'h1b4 == io_sel ? io_ins_436 : _GEN_435; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_437 = 10'h1b5 == io_sel ? io_ins_437 : _GEN_436; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_438 = 10'h1b6 == io_sel ? io_ins_438 : _GEN_437; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_439 = 10'h1b7 == io_sel ? io_ins_439 : _GEN_438; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_440 = 10'h1b8 == io_sel ? io_ins_440 : _GEN_439; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_441 = 10'h1b9 == io_sel ? io_ins_441 : _GEN_440; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_442 = 10'h1ba == io_sel ? io_ins_442 : _GEN_441; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_443 = 10'h1bb == io_sel ? io_ins_443 : _GEN_442; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_444 = 10'h1bc == io_sel ? io_ins_444 : _GEN_443; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_445 = 10'h1bd == io_sel ? io_ins_445 : _GEN_444; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_446 = 10'h1be == io_sel ? io_ins_446 : _GEN_445; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_447 = 10'h1bf == io_sel ? io_ins_447 : _GEN_446; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_448 = 10'h1c0 == io_sel ? io_ins_448 : _GEN_447; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_449 = 10'h1c1 == io_sel ? io_ins_449 : _GEN_448; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_450 = 10'h1c2 == io_sel ? io_ins_450 : _GEN_449; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_451 = 10'h1c3 == io_sel ? io_ins_451 : _GEN_450; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_452 = 10'h1c4 == io_sel ? io_ins_452 : _GEN_451; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_453 = 10'h1c5 == io_sel ? io_ins_453 : _GEN_452; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_454 = 10'h1c6 == io_sel ? io_ins_454 : _GEN_453; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_455 = 10'h1c7 == io_sel ? io_ins_455 : _GEN_454; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_456 = 10'h1c8 == io_sel ? io_ins_456 : _GEN_455; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_457 = 10'h1c9 == io_sel ? io_ins_457 : _GEN_456; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_458 = 10'h1ca == io_sel ? io_ins_458 : _GEN_457; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_459 = 10'h1cb == io_sel ? io_ins_459 : _GEN_458; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_460 = 10'h1cc == io_sel ? io_ins_460 : _GEN_459; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_461 = 10'h1cd == io_sel ? io_ins_461 : _GEN_460; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_462 = 10'h1ce == io_sel ? io_ins_462 : _GEN_461; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_463 = 10'h1cf == io_sel ? io_ins_463 : _GEN_462; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_464 = 10'h1d0 == io_sel ? io_ins_464 : _GEN_463; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_465 = 10'h1d1 == io_sel ? io_ins_465 : _GEN_464; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_466 = 10'h1d2 == io_sel ? io_ins_466 : _GEN_465; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_467 = 10'h1d3 == io_sel ? io_ins_467 : _GEN_466; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_468 = 10'h1d4 == io_sel ? io_ins_468 : _GEN_467; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_469 = 10'h1d5 == io_sel ? io_ins_469 : _GEN_468; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_470 = 10'h1d6 == io_sel ? io_ins_470 : _GEN_469; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_471 = 10'h1d7 == io_sel ? io_ins_471 : _GEN_470; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_472 = 10'h1d8 == io_sel ? io_ins_472 : _GEN_471; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_473 = 10'h1d9 == io_sel ? io_ins_473 : _GEN_472; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_474 = 10'h1da == io_sel ? io_ins_474 : _GEN_473; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_475 = 10'h1db == io_sel ? io_ins_475 : _GEN_474; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_476 = 10'h1dc == io_sel ? io_ins_476 : _GEN_475; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_477 = 10'h1dd == io_sel ? io_ins_477 : _GEN_476; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_478 = 10'h1de == io_sel ? io_ins_478 : _GEN_477; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_479 = 10'h1df == io_sel ? io_ins_479 : _GEN_478; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_480 = 10'h1e0 == io_sel ? io_ins_480 : _GEN_479; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_481 = 10'h1e1 == io_sel ? io_ins_481 : _GEN_480; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_482 = 10'h1e2 == io_sel ? io_ins_482 : _GEN_481; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_483 = 10'h1e3 == io_sel ? io_ins_483 : _GEN_482; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_484 = 10'h1e4 == io_sel ? io_ins_484 : _GEN_483; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_485 = 10'h1e5 == io_sel ? io_ins_485 : _GEN_484; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_486 = 10'h1e6 == io_sel ? io_ins_486 : _GEN_485; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_487 = 10'h1e7 == io_sel ? io_ins_487 : _GEN_486; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_488 = 10'h1e8 == io_sel ? io_ins_488 : _GEN_487; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_489 = 10'h1e9 == io_sel ? io_ins_489 : _GEN_488; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_490 = 10'h1ea == io_sel ? io_ins_490 : _GEN_489; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_491 = 10'h1eb == io_sel ? io_ins_491 : _GEN_490; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_492 = 10'h1ec == io_sel ? io_ins_492 : _GEN_491; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_493 = 10'h1ed == io_sel ? io_ins_493 : _GEN_492; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_494 = 10'h1ee == io_sel ? io_ins_494 : _GEN_493; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_495 = 10'h1ef == io_sel ? io_ins_495 : _GEN_494; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_496 = 10'h1f0 == io_sel ? io_ins_496 : _GEN_495; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_497 = 10'h1f1 == io_sel ? io_ins_497 : _GEN_496; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_498 = 10'h1f2 == io_sel ? io_ins_498 : _GEN_497; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_499 = 10'h1f3 == io_sel ? io_ins_499 : _GEN_498; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_500 = 10'h1f4 == io_sel ? io_ins_500 : _GEN_499; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_501 = 10'h1f5 == io_sel ? io_ins_501 : _GEN_500; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_502 = 10'h1f6 == io_sel ? io_ins_502 : _GEN_501; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_503 = 10'h1f7 == io_sel ? io_ins_503 : _GEN_502; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_504 = 10'h1f8 == io_sel ? io_ins_504 : _GEN_503; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_505 = 10'h1f9 == io_sel ? io_ins_505 : _GEN_504; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_506 = 10'h1fa == io_sel ? io_ins_506 : _GEN_505; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_507 = 10'h1fb == io_sel ? io_ins_507 : _GEN_506; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_508 = 10'h1fc == io_sel ? io_ins_508 : _GEN_507; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_509 = 10'h1fd == io_sel ? io_ins_509 : _GEN_508; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_510 = 10'h1fe == io_sel ? io_ins_510 : _GEN_509; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_511 = 10'h1ff == io_sel ? io_ins_511 : _GEN_510; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_512 = 10'h200 == io_sel ? io_ins_512 : _GEN_511; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_513 = 10'h201 == io_sel ? io_ins_513 : _GEN_512; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_514 = 10'h202 == io_sel ? io_ins_514 : _GEN_513; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_515 = 10'h203 == io_sel ? io_ins_515 : _GEN_514; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_516 = 10'h204 == io_sel ? io_ins_516 : _GEN_515; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_517 = 10'h205 == io_sel ? io_ins_517 : _GEN_516; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_518 = 10'h206 == io_sel ? io_ins_518 : _GEN_517; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_519 = 10'h207 == io_sel ? io_ins_519 : _GEN_518; // @[MuxN.scala 16:10:@39796.4]
  assign _GEN_520 = 10'h208 == io_sel ? io_ins_520 : _GEN_519; // @[MuxN.scala 16:10:@39796.4]
  assign io_out = 10'h209 == io_sel ? io_ins_521 : _GEN_520; // @[MuxN.scala 16:10:@39796.4]
endmodule
module RegFile( // @[:@39798.2]
  input         clock, // @[:@39799.4]
  input         reset, // @[:@39800.4]
  input  [31:0] io_raddr, // @[:@39801.4]
  input         io_wen, // @[:@39801.4]
  input  [31:0] io_waddr, // @[:@39801.4]
  input  [63:0] io_wdata, // @[:@39801.4]
  output [63:0] io_rdata, // @[:@39801.4]
  input         io_reset, // @[:@39801.4]
  output [63:0] io_argIns_0, // @[:@39801.4]
  output [63:0] io_argIns_1, // @[:@39801.4]
  output [63:0] io_argIns_2, // @[:@39801.4]
  input         io_argOuts_0_valid, // @[:@39801.4]
  input  [63:0] io_argOuts_0_bits, // @[:@39801.4]
  input         io_argOuts_1_valid, // @[:@39801.4]
  input  [63:0] io_argOuts_1_bits, // @[:@39801.4]
  input         io_argOuts_2_valid, // @[:@39801.4]
  input  [63:0] io_argOuts_2_bits, // @[:@39801.4]
  input         io_argOuts_3_valid, // @[:@39801.4]
  input  [63:0] io_argOuts_3_bits, // @[:@39801.4]
  input         io_argOuts_4_valid, // @[:@39801.4]
  input  [63:0] io_argOuts_4_bits, // @[:@39801.4]
  input         io_argOuts_5_valid, // @[:@39801.4]
  input  [63:0] io_argOuts_5_bits, // @[:@39801.4]
  input         io_argOuts_6_valid, // @[:@39801.4]
  input  [63:0] io_argOuts_6_bits, // @[:@39801.4]
  input         io_argOuts_7_valid, // @[:@39801.4]
  input  [63:0] io_argOuts_7_bits, // @[:@39801.4]
  input         io_argOuts_8_valid, // @[:@39801.4]
  input  [63:0] io_argOuts_8_bits, // @[:@39801.4]
  input         io_argOuts_9_valid, // @[:@39801.4]
  input  [63:0] io_argOuts_9_bits, // @[:@39801.4]
  input         io_argOuts_10_valid, // @[:@39801.4]
  input  [63:0] io_argOuts_10_bits, // @[:@39801.4]
  input         io_argOuts_11_valid, // @[:@39801.4]
  input  [63:0] io_argOuts_11_bits, // @[:@39801.4]
  input         io_argOuts_12_valid, // @[:@39801.4]
  input  [63:0] io_argOuts_12_bits, // @[:@39801.4]
  input         io_argOuts_13_valid, // @[:@39801.4]
  input  [63:0] io_argOuts_13_bits, // @[:@39801.4]
  input         io_argOuts_14_valid, // @[:@39801.4]
  input  [63:0] io_argOuts_14_bits, // @[:@39801.4]
  input         io_argOuts_15_valid, // @[:@39801.4]
  input  [63:0] io_argOuts_15_bits, // @[:@39801.4]
  input         io_argOuts_16_valid, // @[:@39801.4]
  input  [63:0] io_argOuts_16_bits, // @[:@39801.4]
  input         io_argOuts_17_valid, // @[:@39801.4]
  input  [63:0] io_argOuts_17_bits, // @[:@39801.4]
  input         io_argOuts_18_valid, // @[:@39801.4]
  input  [63:0] io_argOuts_18_bits, // @[:@39801.4]
  input         io_argOuts_19_valid, // @[:@39801.4]
  input  [63:0] io_argOuts_19_bits, // @[:@39801.4]
  input         io_argOuts_20_valid, // @[:@39801.4]
  input  [63:0] io_argOuts_20_bits // @[:@39801.4]
);
  wire  regs_0_clock; // @[RegFile.scala 66:20:@41887.4]
  wire  regs_0_reset; // @[RegFile.scala 66:20:@41887.4]
  wire [63:0] regs_0_io_in; // @[RegFile.scala 66:20:@41887.4]
  wire  regs_0_io_reset; // @[RegFile.scala 66:20:@41887.4]
  wire [63:0] regs_0_io_out; // @[RegFile.scala 66:20:@41887.4]
  wire  regs_0_io_enable; // @[RegFile.scala 66:20:@41887.4]
  wire  regs_1_clock; // @[RegFile.scala 66:20:@41899.4]
  wire  regs_1_reset; // @[RegFile.scala 66:20:@41899.4]
  wire [63:0] regs_1_io_in; // @[RegFile.scala 66:20:@41899.4]
  wire  regs_1_io_reset; // @[RegFile.scala 66:20:@41899.4]
  wire [63:0] regs_1_io_out; // @[RegFile.scala 66:20:@41899.4]
  wire  regs_1_io_enable; // @[RegFile.scala 66:20:@41899.4]
  wire  regs_2_clock; // @[RegFile.scala 66:20:@41918.4]
  wire  regs_2_reset; // @[RegFile.scala 66:20:@41918.4]
  wire [63:0] regs_2_io_in; // @[RegFile.scala 66:20:@41918.4]
  wire  regs_2_io_reset; // @[RegFile.scala 66:20:@41918.4]
  wire [63:0] regs_2_io_out; // @[RegFile.scala 66:20:@41918.4]
  wire  regs_2_io_enable; // @[RegFile.scala 66:20:@41918.4]
  wire  regs_3_clock; // @[RegFile.scala 66:20:@41930.4]
  wire  regs_3_reset; // @[RegFile.scala 66:20:@41930.4]
  wire [63:0] regs_3_io_in; // @[RegFile.scala 66:20:@41930.4]
  wire  regs_3_io_reset; // @[RegFile.scala 66:20:@41930.4]
  wire [63:0] regs_3_io_out; // @[RegFile.scala 66:20:@41930.4]
  wire  regs_3_io_enable; // @[RegFile.scala 66:20:@41930.4]
  wire  regs_4_clock; // @[RegFile.scala 66:20:@41944.4]
  wire  regs_4_reset; // @[RegFile.scala 66:20:@41944.4]
  wire [63:0] regs_4_io_in; // @[RegFile.scala 66:20:@41944.4]
  wire  regs_4_io_reset; // @[RegFile.scala 66:20:@41944.4]
  wire [63:0] regs_4_io_out; // @[RegFile.scala 66:20:@41944.4]
  wire  regs_4_io_enable; // @[RegFile.scala 66:20:@41944.4]
  wire  regs_5_clock; // @[RegFile.scala 66:20:@41958.4]
  wire  regs_5_reset; // @[RegFile.scala 66:20:@41958.4]
  wire [63:0] regs_5_io_in; // @[RegFile.scala 66:20:@41958.4]
  wire  regs_5_io_reset; // @[RegFile.scala 66:20:@41958.4]
  wire [63:0] regs_5_io_out; // @[RegFile.scala 66:20:@41958.4]
  wire  regs_5_io_enable; // @[RegFile.scala 66:20:@41958.4]
  wire  regs_6_clock; // @[RegFile.scala 66:20:@41972.4]
  wire  regs_6_reset; // @[RegFile.scala 66:20:@41972.4]
  wire [63:0] regs_6_io_in; // @[RegFile.scala 66:20:@41972.4]
  wire  regs_6_io_reset; // @[RegFile.scala 66:20:@41972.4]
  wire [63:0] regs_6_io_out; // @[RegFile.scala 66:20:@41972.4]
  wire  regs_6_io_enable; // @[RegFile.scala 66:20:@41972.4]
  wire  regs_7_clock; // @[RegFile.scala 66:20:@41986.4]
  wire  regs_7_reset; // @[RegFile.scala 66:20:@41986.4]
  wire [63:0] regs_7_io_in; // @[RegFile.scala 66:20:@41986.4]
  wire  regs_7_io_reset; // @[RegFile.scala 66:20:@41986.4]
  wire [63:0] regs_7_io_out; // @[RegFile.scala 66:20:@41986.4]
  wire  regs_7_io_enable; // @[RegFile.scala 66:20:@41986.4]
  wire  regs_8_clock; // @[RegFile.scala 66:20:@42000.4]
  wire  regs_8_reset; // @[RegFile.scala 66:20:@42000.4]
  wire [63:0] regs_8_io_in; // @[RegFile.scala 66:20:@42000.4]
  wire  regs_8_io_reset; // @[RegFile.scala 66:20:@42000.4]
  wire [63:0] regs_8_io_out; // @[RegFile.scala 66:20:@42000.4]
  wire  regs_8_io_enable; // @[RegFile.scala 66:20:@42000.4]
  wire  regs_9_clock; // @[RegFile.scala 66:20:@42014.4]
  wire  regs_9_reset; // @[RegFile.scala 66:20:@42014.4]
  wire [63:0] regs_9_io_in; // @[RegFile.scala 66:20:@42014.4]
  wire  regs_9_io_reset; // @[RegFile.scala 66:20:@42014.4]
  wire [63:0] regs_9_io_out; // @[RegFile.scala 66:20:@42014.4]
  wire  regs_9_io_enable; // @[RegFile.scala 66:20:@42014.4]
  wire  regs_10_clock; // @[RegFile.scala 66:20:@42028.4]
  wire  regs_10_reset; // @[RegFile.scala 66:20:@42028.4]
  wire [63:0] regs_10_io_in; // @[RegFile.scala 66:20:@42028.4]
  wire  regs_10_io_reset; // @[RegFile.scala 66:20:@42028.4]
  wire [63:0] regs_10_io_out; // @[RegFile.scala 66:20:@42028.4]
  wire  regs_10_io_enable; // @[RegFile.scala 66:20:@42028.4]
  wire  regs_11_clock; // @[RegFile.scala 66:20:@42042.4]
  wire  regs_11_reset; // @[RegFile.scala 66:20:@42042.4]
  wire [63:0] regs_11_io_in; // @[RegFile.scala 66:20:@42042.4]
  wire  regs_11_io_reset; // @[RegFile.scala 66:20:@42042.4]
  wire [63:0] regs_11_io_out; // @[RegFile.scala 66:20:@42042.4]
  wire  regs_11_io_enable; // @[RegFile.scala 66:20:@42042.4]
  wire  regs_12_clock; // @[RegFile.scala 66:20:@42056.4]
  wire  regs_12_reset; // @[RegFile.scala 66:20:@42056.4]
  wire [63:0] regs_12_io_in; // @[RegFile.scala 66:20:@42056.4]
  wire  regs_12_io_reset; // @[RegFile.scala 66:20:@42056.4]
  wire [63:0] regs_12_io_out; // @[RegFile.scala 66:20:@42056.4]
  wire  regs_12_io_enable; // @[RegFile.scala 66:20:@42056.4]
  wire  regs_13_clock; // @[RegFile.scala 66:20:@42070.4]
  wire  regs_13_reset; // @[RegFile.scala 66:20:@42070.4]
  wire [63:0] regs_13_io_in; // @[RegFile.scala 66:20:@42070.4]
  wire  regs_13_io_reset; // @[RegFile.scala 66:20:@42070.4]
  wire [63:0] regs_13_io_out; // @[RegFile.scala 66:20:@42070.4]
  wire  regs_13_io_enable; // @[RegFile.scala 66:20:@42070.4]
  wire  regs_14_clock; // @[RegFile.scala 66:20:@42084.4]
  wire  regs_14_reset; // @[RegFile.scala 66:20:@42084.4]
  wire [63:0] regs_14_io_in; // @[RegFile.scala 66:20:@42084.4]
  wire  regs_14_io_reset; // @[RegFile.scala 66:20:@42084.4]
  wire [63:0] regs_14_io_out; // @[RegFile.scala 66:20:@42084.4]
  wire  regs_14_io_enable; // @[RegFile.scala 66:20:@42084.4]
  wire  regs_15_clock; // @[RegFile.scala 66:20:@42098.4]
  wire  regs_15_reset; // @[RegFile.scala 66:20:@42098.4]
  wire [63:0] regs_15_io_in; // @[RegFile.scala 66:20:@42098.4]
  wire  regs_15_io_reset; // @[RegFile.scala 66:20:@42098.4]
  wire [63:0] regs_15_io_out; // @[RegFile.scala 66:20:@42098.4]
  wire  regs_15_io_enable; // @[RegFile.scala 66:20:@42098.4]
  wire  regs_16_clock; // @[RegFile.scala 66:20:@42112.4]
  wire  regs_16_reset; // @[RegFile.scala 66:20:@42112.4]
  wire [63:0] regs_16_io_in; // @[RegFile.scala 66:20:@42112.4]
  wire  regs_16_io_reset; // @[RegFile.scala 66:20:@42112.4]
  wire [63:0] regs_16_io_out; // @[RegFile.scala 66:20:@42112.4]
  wire  regs_16_io_enable; // @[RegFile.scala 66:20:@42112.4]
  wire  regs_17_clock; // @[RegFile.scala 66:20:@42126.4]
  wire  regs_17_reset; // @[RegFile.scala 66:20:@42126.4]
  wire [63:0] regs_17_io_in; // @[RegFile.scala 66:20:@42126.4]
  wire  regs_17_io_reset; // @[RegFile.scala 66:20:@42126.4]
  wire [63:0] regs_17_io_out; // @[RegFile.scala 66:20:@42126.4]
  wire  regs_17_io_enable; // @[RegFile.scala 66:20:@42126.4]
  wire  regs_18_clock; // @[RegFile.scala 66:20:@42140.4]
  wire  regs_18_reset; // @[RegFile.scala 66:20:@42140.4]
  wire [63:0] regs_18_io_in; // @[RegFile.scala 66:20:@42140.4]
  wire  regs_18_io_reset; // @[RegFile.scala 66:20:@42140.4]
  wire [63:0] regs_18_io_out; // @[RegFile.scala 66:20:@42140.4]
  wire  regs_18_io_enable; // @[RegFile.scala 66:20:@42140.4]
  wire  regs_19_clock; // @[RegFile.scala 66:20:@42154.4]
  wire  regs_19_reset; // @[RegFile.scala 66:20:@42154.4]
  wire [63:0] regs_19_io_in; // @[RegFile.scala 66:20:@42154.4]
  wire  regs_19_io_reset; // @[RegFile.scala 66:20:@42154.4]
  wire [63:0] regs_19_io_out; // @[RegFile.scala 66:20:@42154.4]
  wire  regs_19_io_enable; // @[RegFile.scala 66:20:@42154.4]
  wire  regs_20_clock; // @[RegFile.scala 66:20:@42168.4]
  wire  regs_20_reset; // @[RegFile.scala 66:20:@42168.4]
  wire [63:0] regs_20_io_in; // @[RegFile.scala 66:20:@42168.4]
  wire  regs_20_io_reset; // @[RegFile.scala 66:20:@42168.4]
  wire [63:0] regs_20_io_out; // @[RegFile.scala 66:20:@42168.4]
  wire  regs_20_io_enable; // @[RegFile.scala 66:20:@42168.4]
  wire  regs_21_clock; // @[RegFile.scala 66:20:@42182.4]
  wire  regs_21_reset; // @[RegFile.scala 66:20:@42182.4]
  wire [63:0] regs_21_io_in; // @[RegFile.scala 66:20:@42182.4]
  wire  regs_21_io_reset; // @[RegFile.scala 66:20:@42182.4]
  wire [63:0] regs_21_io_out; // @[RegFile.scala 66:20:@42182.4]
  wire  regs_21_io_enable; // @[RegFile.scala 66:20:@42182.4]
  wire  regs_22_clock; // @[RegFile.scala 66:20:@42196.4]
  wire  regs_22_reset; // @[RegFile.scala 66:20:@42196.4]
  wire [63:0] regs_22_io_in; // @[RegFile.scala 66:20:@42196.4]
  wire  regs_22_io_reset; // @[RegFile.scala 66:20:@42196.4]
  wire [63:0] regs_22_io_out; // @[RegFile.scala 66:20:@42196.4]
  wire  regs_22_io_enable; // @[RegFile.scala 66:20:@42196.4]
  wire  regs_23_clock; // @[RegFile.scala 66:20:@42210.4]
  wire  regs_23_reset; // @[RegFile.scala 66:20:@42210.4]
  wire [63:0] regs_23_io_in; // @[RegFile.scala 66:20:@42210.4]
  wire  regs_23_io_reset; // @[RegFile.scala 66:20:@42210.4]
  wire [63:0] regs_23_io_out; // @[RegFile.scala 66:20:@42210.4]
  wire  regs_23_io_enable; // @[RegFile.scala 66:20:@42210.4]
  wire  regs_24_clock; // @[RegFile.scala 66:20:@42224.4]
  wire  regs_24_reset; // @[RegFile.scala 66:20:@42224.4]
  wire [63:0] regs_24_io_in; // @[RegFile.scala 66:20:@42224.4]
  wire  regs_24_io_reset; // @[RegFile.scala 66:20:@42224.4]
  wire [63:0] regs_24_io_out; // @[RegFile.scala 66:20:@42224.4]
  wire  regs_24_io_enable; // @[RegFile.scala 66:20:@42224.4]
  wire  regs_25_clock; // @[RegFile.scala 66:20:@42238.4]
  wire  regs_25_reset; // @[RegFile.scala 66:20:@42238.4]
  wire [63:0] regs_25_io_in; // @[RegFile.scala 66:20:@42238.4]
  wire  regs_25_io_reset; // @[RegFile.scala 66:20:@42238.4]
  wire [63:0] regs_25_io_out; // @[RegFile.scala 66:20:@42238.4]
  wire  regs_25_io_enable; // @[RegFile.scala 66:20:@42238.4]
  wire  regs_26_clock; // @[RegFile.scala 66:20:@42252.4]
  wire  regs_26_reset; // @[RegFile.scala 66:20:@42252.4]
  wire [63:0] regs_26_io_in; // @[RegFile.scala 66:20:@42252.4]
  wire  regs_26_io_reset; // @[RegFile.scala 66:20:@42252.4]
  wire [63:0] regs_26_io_out; // @[RegFile.scala 66:20:@42252.4]
  wire  regs_26_io_enable; // @[RegFile.scala 66:20:@42252.4]
  wire  regs_27_clock; // @[RegFile.scala 66:20:@42266.4]
  wire  regs_27_reset; // @[RegFile.scala 66:20:@42266.4]
  wire [63:0] regs_27_io_in; // @[RegFile.scala 66:20:@42266.4]
  wire  regs_27_io_reset; // @[RegFile.scala 66:20:@42266.4]
  wire [63:0] regs_27_io_out; // @[RegFile.scala 66:20:@42266.4]
  wire  regs_27_io_enable; // @[RegFile.scala 66:20:@42266.4]
  wire  regs_28_clock; // @[RegFile.scala 66:20:@42280.4]
  wire  regs_28_reset; // @[RegFile.scala 66:20:@42280.4]
  wire [63:0] regs_28_io_in; // @[RegFile.scala 66:20:@42280.4]
  wire  regs_28_io_reset; // @[RegFile.scala 66:20:@42280.4]
  wire [63:0] regs_28_io_out; // @[RegFile.scala 66:20:@42280.4]
  wire  regs_28_io_enable; // @[RegFile.scala 66:20:@42280.4]
  wire  regs_29_clock; // @[RegFile.scala 66:20:@42294.4]
  wire  regs_29_reset; // @[RegFile.scala 66:20:@42294.4]
  wire [63:0] regs_29_io_in; // @[RegFile.scala 66:20:@42294.4]
  wire  regs_29_io_reset; // @[RegFile.scala 66:20:@42294.4]
  wire [63:0] regs_29_io_out; // @[RegFile.scala 66:20:@42294.4]
  wire  regs_29_io_enable; // @[RegFile.scala 66:20:@42294.4]
  wire  regs_30_clock; // @[RegFile.scala 66:20:@42308.4]
  wire  regs_30_reset; // @[RegFile.scala 66:20:@42308.4]
  wire [63:0] regs_30_io_in; // @[RegFile.scala 66:20:@42308.4]
  wire  regs_30_io_reset; // @[RegFile.scala 66:20:@42308.4]
  wire [63:0] regs_30_io_out; // @[RegFile.scala 66:20:@42308.4]
  wire  regs_30_io_enable; // @[RegFile.scala 66:20:@42308.4]
  wire  regs_31_clock; // @[RegFile.scala 66:20:@42322.4]
  wire  regs_31_reset; // @[RegFile.scala 66:20:@42322.4]
  wire [63:0] regs_31_io_in; // @[RegFile.scala 66:20:@42322.4]
  wire  regs_31_io_reset; // @[RegFile.scala 66:20:@42322.4]
  wire [63:0] regs_31_io_out; // @[RegFile.scala 66:20:@42322.4]
  wire  regs_31_io_enable; // @[RegFile.scala 66:20:@42322.4]
  wire  regs_32_clock; // @[RegFile.scala 66:20:@42336.4]
  wire  regs_32_reset; // @[RegFile.scala 66:20:@42336.4]
  wire [63:0] regs_32_io_in; // @[RegFile.scala 66:20:@42336.4]
  wire  regs_32_io_reset; // @[RegFile.scala 66:20:@42336.4]
  wire [63:0] regs_32_io_out; // @[RegFile.scala 66:20:@42336.4]
  wire  regs_32_io_enable; // @[RegFile.scala 66:20:@42336.4]
  wire  regs_33_clock; // @[RegFile.scala 66:20:@42350.4]
  wire  regs_33_reset; // @[RegFile.scala 66:20:@42350.4]
  wire [63:0] regs_33_io_in; // @[RegFile.scala 66:20:@42350.4]
  wire  regs_33_io_reset; // @[RegFile.scala 66:20:@42350.4]
  wire [63:0] regs_33_io_out; // @[RegFile.scala 66:20:@42350.4]
  wire  regs_33_io_enable; // @[RegFile.scala 66:20:@42350.4]
  wire  regs_34_clock; // @[RegFile.scala 66:20:@42364.4]
  wire  regs_34_reset; // @[RegFile.scala 66:20:@42364.4]
  wire [63:0] regs_34_io_in; // @[RegFile.scala 66:20:@42364.4]
  wire  regs_34_io_reset; // @[RegFile.scala 66:20:@42364.4]
  wire [63:0] regs_34_io_out; // @[RegFile.scala 66:20:@42364.4]
  wire  regs_34_io_enable; // @[RegFile.scala 66:20:@42364.4]
  wire  regs_35_clock; // @[RegFile.scala 66:20:@42378.4]
  wire  regs_35_reset; // @[RegFile.scala 66:20:@42378.4]
  wire [63:0] regs_35_io_in; // @[RegFile.scala 66:20:@42378.4]
  wire  regs_35_io_reset; // @[RegFile.scala 66:20:@42378.4]
  wire [63:0] regs_35_io_out; // @[RegFile.scala 66:20:@42378.4]
  wire  regs_35_io_enable; // @[RegFile.scala 66:20:@42378.4]
  wire  regs_36_clock; // @[RegFile.scala 66:20:@42392.4]
  wire  regs_36_reset; // @[RegFile.scala 66:20:@42392.4]
  wire [63:0] regs_36_io_in; // @[RegFile.scala 66:20:@42392.4]
  wire  regs_36_io_reset; // @[RegFile.scala 66:20:@42392.4]
  wire [63:0] regs_36_io_out; // @[RegFile.scala 66:20:@42392.4]
  wire  regs_36_io_enable; // @[RegFile.scala 66:20:@42392.4]
  wire  regs_37_clock; // @[RegFile.scala 66:20:@42406.4]
  wire  regs_37_reset; // @[RegFile.scala 66:20:@42406.4]
  wire [63:0] regs_37_io_in; // @[RegFile.scala 66:20:@42406.4]
  wire  regs_37_io_reset; // @[RegFile.scala 66:20:@42406.4]
  wire [63:0] regs_37_io_out; // @[RegFile.scala 66:20:@42406.4]
  wire  regs_37_io_enable; // @[RegFile.scala 66:20:@42406.4]
  wire  regs_38_clock; // @[RegFile.scala 66:20:@42420.4]
  wire  regs_38_reset; // @[RegFile.scala 66:20:@42420.4]
  wire [63:0] regs_38_io_in; // @[RegFile.scala 66:20:@42420.4]
  wire  regs_38_io_reset; // @[RegFile.scala 66:20:@42420.4]
  wire [63:0] regs_38_io_out; // @[RegFile.scala 66:20:@42420.4]
  wire  regs_38_io_enable; // @[RegFile.scala 66:20:@42420.4]
  wire  regs_39_clock; // @[RegFile.scala 66:20:@42434.4]
  wire  regs_39_reset; // @[RegFile.scala 66:20:@42434.4]
  wire [63:0] regs_39_io_in; // @[RegFile.scala 66:20:@42434.4]
  wire  regs_39_io_reset; // @[RegFile.scala 66:20:@42434.4]
  wire [63:0] regs_39_io_out; // @[RegFile.scala 66:20:@42434.4]
  wire  regs_39_io_enable; // @[RegFile.scala 66:20:@42434.4]
  wire  regs_40_clock; // @[RegFile.scala 66:20:@42448.4]
  wire  regs_40_reset; // @[RegFile.scala 66:20:@42448.4]
  wire [63:0] regs_40_io_in; // @[RegFile.scala 66:20:@42448.4]
  wire  regs_40_io_reset; // @[RegFile.scala 66:20:@42448.4]
  wire [63:0] regs_40_io_out; // @[RegFile.scala 66:20:@42448.4]
  wire  regs_40_io_enable; // @[RegFile.scala 66:20:@42448.4]
  wire  regs_41_clock; // @[RegFile.scala 66:20:@42462.4]
  wire  regs_41_reset; // @[RegFile.scala 66:20:@42462.4]
  wire [63:0] regs_41_io_in; // @[RegFile.scala 66:20:@42462.4]
  wire  regs_41_io_reset; // @[RegFile.scala 66:20:@42462.4]
  wire [63:0] regs_41_io_out; // @[RegFile.scala 66:20:@42462.4]
  wire  regs_41_io_enable; // @[RegFile.scala 66:20:@42462.4]
  wire  regs_42_clock; // @[RegFile.scala 66:20:@42476.4]
  wire  regs_42_reset; // @[RegFile.scala 66:20:@42476.4]
  wire [63:0] regs_42_io_in; // @[RegFile.scala 66:20:@42476.4]
  wire  regs_42_io_reset; // @[RegFile.scala 66:20:@42476.4]
  wire [63:0] regs_42_io_out; // @[RegFile.scala 66:20:@42476.4]
  wire  regs_42_io_enable; // @[RegFile.scala 66:20:@42476.4]
  wire  regs_43_clock; // @[RegFile.scala 66:20:@42490.4]
  wire  regs_43_reset; // @[RegFile.scala 66:20:@42490.4]
  wire [63:0] regs_43_io_in; // @[RegFile.scala 66:20:@42490.4]
  wire  regs_43_io_reset; // @[RegFile.scala 66:20:@42490.4]
  wire [63:0] regs_43_io_out; // @[RegFile.scala 66:20:@42490.4]
  wire  regs_43_io_enable; // @[RegFile.scala 66:20:@42490.4]
  wire  regs_44_clock; // @[RegFile.scala 66:20:@42504.4]
  wire  regs_44_reset; // @[RegFile.scala 66:20:@42504.4]
  wire [63:0] regs_44_io_in; // @[RegFile.scala 66:20:@42504.4]
  wire  regs_44_io_reset; // @[RegFile.scala 66:20:@42504.4]
  wire [63:0] regs_44_io_out; // @[RegFile.scala 66:20:@42504.4]
  wire  regs_44_io_enable; // @[RegFile.scala 66:20:@42504.4]
  wire  regs_45_clock; // @[RegFile.scala 66:20:@42518.4]
  wire  regs_45_reset; // @[RegFile.scala 66:20:@42518.4]
  wire [63:0] regs_45_io_in; // @[RegFile.scala 66:20:@42518.4]
  wire  regs_45_io_reset; // @[RegFile.scala 66:20:@42518.4]
  wire [63:0] regs_45_io_out; // @[RegFile.scala 66:20:@42518.4]
  wire  regs_45_io_enable; // @[RegFile.scala 66:20:@42518.4]
  wire  regs_46_clock; // @[RegFile.scala 66:20:@42532.4]
  wire  regs_46_reset; // @[RegFile.scala 66:20:@42532.4]
  wire [63:0] regs_46_io_in; // @[RegFile.scala 66:20:@42532.4]
  wire  regs_46_io_reset; // @[RegFile.scala 66:20:@42532.4]
  wire [63:0] regs_46_io_out; // @[RegFile.scala 66:20:@42532.4]
  wire  regs_46_io_enable; // @[RegFile.scala 66:20:@42532.4]
  wire  regs_47_clock; // @[RegFile.scala 66:20:@42546.4]
  wire  regs_47_reset; // @[RegFile.scala 66:20:@42546.4]
  wire [63:0] regs_47_io_in; // @[RegFile.scala 66:20:@42546.4]
  wire  regs_47_io_reset; // @[RegFile.scala 66:20:@42546.4]
  wire [63:0] regs_47_io_out; // @[RegFile.scala 66:20:@42546.4]
  wire  regs_47_io_enable; // @[RegFile.scala 66:20:@42546.4]
  wire  regs_48_clock; // @[RegFile.scala 66:20:@42560.4]
  wire  regs_48_reset; // @[RegFile.scala 66:20:@42560.4]
  wire [63:0] regs_48_io_in; // @[RegFile.scala 66:20:@42560.4]
  wire  regs_48_io_reset; // @[RegFile.scala 66:20:@42560.4]
  wire [63:0] regs_48_io_out; // @[RegFile.scala 66:20:@42560.4]
  wire  regs_48_io_enable; // @[RegFile.scala 66:20:@42560.4]
  wire  regs_49_clock; // @[RegFile.scala 66:20:@42574.4]
  wire  regs_49_reset; // @[RegFile.scala 66:20:@42574.4]
  wire [63:0] regs_49_io_in; // @[RegFile.scala 66:20:@42574.4]
  wire  regs_49_io_reset; // @[RegFile.scala 66:20:@42574.4]
  wire [63:0] regs_49_io_out; // @[RegFile.scala 66:20:@42574.4]
  wire  regs_49_io_enable; // @[RegFile.scala 66:20:@42574.4]
  wire  regs_50_clock; // @[RegFile.scala 66:20:@42588.4]
  wire  regs_50_reset; // @[RegFile.scala 66:20:@42588.4]
  wire [63:0] regs_50_io_in; // @[RegFile.scala 66:20:@42588.4]
  wire  regs_50_io_reset; // @[RegFile.scala 66:20:@42588.4]
  wire [63:0] regs_50_io_out; // @[RegFile.scala 66:20:@42588.4]
  wire  regs_50_io_enable; // @[RegFile.scala 66:20:@42588.4]
  wire  regs_51_clock; // @[RegFile.scala 66:20:@42602.4]
  wire  regs_51_reset; // @[RegFile.scala 66:20:@42602.4]
  wire [63:0] regs_51_io_in; // @[RegFile.scala 66:20:@42602.4]
  wire  regs_51_io_reset; // @[RegFile.scala 66:20:@42602.4]
  wire [63:0] regs_51_io_out; // @[RegFile.scala 66:20:@42602.4]
  wire  regs_51_io_enable; // @[RegFile.scala 66:20:@42602.4]
  wire  regs_52_clock; // @[RegFile.scala 66:20:@42616.4]
  wire  regs_52_reset; // @[RegFile.scala 66:20:@42616.4]
  wire [63:0] regs_52_io_in; // @[RegFile.scala 66:20:@42616.4]
  wire  regs_52_io_reset; // @[RegFile.scala 66:20:@42616.4]
  wire [63:0] regs_52_io_out; // @[RegFile.scala 66:20:@42616.4]
  wire  regs_52_io_enable; // @[RegFile.scala 66:20:@42616.4]
  wire  regs_53_clock; // @[RegFile.scala 66:20:@42630.4]
  wire  regs_53_reset; // @[RegFile.scala 66:20:@42630.4]
  wire [63:0] regs_53_io_in; // @[RegFile.scala 66:20:@42630.4]
  wire  regs_53_io_reset; // @[RegFile.scala 66:20:@42630.4]
  wire [63:0] regs_53_io_out; // @[RegFile.scala 66:20:@42630.4]
  wire  regs_53_io_enable; // @[RegFile.scala 66:20:@42630.4]
  wire  regs_54_clock; // @[RegFile.scala 66:20:@42644.4]
  wire  regs_54_reset; // @[RegFile.scala 66:20:@42644.4]
  wire [63:0] regs_54_io_in; // @[RegFile.scala 66:20:@42644.4]
  wire  regs_54_io_reset; // @[RegFile.scala 66:20:@42644.4]
  wire [63:0] regs_54_io_out; // @[RegFile.scala 66:20:@42644.4]
  wire  regs_54_io_enable; // @[RegFile.scala 66:20:@42644.4]
  wire  regs_55_clock; // @[RegFile.scala 66:20:@42658.4]
  wire  regs_55_reset; // @[RegFile.scala 66:20:@42658.4]
  wire [63:0] regs_55_io_in; // @[RegFile.scala 66:20:@42658.4]
  wire  regs_55_io_reset; // @[RegFile.scala 66:20:@42658.4]
  wire [63:0] regs_55_io_out; // @[RegFile.scala 66:20:@42658.4]
  wire  regs_55_io_enable; // @[RegFile.scala 66:20:@42658.4]
  wire  regs_56_clock; // @[RegFile.scala 66:20:@42672.4]
  wire  regs_56_reset; // @[RegFile.scala 66:20:@42672.4]
  wire [63:0] regs_56_io_in; // @[RegFile.scala 66:20:@42672.4]
  wire  regs_56_io_reset; // @[RegFile.scala 66:20:@42672.4]
  wire [63:0] regs_56_io_out; // @[RegFile.scala 66:20:@42672.4]
  wire  regs_56_io_enable; // @[RegFile.scala 66:20:@42672.4]
  wire  regs_57_clock; // @[RegFile.scala 66:20:@42686.4]
  wire  regs_57_reset; // @[RegFile.scala 66:20:@42686.4]
  wire [63:0] regs_57_io_in; // @[RegFile.scala 66:20:@42686.4]
  wire  regs_57_io_reset; // @[RegFile.scala 66:20:@42686.4]
  wire [63:0] regs_57_io_out; // @[RegFile.scala 66:20:@42686.4]
  wire  regs_57_io_enable; // @[RegFile.scala 66:20:@42686.4]
  wire  regs_58_clock; // @[RegFile.scala 66:20:@42700.4]
  wire  regs_58_reset; // @[RegFile.scala 66:20:@42700.4]
  wire [63:0] regs_58_io_in; // @[RegFile.scala 66:20:@42700.4]
  wire  regs_58_io_reset; // @[RegFile.scala 66:20:@42700.4]
  wire [63:0] regs_58_io_out; // @[RegFile.scala 66:20:@42700.4]
  wire  regs_58_io_enable; // @[RegFile.scala 66:20:@42700.4]
  wire  regs_59_clock; // @[RegFile.scala 66:20:@42714.4]
  wire  regs_59_reset; // @[RegFile.scala 66:20:@42714.4]
  wire [63:0] regs_59_io_in; // @[RegFile.scala 66:20:@42714.4]
  wire  regs_59_io_reset; // @[RegFile.scala 66:20:@42714.4]
  wire [63:0] regs_59_io_out; // @[RegFile.scala 66:20:@42714.4]
  wire  regs_59_io_enable; // @[RegFile.scala 66:20:@42714.4]
  wire  regs_60_clock; // @[RegFile.scala 66:20:@42728.4]
  wire  regs_60_reset; // @[RegFile.scala 66:20:@42728.4]
  wire [63:0] regs_60_io_in; // @[RegFile.scala 66:20:@42728.4]
  wire  regs_60_io_reset; // @[RegFile.scala 66:20:@42728.4]
  wire [63:0] regs_60_io_out; // @[RegFile.scala 66:20:@42728.4]
  wire  regs_60_io_enable; // @[RegFile.scala 66:20:@42728.4]
  wire  regs_61_clock; // @[RegFile.scala 66:20:@42742.4]
  wire  regs_61_reset; // @[RegFile.scala 66:20:@42742.4]
  wire [63:0] regs_61_io_in; // @[RegFile.scala 66:20:@42742.4]
  wire  regs_61_io_reset; // @[RegFile.scala 66:20:@42742.4]
  wire [63:0] regs_61_io_out; // @[RegFile.scala 66:20:@42742.4]
  wire  regs_61_io_enable; // @[RegFile.scala 66:20:@42742.4]
  wire  regs_62_clock; // @[RegFile.scala 66:20:@42756.4]
  wire  regs_62_reset; // @[RegFile.scala 66:20:@42756.4]
  wire [63:0] regs_62_io_in; // @[RegFile.scala 66:20:@42756.4]
  wire  regs_62_io_reset; // @[RegFile.scala 66:20:@42756.4]
  wire [63:0] regs_62_io_out; // @[RegFile.scala 66:20:@42756.4]
  wire  regs_62_io_enable; // @[RegFile.scala 66:20:@42756.4]
  wire  regs_63_clock; // @[RegFile.scala 66:20:@42770.4]
  wire  regs_63_reset; // @[RegFile.scala 66:20:@42770.4]
  wire [63:0] regs_63_io_in; // @[RegFile.scala 66:20:@42770.4]
  wire  regs_63_io_reset; // @[RegFile.scala 66:20:@42770.4]
  wire [63:0] regs_63_io_out; // @[RegFile.scala 66:20:@42770.4]
  wire  regs_63_io_enable; // @[RegFile.scala 66:20:@42770.4]
  wire  regs_64_clock; // @[RegFile.scala 66:20:@42784.4]
  wire  regs_64_reset; // @[RegFile.scala 66:20:@42784.4]
  wire [63:0] regs_64_io_in; // @[RegFile.scala 66:20:@42784.4]
  wire  regs_64_io_reset; // @[RegFile.scala 66:20:@42784.4]
  wire [63:0] regs_64_io_out; // @[RegFile.scala 66:20:@42784.4]
  wire  regs_64_io_enable; // @[RegFile.scala 66:20:@42784.4]
  wire  regs_65_clock; // @[RegFile.scala 66:20:@42798.4]
  wire  regs_65_reset; // @[RegFile.scala 66:20:@42798.4]
  wire [63:0] regs_65_io_in; // @[RegFile.scala 66:20:@42798.4]
  wire  regs_65_io_reset; // @[RegFile.scala 66:20:@42798.4]
  wire [63:0] regs_65_io_out; // @[RegFile.scala 66:20:@42798.4]
  wire  regs_65_io_enable; // @[RegFile.scala 66:20:@42798.4]
  wire  regs_66_clock; // @[RegFile.scala 66:20:@42812.4]
  wire  regs_66_reset; // @[RegFile.scala 66:20:@42812.4]
  wire [63:0] regs_66_io_in; // @[RegFile.scala 66:20:@42812.4]
  wire  regs_66_io_reset; // @[RegFile.scala 66:20:@42812.4]
  wire [63:0] regs_66_io_out; // @[RegFile.scala 66:20:@42812.4]
  wire  regs_66_io_enable; // @[RegFile.scala 66:20:@42812.4]
  wire  regs_67_clock; // @[RegFile.scala 66:20:@42826.4]
  wire  regs_67_reset; // @[RegFile.scala 66:20:@42826.4]
  wire [63:0] regs_67_io_in; // @[RegFile.scala 66:20:@42826.4]
  wire  regs_67_io_reset; // @[RegFile.scala 66:20:@42826.4]
  wire [63:0] regs_67_io_out; // @[RegFile.scala 66:20:@42826.4]
  wire  regs_67_io_enable; // @[RegFile.scala 66:20:@42826.4]
  wire  regs_68_clock; // @[RegFile.scala 66:20:@42840.4]
  wire  regs_68_reset; // @[RegFile.scala 66:20:@42840.4]
  wire [63:0] regs_68_io_in; // @[RegFile.scala 66:20:@42840.4]
  wire  regs_68_io_reset; // @[RegFile.scala 66:20:@42840.4]
  wire [63:0] regs_68_io_out; // @[RegFile.scala 66:20:@42840.4]
  wire  regs_68_io_enable; // @[RegFile.scala 66:20:@42840.4]
  wire  regs_69_clock; // @[RegFile.scala 66:20:@42854.4]
  wire  regs_69_reset; // @[RegFile.scala 66:20:@42854.4]
  wire [63:0] regs_69_io_in; // @[RegFile.scala 66:20:@42854.4]
  wire  regs_69_io_reset; // @[RegFile.scala 66:20:@42854.4]
  wire [63:0] regs_69_io_out; // @[RegFile.scala 66:20:@42854.4]
  wire  regs_69_io_enable; // @[RegFile.scala 66:20:@42854.4]
  wire  regs_70_clock; // @[RegFile.scala 66:20:@42868.4]
  wire  regs_70_reset; // @[RegFile.scala 66:20:@42868.4]
  wire [63:0] regs_70_io_in; // @[RegFile.scala 66:20:@42868.4]
  wire  regs_70_io_reset; // @[RegFile.scala 66:20:@42868.4]
  wire [63:0] regs_70_io_out; // @[RegFile.scala 66:20:@42868.4]
  wire  regs_70_io_enable; // @[RegFile.scala 66:20:@42868.4]
  wire  regs_71_clock; // @[RegFile.scala 66:20:@42882.4]
  wire  regs_71_reset; // @[RegFile.scala 66:20:@42882.4]
  wire [63:0] regs_71_io_in; // @[RegFile.scala 66:20:@42882.4]
  wire  regs_71_io_reset; // @[RegFile.scala 66:20:@42882.4]
  wire [63:0] regs_71_io_out; // @[RegFile.scala 66:20:@42882.4]
  wire  regs_71_io_enable; // @[RegFile.scala 66:20:@42882.4]
  wire  regs_72_clock; // @[RegFile.scala 66:20:@42896.4]
  wire  regs_72_reset; // @[RegFile.scala 66:20:@42896.4]
  wire [63:0] regs_72_io_in; // @[RegFile.scala 66:20:@42896.4]
  wire  regs_72_io_reset; // @[RegFile.scala 66:20:@42896.4]
  wire [63:0] regs_72_io_out; // @[RegFile.scala 66:20:@42896.4]
  wire  regs_72_io_enable; // @[RegFile.scala 66:20:@42896.4]
  wire  regs_73_clock; // @[RegFile.scala 66:20:@42910.4]
  wire  regs_73_reset; // @[RegFile.scala 66:20:@42910.4]
  wire [63:0] regs_73_io_in; // @[RegFile.scala 66:20:@42910.4]
  wire  regs_73_io_reset; // @[RegFile.scala 66:20:@42910.4]
  wire [63:0] regs_73_io_out; // @[RegFile.scala 66:20:@42910.4]
  wire  regs_73_io_enable; // @[RegFile.scala 66:20:@42910.4]
  wire  regs_74_clock; // @[RegFile.scala 66:20:@42924.4]
  wire  regs_74_reset; // @[RegFile.scala 66:20:@42924.4]
  wire [63:0] regs_74_io_in; // @[RegFile.scala 66:20:@42924.4]
  wire  regs_74_io_reset; // @[RegFile.scala 66:20:@42924.4]
  wire [63:0] regs_74_io_out; // @[RegFile.scala 66:20:@42924.4]
  wire  regs_74_io_enable; // @[RegFile.scala 66:20:@42924.4]
  wire  regs_75_clock; // @[RegFile.scala 66:20:@42938.4]
  wire  regs_75_reset; // @[RegFile.scala 66:20:@42938.4]
  wire [63:0] regs_75_io_in; // @[RegFile.scala 66:20:@42938.4]
  wire  regs_75_io_reset; // @[RegFile.scala 66:20:@42938.4]
  wire [63:0] regs_75_io_out; // @[RegFile.scala 66:20:@42938.4]
  wire  regs_75_io_enable; // @[RegFile.scala 66:20:@42938.4]
  wire  regs_76_clock; // @[RegFile.scala 66:20:@42952.4]
  wire  regs_76_reset; // @[RegFile.scala 66:20:@42952.4]
  wire [63:0] regs_76_io_in; // @[RegFile.scala 66:20:@42952.4]
  wire  regs_76_io_reset; // @[RegFile.scala 66:20:@42952.4]
  wire [63:0] regs_76_io_out; // @[RegFile.scala 66:20:@42952.4]
  wire  regs_76_io_enable; // @[RegFile.scala 66:20:@42952.4]
  wire  regs_77_clock; // @[RegFile.scala 66:20:@42966.4]
  wire  regs_77_reset; // @[RegFile.scala 66:20:@42966.4]
  wire [63:0] regs_77_io_in; // @[RegFile.scala 66:20:@42966.4]
  wire  regs_77_io_reset; // @[RegFile.scala 66:20:@42966.4]
  wire [63:0] regs_77_io_out; // @[RegFile.scala 66:20:@42966.4]
  wire  regs_77_io_enable; // @[RegFile.scala 66:20:@42966.4]
  wire  regs_78_clock; // @[RegFile.scala 66:20:@42980.4]
  wire  regs_78_reset; // @[RegFile.scala 66:20:@42980.4]
  wire [63:0] regs_78_io_in; // @[RegFile.scala 66:20:@42980.4]
  wire  regs_78_io_reset; // @[RegFile.scala 66:20:@42980.4]
  wire [63:0] regs_78_io_out; // @[RegFile.scala 66:20:@42980.4]
  wire  regs_78_io_enable; // @[RegFile.scala 66:20:@42980.4]
  wire  regs_79_clock; // @[RegFile.scala 66:20:@42994.4]
  wire  regs_79_reset; // @[RegFile.scala 66:20:@42994.4]
  wire [63:0] regs_79_io_in; // @[RegFile.scala 66:20:@42994.4]
  wire  regs_79_io_reset; // @[RegFile.scala 66:20:@42994.4]
  wire [63:0] regs_79_io_out; // @[RegFile.scala 66:20:@42994.4]
  wire  regs_79_io_enable; // @[RegFile.scala 66:20:@42994.4]
  wire  regs_80_clock; // @[RegFile.scala 66:20:@43008.4]
  wire  regs_80_reset; // @[RegFile.scala 66:20:@43008.4]
  wire [63:0] regs_80_io_in; // @[RegFile.scala 66:20:@43008.4]
  wire  regs_80_io_reset; // @[RegFile.scala 66:20:@43008.4]
  wire [63:0] regs_80_io_out; // @[RegFile.scala 66:20:@43008.4]
  wire  regs_80_io_enable; // @[RegFile.scala 66:20:@43008.4]
  wire  regs_81_clock; // @[RegFile.scala 66:20:@43022.4]
  wire  regs_81_reset; // @[RegFile.scala 66:20:@43022.4]
  wire [63:0] regs_81_io_in; // @[RegFile.scala 66:20:@43022.4]
  wire  regs_81_io_reset; // @[RegFile.scala 66:20:@43022.4]
  wire [63:0] regs_81_io_out; // @[RegFile.scala 66:20:@43022.4]
  wire  regs_81_io_enable; // @[RegFile.scala 66:20:@43022.4]
  wire  regs_82_clock; // @[RegFile.scala 66:20:@43036.4]
  wire  regs_82_reset; // @[RegFile.scala 66:20:@43036.4]
  wire [63:0] regs_82_io_in; // @[RegFile.scala 66:20:@43036.4]
  wire  regs_82_io_reset; // @[RegFile.scala 66:20:@43036.4]
  wire [63:0] regs_82_io_out; // @[RegFile.scala 66:20:@43036.4]
  wire  regs_82_io_enable; // @[RegFile.scala 66:20:@43036.4]
  wire  regs_83_clock; // @[RegFile.scala 66:20:@43050.4]
  wire  regs_83_reset; // @[RegFile.scala 66:20:@43050.4]
  wire [63:0] regs_83_io_in; // @[RegFile.scala 66:20:@43050.4]
  wire  regs_83_io_reset; // @[RegFile.scala 66:20:@43050.4]
  wire [63:0] regs_83_io_out; // @[RegFile.scala 66:20:@43050.4]
  wire  regs_83_io_enable; // @[RegFile.scala 66:20:@43050.4]
  wire  regs_84_clock; // @[RegFile.scala 66:20:@43064.4]
  wire  regs_84_reset; // @[RegFile.scala 66:20:@43064.4]
  wire [63:0] regs_84_io_in; // @[RegFile.scala 66:20:@43064.4]
  wire  regs_84_io_reset; // @[RegFile.scala 66:20:@43064.4]
  wire [63:0] regs_84_io_out; // @[RegFile.scala 66:20:@43064.4]
  wire  regs_84_io_enable; // @[RegFile.scala 66:20:@43064.4]
  wire  regs_85_clock; // @[RegFile.scala 66:20:@43078.4]
  wire  regs_85_reset; // @[RegFile.scala 66:20:@43078.4]
  wire [63:0] regs_85_io_in; // @[RegFile.scala 66:20:@43078.4]
  wire  regs_85_io_reset; // @[RegFile.scala 66:20:@43078.4]
  wire [63:0] regs_85_io_out; // @[RegFile.scala 66:20:@43078.4]
  wire  regs_85_io_enable; // @[RegFile.scala 66:20:@43078.4]
  wire  regs_86_clock; // @[RegFile.scala 66:20:@43092.4]
  wire  regs_86_reset; // @[RegFile.scala 66:20:@43092.4]
  wire [63:0] regs_86_io_in; // @[RegFile.scala 66:20:@43092.4]
  wire  regs_86_io_reset; // @[RegFile.scala 66:20:@43092.4]
  wire [63:0] regs_86_io_out; // @[RegFile.scala 66:20:@43092.4]
  wire  regs_86_io_enable; // @[RegFile.scala 66:20:@43092.4]
  wire  regs_87_clock; // @[RegFile.scala 66:20:@43106.4]
  wire  regs_87_reset; // @[RegFile.scala 66:20:@43106.4]
  wire [63:0] regs_87_io_in; // @[RegFile.scala 66:20:@43106.4]
  wire  regs_87_io_reset; // @[RegFile.scala 66:20:@43106.4]
  wire [63:0] regs_87_io_out; // @[RegFile.scala 66:20:@43106.4]
  wire  regs_87_io_enable; // @[RegFile.scala 66:20:@43106.4]
  wire  regs_88_clock; // @[RegFile.scala 66:20:@43120.4]
  wire  regs_88_reset; // @[RegFile.scala 66:20:@43120.4]
  wire [63:0] regs_88_io_in; // @[RegFile.scala 66:20:@43120.4]
  wire  regs_88_io_reset; // @[RegFile.scala 66:20:@43120.4]
  wire [63:0] regs_88_io_out; // @[RegFile.scala 66:20:@43120.4]
  wire  regs_88_io_enable; // @[RegFile.scala 66:20:@43120.4]
  wire  regs_89_clock; // @[RegFile.scala 66:20:@43134.4]
  wire  regs_89_reset; // @[RegFile.scala 66:20:@43134.4]
  wire [63:0] regs_89_io_in; // @[RegFile.scala 66:20:@43134.4]
  wire  regs_89_io_reset; // @[RegFile.scala 66:20:@43134.4]
  wire [63:0] regs_89_io_out; // @[RegFile.scala 66:20:@43134.4]
  wire  regs_89_io_enable; // @[RegFile.scala 66:20:@43134.4]
  wire  regs_90_clock; // @[RegFile.scala 66:20:@43148.4]
  wire  regs_90_reset; // @[RegFile.scala 66:20:@43148.4]
  wire [63:0] regs_90_io_in; // @[RegFile.scala 66:20:@43148.4]
  wire  regs_90_io_reset; // @[RegFile.scala 66:20:@43148.4]
  wire [63:0] regs_90_io_out; // @[RegFile.scala 66:20:@43148.4]
  wire  regs_90_io_enable; // @[RegFile.scala 66:20:@43148.4]
  wire  regs_91_clock; // @[RegFile.scala 66:20:@43162.4]
  wire  regs_91_reset; // @[RegFile.scala 66:20:@43162.4]
  wire [63:0] regs_91_io_in; // @[RegFile.scala 66:20:@43162.4]
  wire  regs_91_io_reset; // @[RegFile.scala 66:20:@43162.4]
  wire [63:0] regs_91_io_out; // @[RegFile.scala 66:20:@43162.4]
  wire  regs_91_io_enable; // @[RegFile.scala 66:20:@43162.4]
  wire  regs_92_clock; // @[RegFile.scala 66:20:@43176.4]
  wire  regs_92_reset; // @[RegFile.scala 66:20:@43176.4]
  wire [63:0] regs_92_io_in; // @[RegFile.scala 66:20:@43176.4]
  wire  regs_92_io_reset; // @[RegFile.scala 66:20:@43176.4]
  wire [63:0] regs_92_io_out; // @[RegFile.scala 66:20:@43176.4]
  wire  regs_92_io_enable; // @[RegFile.scala 66:20:@43176.4]
  wire  regs_93_clock; // @[RegFile.scala 66:20:@43190.4]
  wire  regs_93_reset; // @[RegFile.scala 66:20:@43190.4]
  wire [63:0] regs_93_io_in; // @[RegFile.scala 66:20:@43190.4]
  wire  regs_93_io_reset; // @[RegFile.scala 66:20:@43190.4]
  wire [63:0] regs_93_io_out; // @[RegFile.scala 66:20:@43190.4]
  wire  regs_93_io_enable; // @[RegFile.scala 66:20:@43190.4]
  wire  regs_94_clock; // @[RegFile.scala 66:20:@43204.4]
  wire  regs_94_reset; // @[RegFile.scala 66:20:@43204.4]
  wire [63:0] regs_94_io_in; // @[RegFile.scala 66:20:@43204.4]
  wire  regs_94_io_reset; // @[RegFile.scala 66:20:@43204.4]
  wire [63:0] regs_94_io_out; // @[RegFile.scala 66:20:@43204.4]
  wire  regs_94_io_enable; // @[RegFile.scala 66:20:@43204.4]
  wire  regs_95_clock; // @[RegFile.scala 66:20:@43218.4]
  wire  regs_95_reset; // @[RegFile.scala 66:20:@43218.4]
  wire [63:0] regs_95_io_in; // @[RegFile.scala 66:20:@43218.4]
  wire  regs_95_io_reset; // @[RegFile.scala 66:20:@43218.4]
  wire [63:0] regs_95_io_out; // @[RegFile.scala 66:20:@43218.4]
  wire  regs_95_io_enable; // @[RegFile.scala 66:20:@43218.4]
  wire  regs_96_clock; // @[RegFile.scala 66:20:@43232.4]
  wire  regs_96_reset; // @[RegFile.scala 66:20:@43232.4]
  wire [63:0] regs_96_io_in; // @[RegFile.scala 66:20:@43232.4]
  wire  regs_96_io_reset; // @[RegFile.scala 66:20:@43232.4]
  wire [63:0] regs_96_io_out; // @[RegFile.scala 66:20:@43232.4]
  wire  regs_96_io_enable; // @[RegFile.scala 66:20:@43232.4]
  wire  regs_97_clock; // @[RegFile.scala 66:20:@43246.4]
  wire  regs_97_reset; // @[RegFile.scala 66:20:@43246.4]
  wire [63:0] regs_97_io_in; // @[RegFile.scala 66:20:@43246.4]
  wire  regs_97_io_reset; // @[RegFile.scala 66:20:@43246.4]
  wire [63:0] regs_97_io_out; // @[RegFile.scala 66:20:@43246.4]
  wire  regs_97_io_enable; // @[RegFile.scala 66:20:@43246.4]
  wire  regs_98_clock; // @[RegFile.scala 66:20:@43260.4]
  wire  regs_98_reset; // @[RegFile.scala 66:20:@43260.4]
  wire [63:0] regs_98_io_in; // @[RegFile.scala 66:20:@43260.4]
  wire  regs_98_io_reset; // @[RegFile.scala 66:20:@43260.4]
  wire [63:0] regs_98_io_out; // @[RegFile.scala 66:20:@43260.4]
  wire  regs_98_io_enable; // @[RegFile.scala 66:20:@43260.4]
  wire  regs_99_clock; // @[RegFile.scala 66:20:@43274.4]
  wire  regs_99_reset; // @[RegFile.scala 66:20:@43274.4]
  wire [63:0] regs_99_io_in; // @[RegFile.scala 66:20:@43274.4]
  wire  regs_99_io_reset; // @[RegFile.scala 66:20:@43274.4]
  wire [63:0] regs_99_io_out; // @[RegFile.scala 66:20:@43274.4]
  wire  regs_99_io_enable; // @[RegFile.scala 66:20:@43274.4]
  wire  regs_100_clock; // @[RegFile.scala 66:20:@43288.4]
  wire  regs_100_reset; // @[RegFile.scala 66:20:@43288.4]
  wire [63:0] regs_100_io_in; // @[RegFile.scala 66:20:@43288.4]
  wire  regs_100_io_reset; // @[RegFile.scala 66:20:@43288.4]
  wire [63:0] regs_100_io_out; // @[RegFile.scala 66:20:@43288.4]
  wire  regs_100_io_enable; // @[RegFile.scala 66:20:@43288.4]
  wire  regs_101_clock; // @[RegFile.scala 66:20:@43302.4]
  wire  regs_101_reset; // @[RegFile.scala 66:20:@43302.4]
  wire [63:0] regs_101_io_in; // @[RegFile.scala 66:20:@43302.4]
  wire  regs_101_io_reset; // @[RegFile.scala 66:20:@43302.4]
  wire [63:0] regs_101_io_out; // @[RegFile.scala 66:20:@43302.4]
  wire  regs_101_io_enable; // @[RegFile.scala 66:20:@43302.4]
  wire  regs_102_clock; // @[RegFile.scala 66:20:@43316.4]
  wire  regs_102_reset; // @[RegFile.scala 66:20:@43316.4]
  wire [63:0] regs_102_io_in; // @[RegFile.scala 66:20:@43316.4]
  wire  regs_102_io_reset; // @[RegFile.scala 66:20:@43316.4]
  wire [63:0] regs_102_io_out; // @[RegFile.scala 66:20:@43316.4]
  wire  regs_102_io_enable; // @[RegFile.scala 66:20:@43316.4]
  wire  regs_103_clock; // @[RegFile.scala 66:20:@43330.4]
  wire  regs_103_reset; // @[RegFile.scala 66:20:@43330.4]
  wire [63:0] regs_103_io_in; // @[RegFile.scala 66:20:@43330.4]
  wire  regs_103_io_reset; // @[RegFile.scala 66:20:@43330.4]
  wire [63:0] regs_103_io_out; // @[RegFile.scala 66:20:@43330.4]
  wire  regs_103_io_enable; // @[RegFile.scala 66:20:@43330.4]
  wire  regs_104_clock; // @[RegFile.scala 66:20:@43344.4]
  wire  regs_104_reset; // @[RegFile.scala 66:20:@43344.4]
  wire [63:0] regs_104_io_in; // @[RegFile.scala 66:20:@43344.4]
  wire  regs_104_io_reset; // @[RegFile.scala 66:20:@43344.4]
  wire [63:0] regs_104_io_out; // @[RegFile.scala 66:20:@43344.4]
  wire  regs_104_io_enable; // @[RegFile.scala 66:20:@43344.4]
  wire  regs_105_clock; // @[RegFile.scala 66:20:@43358.4]
  wire  regs_105_reset; // @[RegFile.scala 66:20:@43358.4]
  wire [63:0] regs_105_io_in; // @[RegFile.scala 66:20:@43358.4]
  wire  regs_105_io_reset; // @[RegFile.scala 66:20:@43358.4]
  wire [63:0] regs_105_io_out; // @[RegFile.scala 66:20:@43358.4]
  wire  regs_105_io_enable; // @[RegFile.scala 66:20:@43358.4]
  wire  regs_106_clock; // @[RegFile.scala 66:20:@43372.4]
  wire  regs_106_reset; // @[RegFile.scala 66:20:@43372.4]
  wire [63:0] regs_106_io_in; // @[RegFile.scala 66:20:@43372.4]
  wire  regs_106_io_reset; // @[RegFile.scala 66:20:@43372.4]
  wire [63:0] regs_106_io_out; // @[RegFile.scala 66:20:@43372.4]
  wire  regs_106_io_enable; // @[RegFile.scala 66:20:@43372.4]
  wire  regs_107_clock; // @[RegFile.scala 66:20:@43386.4]
  wire  regs_107_reset; // @[RegFile.scala 66:20:@43386.4]
  wire [63:0] regs_107_io_in; // @[RegFile.scala 66:20:@43386.4]
  wire  regs_107_io_reset; // @[RegFile.scala 66:20:@43386.4]
  wire [63:0] regs_107_io_out; // @[RegFile.scala 66:20:@43386.4]
  wire  regs_107_io_enable; // @[RegFile.scala 66:20:@43386.4]
  wire  regs_108_clock; // @[RegFile.scala 66:20:@43400.4]
  wire  regs_108_reset; // @[RegFile.scala 66:20:@43400.4]
  wire [63:0] regs_108_io_in; // @[RegFile.scala 66:20:@43400.4]
  wire  regs_108_io_reset; // @[RegFile.scala 66:20:@43400.4]
  wire [63:0] regs_108_io_out; // @[RegFile.scala 66:20:@43400.4]
  wire  regs_108_io_enable; // @[RegFile.scala 66:20:@43400.4]
  wire  regs_109_clock; // @[RegFile.scala 66:20:@43414.4]
  wire  regs_109_reset; // @[RegFile.scala 66:20:@43414.4]
  wire [63:0] regs_109_io_in; // @[RegFile.scala 66:20:@43414.4]
  wire  regs_109_io_reset; // @[RegFile.scala 66:20:@43414.4]
  wire [63:0] regs_109_io_out; // @[RegFile.scala 66:20:@43414.4]
  wire  regs_109_io_enable; // @[RegFile.scala 66:20:@43414.4]
  wire  regs_110_clock; // @[RegFile.scala 66:20:@43428.4]
  wire  regs_110_reset; // @[RegFile.scala 66:20:@43428.4]
  wire [63:0] regs_110_io_in; // @[RegFile.scala 66:20:@43428.4]
  wire  regs_110_io_reset; // @[RegFile.scala 66:20:@43428.4]
  wire [63:0] regs_110_io_out; // @[RegFile.scala 66:20:@43428.4]
  wire  regs_110_io_enable; // @[RegFile.scala 66:20:@43428.4]
  wire  regs_111_clock; // @[RegFile.scala 66:20:@43442.4]
  wire  regs_111_reset; // @[RegFile.scala 66:20:@43442.4]
  wire [63:0] regs_111_io_in; // @[RegFile.scala 66:20:@43442.4]
  wire  regs_111_io_reset; // @[RegFile.scala 66:20:@43442.4]
  wire [63:0] regs_111_io_out; // @[RegFile.scala 66:20:@43442.4]
  wire  regs_111_io_enable; // @[RegFile.scala 66:20:@43442.4]
  wire  regs_112_clock; // @[RegFile.scala 66:20:@43456.4]
  wire  regs_112_reset; // @[RegFile.scala 66:20:@43456.4]
  wire [63:0] regs_112_io_in; // @[RegFile.scala 66:20:@43456.4]
  wire  regs_112_io_reset; // @[RegFile.scala 66:20:@43456.4]
  wire [63:0] regs_112_io_out; // @[RegFile.scala 66:20:@43456.4]
  wire  regs_112_io_enable; // @[RegFile.scala 66:20:@43456.4]
  wire  regs_113_clock; // @[RegFile.scala 66:20:@43470.4]
  wire  regs_113_reset; // @[RegFile.scala 66:20:@43470.4]
  wire [63:0] regs_113_io_in; // @[RegFile.scala 66:20:@43470.4]
  wire  regs_113_io_reset; // @[RegFile.scala 66:20:@43470.4]
  wire [63:0] regs_113_io_out; // @[RegFile.scala 66:20:@43470.4]
  wire  regs_113_io_enable; // @[RegFile.scala 66:20:@43470.4]
  wire  regs_114_clock; // @[RegFile.scala 66:20:@43484.4]
  wire  regs_114_reset; // @[RegFile.scala 66:20:@43484.4]
  wire [63:0] regs_114_io_in; // @[RegFile.scala 66:20:@43484.4]
  wire  regs_114_io_reset; // @[RegFile.scala 66:20:@43484.4]
  wire [63:0] regs_114_io_out; // @[RegFile.scala 66:20:@43484.4]
  wire  regs_114_io_enable; // @[RegFile.scala 66:20:@43484.4]
  wire  regs_115_clock; // @[RegFile.scala 66:20:@43498.4]
  wire  regs_115_reset; // @[RegFile.scala 66:20:@43498.4]
  wire [63:0] regs_115_io_in; // @[RegFile.scala 66:20:@43498.4]
  wire  regs_115_io_reset; // @[RegFile.scala 66:20:@43498.4]
  wire [63:0] regs_115_io_out; // @[RegFile.scala 66:20:@43498.4]
  wire  regs_115_io_enable; // @[RegFile.scala 66:20:@43498.4]
  wire  regs_116_clock; // @[RegFile.scala 66:20:@43512.4]
  wire  regs_116_reset; // @[RegFile.scala 66:20:@43512.4]
  wire [63:0] regs_116_io_in; // @[RegFile.scala 66:20:@43512.4]
  wire  regs_116_io_reset; // @[RegFile.scala 66:20:@43512.4]
  wire [63:0] regs_116_io_out; // @[RegFile.scala 66:20:@43512.4]
  wire  regs_116_io_enable; // @[RegFile.scala 66:20:@43512.4]
  wire  regs_117_clock; // @[RegFile.scala 66:20:@43526.4]
  wire  regs_117_reset; // @[RegFile.scala 66:20:@43526.4]
  wire [63:0] regs_117_io_in; // @[RegFile.scala 66:20:@43526.4]
  wire  regs_117_io_reset; // @[RegFile.scala 66:20:@43526.4]
  wire [63:0] regs_117_io_out; // @[RegFile.scala 66:20:@43526.4]
  wire  regs_117_io_enable; // @[RegFile.scala 66:20:@43526.4]
  wire  regs_118_clock; // @[RegFile.scala 66:20:@43540.4]
  wire  regs_118_reset; // @[RegFile.scala 66:20:@43540.4]
  wire [63:0] regs_118_io_in; // @[RegFile.scala 66:20:@43540.4]
  wire  regs_118_io_reset; // @[RegFile.scala 66:20:@43540.4]
  wire [63:0] regs_118_io_out; // @[RegFile.scala 66:20:@43540.4]
  wire  regs_118_io_enable; // @[RegFile.scala 66:20:@43540.4]
  wire  regs_119_clock; // @[RegFile.scala 66:20:@43554.4]
  wire  regs_119_reset; // @[RegFile.scala 66:20:@43554.4]
  wire [63:0] regs_119_io_in; // @[RegFile.scala 66:20:@43554.4]
  wire  regs_119_io_reset; // @[RegFile.scala 66:20:@43554.4]
  wire [63:0] regs_119_io_out; // @[RegFile.scala 66:20:@43554.4]
  wire  regs_119_io_enable; // @[RegFile.scala 66:20:@43554.4]
  wire  regs_120_clock; // @[RegFile.scala 66:20:@43568.4]
  wire  regs_120_reset; // @[RegFile.scala 66:20:@43568.4]
  wire [63:0] regs_120_io_in; // @[RegFile.scala 66:20:@43568.4]
  wire  regs_120_io_reset; // @[RegFile.scala 66:20:@43568.4]
  wire [63:0] regs_120_io_out; // @[RegFile.scala 66:20:@43568.4]
  wire  regs_120_io_enable; // @[RegFile.scala 66:20:@43568.4]
  wire  regs_121_clock; // @[RegFile.scala 66:20:@43582.4]
  wire  regs_121_reset; // @[RegFile.scala 66:20:@43582.4]
  wire [63:0] regs_121_io_in; // @[RegFile.scala 66:20:@43582.4]
  wire  regs_121_io_reset; // @[RegFile.scala 66:20:@43582.4]
  wire [63:0] regs_121_io_out; // @[RegFile.scala 66:20:@43582.4]
  wire  regs_121_io_enable; // @[RegFile.scala 66:20:@43582.4]
  wire  regs_122_clock; // @[RegFile.scala 66:20:@43596.4]
  wire  regs_122_reset; // @[RegFile.scala 66:20:@43596.4]
  wire [63:0] regs_122_io_in; // @[RegFile.scala 66:20:@43596.4]
  wire  regs_122_io_reset; // @[RegFile.scala 66:20:@43596.4]
  wire [63:0] regs_122_io_out; // @[RegFile.scala 66:20:@43596.4]
  wire  regs_122_io_enable; // @[RegFile.scala 66:20:@43596.4]
  wire  regs_123_clock; // @[RegFile.scala 66:20:@43610.4]
  wire  regs_123_reset; // @[RegFile.scala 66:20:@43610.4]
  wire [63:0] regs_123_io_in; // @[RegFile.scala 66:20:@43610.4]
  wire  regs_123_io_reset; // @[RegFile.scala 66:20:@43610.4]
  wire [63:0] regs_123_io_out; // @[RegFile.scala 66:20:@43610.4]
  wire  regs_123_io_enable; // @[RegFile.scala 66:20:@43610.4]
  wire  regs_124_clock; // @[RegFile.scala 66:20:@43624.4]
  wire  regs_124_reset; // @[RegFile.scala 66:20:@43624.4]
  wire [63:0] regs_124_io_in; // @[RegFile.scala 66:20:@43624.4]
  wire  regs_124_io_reset; // @[RegFile.scala 66:20:@43624.4]
  wire [63:0] regs_124_io_out; // @[RegFile.scala 66:20:@43624.4]
  wire  regs_124_io_enable; // @[RegFile.scala 66:20:@43624.4]
  wire  regs_125_clock; // @[RegFile.scala 66:20:@43638.4]
  wire  regs_125_reset; // @[RegFile.scala 66:20:@43638.4]
  wire [63:0] regs_125_io_in; // @[RegFile.scala 66:20:@43638.4]
  wire  regs_125_io_reset; // @[RegFile.scala 66:20:@43638.4]
  wire [63:0] regs_125_io_out; // @[RegFile.scala 66:20:@43638.4]
  wire  regs_125_io_enable; // @[RegFile.scala 66:20:@43638.4]
  wire  regs_126_clock; // @[RegFile.scala 66:20:@43652.4]
  wire  regs_126_reset; // @[RegFile.scala 66:20:@43652.4]
  wire [63:0] regs_126_io_in; // @[RegFile.scala 66:20:@43652.4]
  wire  regs_126_io_reset; // @[RegFile.scala 66:20:@43652.4]
  wire [63:0] regs_126_io_out; // @[RegFile.scala 66:20:@43652.4]
  wire  regs_126_io_enable; // @[RegFile.scala 66:20:@43652.4]
  wire  regs_127_clock; // @[RegFile.scala 66:20:@43666.4]
  wire  regs_127_reset; // @[RegFile.scala 66:20:@43666.4]
  wire [63:0] regs_127_io_in; // @[RegFile.scala 66:20:@43666.4]
  wire  regs_127_io_reset; // @[RegFile.scala 66:20:@43666.4]
  wire [63:0] regs_127_io_out; // @[RegFile.scala 66:20:@43666.4]
  wire  regs_127_io_enable; // @[RegFile.scala 66:20:@43666.4]
  wire  regs_128_clock; // @[RegFile.scala 66:20:@43680.4]
  wire  regs_128_reset; // @[RegFile.scala 66:20:@43680.4]
  wire [63:0] regs_128_io_in; // @[RegFile.scala 66:20:@43680.4]
  wire  regs_128_io_reset; // @[RegFile.scala 66:20:@43680.4]
  wire [63:0] regs_128_io_out; // @[RegFile.scala 66:20:@43680.4]
  wire  regs_128_io_enable; // @[RegFile.scala 66:20:@43680.4]
  wire  regs_129_clock; // @[RegFile.scala 66:20:@43694.4]
  wire  regs_129_reset; // @[RegFile.scala 66:20:@43694.4]
  wire [63:0] regs_129_io_in; // @[RegFile.scala 66:20:@43694.4]
  wire  regs_129_io_reset; // @[RegFile.scala 66:20:@43694.4]
  wire [63:0] regs_129_io_out; // @[RegFile.scala 66:20:@43694.4]
  wire  regs_129_io_enable; // @[RegFile.scala 66:20:@43694.4]
  wire  regs_130_clock; // @[RegFile.scala 66:20:@43708.4]
  wire  regs_130_reset; // @[RegFile.scala 66:20:@43708.4]
  wire [63:0] regs_130_io_in; // @[RegFile.scala 66:20:@43708.4]
  wire  regs_130_io_reset; // @[RegFile.scala 66:20:@43708.4]
  wire [63:0] regs_130_io_out; // @[RegFile.scala 66:20:@43708.4]
  wire  regs_130_io_enable; // @[RegFile.scala 66:20:@43708.4]
  wire  regs_131_clock; // @[RegFile.scala 66:20:@43722.4]
  wire  regs_131_reset; // @[RegFile.scala 66:20:@43722.4]
  wire [63:0] regs_131_io_in; // @[RegFile.scala 66:20:@43722.4]
  wire  regs_131_io_reset; // @[RegFile.scala 66:20:@43722.4]
  wire [63:0] regs_131_io_out; // @[RegFile.scala 66:20:@43722.4]
  wire  regs_131_io_enable; // @[RegFile.scala 66:20:@43722.4]
  wire  regs_132_clock; // @[RegFile.scala 66:20:@43736.4]
  wire  regs_132_reset; // @[RegFile.scala 66:20:@43736.4]
  wire [63:0] regs_132_io_in; // @[RegFile.scala 66:20:@43736.4]
  wire  regs_132_io_reset; // @[RegFile.scala 66:20:@43736.4]
  wire [63:0] regs_132_io_out; // @[RegFile.scala 66:20:@43736.4]
  wire  regs_132_io_enable; // @[RegFile.scala 66:20:@43736.4]
  wire  regs_133_clock; // @[RegFile.scala 66:20:@43750.4]
  wire  regs_133_reset; // @[RegFile.scala 66:20:@43750.4]
  wire [63:0] regs_133_io_in; // @[RegFile.scala 66:20:@43750.4]
  wire  regs_133_io_reset; // @[RegFile.scala 66:20:@43750.4]
  wire [63:0] regs_133_io_out; // @[RegFile.scala 66:20:@43750.4]
  wire  regs_133_io_enable; // @[RegFile.scala 66:20:@43750.4]
  wire  regs_134_clock; // @[RegFile.scala 66:20:@43764.4]
  wire  regs_134_reset; // @[RegFile.scala 66:20:@43764.4]
  wire [63:0] regs_134_io_in; // @[RegFile.scala 66:20:@43764.4]
  wire  regs_134_io_reset; // @[RegFile.scala 66:20:@43764.4]
  wire [63:0] regs_134_io_out; // @[RegFile.scala 66:20:@43764.4]
  wire  regs_134_io_enable; // @[RegFile.scala 66:20:@43764.4]
  wire  regs_135_clock; // @[RegFile.scala 66:20:@43778.4]
  wire  regs_135_reset; // @[RegFile.scala 66:20:@43778.4]
  wire [63:0] regs_135_io_in; // @[RegFile.scala 66:20:@43778.4]
  wire  regs_135_io_reset; // @[RegFile.scala 66:20:@43778.4]
  wire [63:0] regs_135_io_out; // @[RegFile.scala 66:20:@43778.4]
  wire  regs_135_io_enable; // @[RegFile.scala 66:20:@43778.4]
  wire  regs_136_clock; // @[RegFile.scala 66:20:@43792.4]
  wire  regs_136_reset; // @[RegFile.scala 66:20:@43792.4]
  wire [63:0] regs_136_io_in; // @[RegFile.scala 66:20:@43792.4]
  wire  regs_136_io_reset; // @[RegFile.scala 66:20:@43792.4]
  wire [63:0] regs_136_io_out; // @[RegFile.scala 66:20:@43792.4]
  wire  regs_136_io_enable; // @[RegFile.scala 66:20:@43792.4]
  wire  regs_137_clock; // @[RegFile.scala 66:20:@43806.4]
  wire  regs_137_reset; // @[RegFile.scala 66:20:@43806.4]
  wire [63:0] regs_137_io_in; // @[RegFile.scala 66:20:@43806.4]
  wire  regs_137_io_reset; // @[RegFile.scala 66:20:@43806.4]
  wire [63:0] regs_137_io_out; // @[RegFile.scala 66:20:@43806.4]
  wire  regs_137_io_enable; // @[RegFile.scala 66:20:@43806.4]
  wire  regs_138_clock; // @[RegFile.scala 66:20:@43820.4]
  wire  regs_138_reset; // @[RegFile.scala 66:20:@43820.4]
  wire [63:0] regs_138_io_in; // @[RegFile.scala 66:20:@43820.4]
  wire  regs_138_io_reset; // @[RegFile.scala 66:20:@43820.4]
  wire [63:0] regs_138_io_out; // @[RegFile.scala 66:20:@43820.4]
  wire  regs_138_io_enable; // @[RegFile.scala 66:20:@43820.4]
  wire  regs_139_clock; // @[RegFile.scala 66:20:@43834.4]
  wire  regs_139_reset; // @[RegFile.scala 66:20:@43834.4]
  wire [63:0] regs_139_io_in; // @[RegFile.scala 66:20:@43834.4]
  wire  regs_139_io_reset; // @[RegFile.scala 66:20:@43834.4]
  wire [63:0] regs_139_io_out; // @[RegFile.scala 66:20:@43834.4]
  wire  regs_139_io_enable; // @[RegFile.scala 66:20:@43834.4]
  wire  regs_140_clock; // @[RegFile.scala 66:20:@43848.4]
  wire  regs_140_reset; // @[RegFile.scala 66:20:@43848.4]
  wire [63:0] regs_140_io_in; // @[RegFile.scala 66:20:@43848.4]
  wire  regs_140_io_reset; // @[RegFile.scala 66:20:@43848.4]
  wire [63:0] regs_140_io_out; // @[RegFile.scala 66:20:@43848.4]
  wire  regs_140_io_enable; // @[RegFile.scala 66:20:@43848.4]
  wire  regs_141_clock; // @[RegFile.scala 66:20:@43862.4]
  wire  regs_141_reset; // @[RegFile.scala 66:20:@43862.4]
  wire [63:0] regs_141_io_in; // @[RegFile.scala 66:20:@43862.4]
  wire  regs_141_io_reset; // @[RegFile.scala 66:20:@43862.4]
  wire [63:0] regs_141_io_out; // @[RegFile.scala 66:20:@43862.4]
  wire  regs_141_io_enable; // @[RegFile.scala 66:20:@43862.4]
  wire  regs_142_clock; // @[RegFile.scala 66:20:@43876.4]
  wire  regs_142_reset; // @[RegFile.scala 66:20:@43876.4]
  wire [63:0] regs_142_io_in; // @[RegFile.scala 66:20:@43876.4]
  wire  regs_142_io_reset; // @[RegFile.scala 66:20:@43876.4]
  wire [63:0] regs_142_io_out; // @[RegFile.scala 66:20:@43876.4]
  wire  regs_142_io_enable; // @[RegFile.scala 66:20:@43876.4]
  wire  regs_143_clock; // @[RegFile.scala 66:20:@43890.4]
  wire  regs_143_reset; // @[RegFile.scala 66:20:@43890.4]
  wire [63:0] regs_143_io_in; // @[RegFile.scala 66:20:@43890.4]
  wire  regs_143_io_reset; // @[RegFile.scala 66:20:@43890.4]
  wire [63:0] regs_143_io_out; // @[RegFile.scala 66:20:@43890.4]
  wire  regs_143_io_enable; // @[RegFile.scala 66:20:@43890.4]
  wire  regs_144_clock; // @[RegFile.scala 66:20:@43904.4]
  wire  regs_144_reset; // @[RegFile.scala 66:20:@43904.4]
  wire [63:0] regs_144_io_in; // @[RegFile.scala 66:20:@43904.4]
  wire  regs_144_io_reset; // @[RegFile.scala 66:20:@43904.4]
  wire [63:0] regs_144_io_out; // @[RegFile.scala 66:20:@43904.4]
  wire  regs_144_io_enable; // @[RegFile.scala 66:20:@43904.4]
  wire  regs_145_clock; // @[RegFile.scala 66:20:@43918.4]
  wire  regs_145_reset; // @[RegFile.scala 66:20:@43918.4]
  wire [63:0] regs_145_io_in; // @[RegFile.scala 66:20:@43918.4]
  wire  regs_145_io_reset; // @[RegFile.scala 66:20:@43918.4]
  wire [63:0] regs_145_io_out; // @[RegFile.scala 66:20:@43918.4]
  wire  regs_145_io_enable; // @[RegFile.scala 66:20:@43918.4]
  wire  regs_146_clock; // @[RegFile.scala 66:20:@43932.4]
  wire  regs_146_reset; // @[RegFile.scala 66:20:@43932.4]
  wire [63:0] regs_146_io_in; // @[RegFile.scala 66:20:@43932.4]
  wire  regs_146_io_reset; // @[RegFile.scala 66:20:@43932.4]
  wire [63:0] regs_146_io_out; // @[RegFile.scala 66:20:@43932.4]
  wire  regs_146_io_enable; // @[RegFile.scala 66:20:@43932.4]
  wire  regs_147_clock; // @[RegFile.scala 66:20:@43946.4]
  wire  regs_147_reset; // @[RegFile.scala 66:20:@43946.4]
  wire [63:0] regs_147_io_in; // @[RegFile.scala 66:20:@43946.4]
  wire  regs_147_io_reset; // @[RegFile.scala 66:20:@43946.4]
  wire [63:0] regs_147_io_out; // @[RegFile.scala 66:20:@43946.4]
  wire  regs_147_io_enable; // @[RegFile.scala 66:20:@43946.4]
  wire  regs_148_clock; // @[RegFile.scala 66:20:@43960.4]
  wire  regs_148_reset; // @[RegFile.scala 66:20:@43960.4]
  wire [63:0] regs_148_io_in; // @[RegFile.scala 66:20:@43960.4]
  wire  regs_148_io_reset; // @[RegFile.scala 66:20:@43960.4]
  wire [63:0] regs_148_io_out; // @[RegFile.scala 66:20:@43960.4]
  wire  regs_148_io_enable; // @[RegFile.scala 66:20:@43960.4]
  wire  regs_149_clock; // @[RegFile.scala 66:20:@43974.4]
  wire  regs_149_reset; // @[RegFile.scala 66:20:@43974.4]
  wire [63:0] regs_149_io_in; // @[RegFile.scala 66:20:@43974.4]
  wire  regs_149_io_reset; // @[RegFile.scala 66:20:@43974.4]
  wire [63:0] regs_149_io_out; // @[RegFile.scala 66:20:@43974.4]
  wire  regs_149_io_enable; // @[RegFile.scala 66:20:@43974.4]
  wire  regs_150_clock; // @[RegFile.scala 66:20:@43988.4]
  wire  regs_150_reset; // @[RegFile.scala 66:20:@43988.4]
  wire [63:0] regs_150_io_in; // @[RegFile.scala 66:20:@43988.4]
  wire  regs_150_io_reset; // @[RegFile.scala 66:20:@43988.4]
  wire [63:0] regs_150_io_out; // @[RegFile.scala 66:20:@43988.4]
  wire  regs_150_io_enable; // @[RegFile.scala 66:20:@43988.4]
  wire  regs_151_clock; // @[RegFile.scala 66:20:@44002.4]
  wire  regs_151_reset; // @[RegFile.scala 66:20:@44002.4]
  wire [63:0] regs_151_io_in; // @[RegFile.scala 66:20:@44002.4]
  wire  regs_151_io_reset; // @[RegFile.scala 66:20:@44002.4]
  wire [63:0] regs_151_io_out; // @[RegFile.scala 66:20:@44002.4]
  wire  regs_151_io_enable; // @[RegFile.scala 66:20:@44002.4]
  wire  regs_152_clock; // @[RegFile.scala 66:20:@44016.4]
  wire  regs_152_reset; // @[RegFile.scala 66:20:@44016.4]
  wire [63:0] regs_152_io_in; // @[RegFile.scala 66:20:@44016.4]
  wire  regs_152_io_reset; // @[RegFile.scala 66:20:@44016.4]
  wire [63:0] regs_152_io_out; // @[RegFile.scala 66:20:@44016.4]
  wire  regs_152_io_enable; // @[RegFile.scala 66:20:@44016.4]
  wire  regs_153_clock; // @[RegFile.scala 66:20:@44030.4]
  wire  regs_153_reset; // @[RegFile.scala 66:20:@44030.4]
  wire [63:0] regs_153_io_in; // @[RegFile.scala 66:20:@44030.4]
  wire  regs_153_io_reset; // @[RegFile.scala 66:20:@44030.4]
  wire [63:0] regs_153_io_out; // @[RegFile.scala 66:20:@44030.4]
  wire  regs_153_io_enable; // @[RegFile.scala 66:20:@44030.4]
  wire  regs_154_clock; // @[RegFile.scala 66:20:@44044.4]
  wire  regs_154_reset; // @[RegFile.scala 66:20:@44044.4]
  wire [63:0] regs_154_io_in; // @[RegFile.scala 66:20:@44044.4]
  wire  regs_154_io_reset; // @[RegFile.scala 66:20:@44044.4]
  wire [63:0] regs_154_io_out; // @[RegFile.scala 66:20:@44044.4]
  wire  regs_154_io_enable; // @[RegFile.scala 66:20:@44044.4]
  wire  regs_155_clock; // @[RegFile.scala 66:20:@44058.4]
  wire  regs_155_reset; // @[RegFile.scala 66:20:@44058.4]
  wire [63:0] regs_155_io_in; // @[RegFile.scala 66:20:@44058.4]
  wire  regs_155_io_reset; // @[RegFile.scala 66:20:@44058.4]
  wire [63:0] regs_155_io_out; // @[RegFile.scala 66:20:@44058.4]
  wire  regs_155_io_enable; // @[RegFile.scala 66:20:@44058.4]
  wire  regs_156_clock; // @[RegFile.scala 66:20:@44072.4]
  wire  regs_156_reset; // @[RegFile.scala 66:20:@44072.4]
  wire [63:0] regs_156_io_in; // @[RegFile.scala 66:20:@44072.4]
  wire  regs_156_io_reset; // @[RegFile.scala 66:20:@44072.4]
  wire [63:0] regs_156_io_out; // @[RegFile.scala 66:20:@44072.4]
  wire  regs_156_io_enable; // @[RegFile.scala 66:20:@44072.4]
  wire  regs_157_clock; // @[RegFile.scala 66:20:@44086.4]
  wire  regs_157_reset; // @[RegFile.scala 66:20:@44086.4]
  wire [63:0] regs_157_io_in; // @[RegFile.scala 66:20:@44086.4]
  wire  regs_157_io_reset; // @[RegFile.scala 66:20:@44086.4]
  wire [63:0] regs_157_io_out; // @[RegFile.scala 66:20:@44086.4]
  wire  regs_157_io_enable; // @[RegFile.scala 66:20:@44086.4]
  wire  regs_158_clock; // @[RegFile.scala 66:20:@44100.4]
  wire  regs_158_reset; // @[RegFile.scala 66:20:@44100.4]
  wire [63:0] regs_158_io_in; // @[RegFile.scala 66:20:@44100.4]
  wire  regs_158_io_reset; // @[RegFile.scala 66:20:@44100.4]
  wire [63:0] regs_158_io_out; // @[RegFile.scala 66:20:@44100.4]
  wire  regs_158_io_enable; // @[RegFile.scala 66:20:@44100.4]
  wire  regs_159_clock; // @[RegFile.scala 66:20:@44114.4]
  wire  regs_159_reset; // @[RegFile.scala 66:20:@44114.4]
  wire [63:0] regs_159_io_in; // @[RegFile.scala 66:20:@44114.4]
  wire  regs_159_io_reset; // @[RegFile.scala 66:20:@44114.4]
  wire [63:0] regs_159_io_out; // @[RegFile.scala 66:20:@44114.4]
  wire  regs_159_io_enable; // @[RegFile.scala 66:20:@44114.4]
  wire  regs_160_clock; // @[RegFile.scala 66:20:@44128.4]
  wire  regs_160_reset; // @[RegFile.scala 66:20:@44128.4]
  wire [63:0] regs_160_io_in; // @[RegFile.scala 66:20:@44128.4]
  wire  regs_160_io_reset; // @[RegFile.scala 66:20:@44128.4]
  wire [63:0] regs_160_io_out; // @[RegFile.scala 66:20:@44128.4]
  wire  regs_160_io_enable; // @[RegFile.scala 66:20:@44128.4]
  wire  regs_161_clock; // @[RegFile.scala 66:20:@44142.4]
  wire  regs_161_reset; // @[RegFile.scala 66:20:@44142.4]
  wire [63:0] regs_161_io_in; // @[RegFile.scala 66:20:@44142.4]
  wire  regs_161_io_reset; // @[RegFile.scala 66:20:@44142.4]
  wire [63:0] regs_161_io_out; // @[RegFile.scala 66:20:@44142.4]
  wire  regs_161_io_enable; // @[RegFile.scala 66:20:@44142.4]
  wire  regs_162_clock; // @[RegFile.scala 66:20:@44156.4]
  wire  regs_162_reset; // @[RegFile.scala 66:20:@44156.4]
  wire [63:0] regs_162_io_in; // @[RegFile.scala 66:20:@44156.4]
  wire  regs_162_io_reset; // @[RegFile.scala 66:20:@44156.4]
  wire [63:0] regs_162_io_out; // @[RegFile.scala 66:20:@44156.4]
  wire  regs_162_io_enable; // @[RegFile.scala 66:20:@44156.4]
  wire  regs_163_clock; // @[RegFile.scala 66:20:@44170.4]
  wire  regs_163_reset; // @[RegFile.scala 66:20:@44170.4]
  wire [63:0] regs_163_io_in; // @[RegFile.scala 66:20:@44170.4]
  wire  regs_163_io_reset; // @[RegFile.scala 66:20:@44170.4]
  wire [63:0] regs_163_io_out; // @[RegFile.scala 66:20:@44170.4]
  wire  regs_163_io_enable; // @[RegFile.scala 66:20:@44170.4]
  wire  regs_164_clock; // @[RegFile.scala 66:20:@44184.4]
  wire  regs_164_reset; // @[RegFile.scala 66:20:@44184.4]
  wire [63:0] regs_164_io_in; // @[RegFile.scala 66:20:@44184.4]
  wire  regs_164_io_reset; // @[RegFile.scala 66:20:@44184.4]
  wire [63:0] regs_164_io_out; // @[RegFile.scala 66:20:@44184.4]
  wire  regs_164_io_enable; // @[RegFile.scala 66:20:@44184.4]
  wire  regs_165_clock; // @[RegFile.scala 66:20:@44198.4]
  wire  regs_165_reset; // @[RegFile.scala 66:20:@44198.4]
  wire [63:0] regs_165_io_in; // @[RegFile.scala 66:20:@44198.4]
  wire  regs_165_io_reset; // @[RegFile.scala 66:20:@44198.4]
  wire [63:0] regs_165_io_out; // @[RegFile.scala 66:20:@44198.4]
  wire  regs_165_io_enable; // @[RegFile.scala 66:20:@44198.4]
  wire  regs_166_clock; // @[RegFile.scala 66:20:@44212.4]
  wire  regs_166_reset; // @[RegFile.scala 66:20:@44212.4]
  wire [63:0] regs_166_io_in; // @[RegFile.scala 66:20:@44212.4]
  wire  regs_166_io_reset; // @[RegFile.scala 66:20:@44212.4]
  wire [63:0] regs_166_io_out; // @[RegFile.scala 66:20:@44212.4]
  wire  regs_166_io_enable; // @[RegFile.scala 66:20:@44212.4]
  wire  regs_167_clock; // @[RegFile.scala 66:20:@44226.4]
  wire  regs_167_reset; // @[RegFile.scala 66:20:@44226.4]
  wire [63:0] regs_167_io_in; // @[RegFile.scala 66:20:@44226.4]
  wire  regs_167_io_reset; // @[RegFile.scala 66:20:@44226.4]
  wire [63:0] regs_167_io_out; // @[RegFile.scala 66:20:@44226.4]
  wire  regs_167_io_enable; // @[RegFile.scala 66:20:@44226.4]
  wire  regs_168_clock; // @[RegFile.scala 66:20:@44240.4]
  wire  regs_168_reset; // @[RegFile.scala 66:20:@44240.4]
  wire [63:0] regs_168_io_in; // @[RegFile.scala 66:20:@44240.4]
  wire  regs_168_io_reset; // @[RegFile.scala 66:20:@44240.4]
  wire [63:0] regs_168_io_out; // @[RegFile.scala 66:20:@44240.4]
  wire  regs_168_io_enable; // @[RegFile.scala 66:20:@44240.4]
  wire  regs_169_clock; // @[RegFile.scala 66:20:@44254.4]
  wire  regs_169_reset; // @[RegFile.scala 66:20:@44254.4]
  wire [63:0] regs_169_io_in; // @[RegFile.scala 66:20:@44254.4]
  wire  regs_169_io_reset; // @[RegFile.scala 66:20:@44254.4]
  wire [63:0] regs_169_io_out; // @[RegFile.scala 66:20:@44254.4]
  wire  regs_169_io_enable; // @[RegFile.scala 66:20:@44254.4]
  wire  regs_170_clock; // @[RegFile.scala 66:20:@44268.4]
  wire  regs_170_reset; // @[RegFile.scala 66:20:@44268.4]
  wire [63:0] regs_170_io_in; // @[RegFile.scala 66:20:@44268.4]
  wire  regs_170_io_reset; // @[RegFile.scala 66:20:@44268.4]
  wire [63:0] regs_170_io_out; // @[RegFile.scala 66:20:@44268.4]
  wire  regs_170_io_enable; // @[RegFile.scala 66:20:@44268.4]
  wire  regs_171_clock; // @[RegFile.scala 66:20:@44282.4]
  wire  regs_171_reset; // @[RegFile.scala 66:20:@44282.4]
  wire [63:0] regs_171_io_in; // @[RegFile.scala 66:20:@44282.4]
  wire  regs_171_io_reset; // @[RegFile.scala 66:20:@44282.4]
  wire [63:0] regs_171_io_out; // @[RegFile.scala 66:20:@44282.4]
  wire  regs_171_io_enable; // @[RegFile.scala 66:20:@44282.4]
  wire  regs_172_clock; // @[RegFile.scala 66:20:@44296.4]
  wire  regs_172_reset; // @[RegFile.scala 66:20:@44296.4]
  wire [63:0] regs_172_io_in; // @[RegFile.scala 66:20:@44296.4]
  wire  regs_172_io_reset; // @[RegFile.scala 66:20:@44296.4]
  wire [63:0] regs_172_io_out; // @[RegFile.scala 66:20:@44296.4]
  wire  regs_172_io_enable; // @[RegFile.scala 66:20:@44296.4]
  wire  regs_173_clock; // @[RegFile.scala 66:20:@44310.4]
  wire  regs_173_reset; // @[RegFile.scala 66:20:@44310.4]
  wire [63:0] regs_173_io_in; // @[RegFile.scala 66:20:@44310.4]
  wire  regs_173_io_reset; // @[RegFile.scala 66:20:@44310.4]
  wire [63:0] regs_173_io_out; // @[RegFile.scala 66:20:@44310.4]
  wire  regs_173_io_enable; // @[RegFile.scala 66:20:@44310.4]
  wire  regs_174_clock; // @[RegFile.scala 66:20:@44324.4]
  wire  regs_174_reset; // @[RegFile.scala 66:20:@44324.4]
  wire [63:0] regs_174_io_in; // @[RegFile.scala 66:20:@44324.4]
  wire  regs_174_io_reset; // @[RegFile.scala 66:20:@44324.4]
  wire [63:0] regs_174_io_out; // @[RegFile.scala 66:20:@44324.4]
  wire  regs_174_io_enable; // @[RegFile.scala 66:20:@44324.4]
  wire  regs_175_clock; // @[RegFile.scala 66:20:@44338.4]
  wire  regs_175_reset; // @[RegFile.scala 66:20:@44338.4]
  wire [63:0] regs_175_io_in; // @[RegFile.scala 66:20:@44338.4]
  wire  regs_175_io_reset; // @[RegFile.scala 66:20:@44338.4]
  wire [63:0] regs_175_io_out; // @[RegFile.scala 66:20:@44338.4]
  wire  regs_175_io_enable; // @[RegFile.scala 66:20:@44338.4]
  wire  regs_176_clock; // @[RegFile.scala 66:20:@44352.4]
  wire  regs_176_reset; // @[RegFile.scala 66:20:@44352.4]
  wire [63:0] regs_176_io_in; // @[RegFile.scala 66:20:@44352.4]
  wire  regs_176_io_reset; // @[RegFile.scala 66:20:@44352.4]
  wire [63:0] regs_176_io_out; // @[RegFile.scala 66:20:@44352.4]
  wire  regs_176_io_enable; // @[RegFile.scala 66:20:@44352.4]
  wire  regs_177_clock; // @[RegFile.scala 66:20:@44366.4]
  wire  regs_177_reset; // @[RegFile.scala 66:20:@44366.4]
  wire [63:0] regs_177_io_in; // @[RegFile.scala 66:20:@44366.4]
  wire  regs_177_io_reset; // @[RegFile.scala 66:20:@44366.4]
  wire [63:0] regs_177_io_out; // @[RegFile.scala 66:20:@44366.4]
  wire  regs_177_io_enable; // @[RegFile.scala 66:20:@44366.4]
  wire  regs_178_clock; // @[RegFile.scala 66:20:@44380.4]
  wire  regs_178_reset; // @[RegFile.scala 66:20:@44380.4]
  wire [63:0] regs_178_io_in; // @[RegFile.scala 66:20:@44380.4]
  wire  regs_178_io_reset; // @[RegFile.scala 66:20:@44380.4]
  wire [63:0] regs_178_io_out; // @[RegFile.scala 66:20:@44380.4]
  wire  regs_178_io_enable; // @[RegFile.scala 66:20:@44380.4]
  wire  regs_179_clock; // @[RegFile.scala 66:20:@44394.4]
  wire  regs_179_reset; // @[RegFile.scala 66:20:@44394.4]
  wire [63:0] regs_179_io_in; // @[RegFile.scala 66:20:@44394.4]
  wire  regs_179_io_reset; // @[RegFile.scala 66:20:@44394.4]
  wire [63:0] regs_179_io_out; // @[RegFile.scala 66:20:@44394.4]
  wire  regs_179_io_enable; // @[RegFile.scala 66:20:@44394.4]
  wire  regs_180_clock; // @[RegFile.scala 66:20:@44408.4]
  wire  regs_180_reset; // @[RegFile.scala 66:20:@44408.4]
  wire [63:0] regs_180_io_in; // @[RegFile.scala 66:20:@44408.4]
  wire  regs_180_io_reset; // @[RegFile.scala 66:20:@44408.4]
  wire [63:0] regs_180_io_out; // @[RegFile.scala 66:20:@44408.4]
  wire  regs_180_io_enable; // @[RegFile.scala 66:20:@44408.4]
  wire  regs_181_clock; // @[RegFile.scala 66:20:@44422.4]
  wire  regs_181_reset; // @[RegFile.scala 66:20:@44422.4]
  wire [63:0] regs_181_io_in; // @[RegFile.scala 66:20:@44422.4]
  wire  regs_181_io_reset; // @[RegFile.scala 66:20:@44422.4]
  wire [63:0] regs_181_io_out; // @[RegFile.scala 66:20:@44422.4]
  wire  regs_181_io_enable; // @[RegFile.scala 66:20:@44422.4]
  wire  regs_182_clock; // @[RegFile.scala 66:20:@44436.4]
  wire  regs_182_reset; // @[RegFile.scala 66:20:@44436.4]
  wire [63:0] regs_182_io_in; // @[RegFile.scala 66:20:@44436.4]
  wire  regs_182_io_reset; // @[RegFile.scala 66:20:@44436.4]
  wire [63:0] regs_182_io_out; // @[RegFile.scala 66:20:@44436.4]
  wire  regs_182_io_enable; // @[RegFile.scala 66:20:@44436.4]
  wire  regs_183_clock; // @[RegFile.scala 66:20:@44450.4]
  wire  regs_183_reset; // @[RegFile.scala 66:20:@44450.4]
  wire [63:0] regs_183_io_in; // @[RegFile.scala 66:20:@44450.4]
  wire  regs_183_io_reset; // @[RegFile.scala 66:20:@44450.4]
  wire [63:0] regs_183_io_out; // @[RegFile.scala 66:20:@44450.4]
  wire  regs_183_io_enable; // @[RegFile.scala 66:20:@44450.4]
  wire  regs_184_clock; // @[RegFile.scala 66:20:@44464.4]
  wire  regs_184_reset; // @[RegFile.scala 66:20:@44464.4]
  wire [63:0] regs_184_io_in; // @[RegFile.scala 66:20:@44464.4]
  wire  regs_184_io_reset; // @[RegFile.scala 66:20:@44464.4]
  wire [63:0] regs_184_io_out; // @[RegFile.scala 66:20:@44464.4]
  wire  regs_184_io_enable; // @[RegFile.scala 66:20:@44464.4]
  wire  regs_185_clock; // @[RegFile.scala 66:20:@44478.4]
  wire  regs_185_reset; // @[RegFile.scala 66:20:@44478.4]
  wire [63:0] regs_185_io_in; // @[RegFile.scala 66:20:@44478.4]
  wire  regs_185_io_reset; // @[RegFile.scala 66:20:@44478.4]
  wire [63:0] regs_185_io_out; // @[RegFile.scala 66:20:@44478.4]
  wire  regs_185_io_enable; // @[RegFile.scala 66:20:@44478.4]
  wire  regs_186_clock; // @[RegFile.scala 66:20:@44492.4]
  wire  regs_186_reset; // @[RegFile.scala 66:20:@44492.4]
  wire [63:0] regs_186_io_in; // @[RegFile.scala 66:20:@44492.4]
  wire  regs_186_io_reset; // @[RegFile.scala 66:20:@44492.4]
  wire [63:0] regs_186_io_out; // @[RegFile.scala 66:20:@44492.4]
  wire  regs_186_io_enable; // @[RegFile.scala 66:20:@44492.4]
  wire  regs_187_clock; // @[RegFile.scala 66:20:@44506.4]
  wire  regs_187_reset; // @[RegFile.scala 66:20:@44506.4]
  wire [63:0] regs_187_io_in; // @[RegFile.scala 66:20:@44506.4]
  wire  regs_187_io_reset; // @[RegFile.scala 66:20:@44506.4]
  wire [63:0] regs_187_io_out; // @[RegFile.scala 66:20:@44506.4]
  wire  regs_187_io_enable; // @[RegFile.scala 66:20:@44506.4]
  wire  regs_188_clock; // @[RegFile.scala 66:20:@44520.4]
  wire  regs_188_reset; // @[RegFile.scala 66:20:@44520.4]
  wire [63:0] regs_188_io_in; // @[RegFile.scala 66:20:@44520.4]
  wire  regs_188_io_reset; // @[RegFile.scala 66:20:@44520.4]
  wire [63:0] regs_188_io_out; // @[RegFile.scala 66:20:@44520.4]
  wire  regs_188_io_enable; // @[RegFile.scala 66:20:@44520.4]
  wire  regs_189_clock; // @[RegFile.scala 66:20:@44534.4]
  wire  regs_189_reset; // @[RegFile.scala 66:20:@44534.4]
  wire [63:0] regs_189_io_in; // @[RegFile.scala 66:20:@44534.4]
  wire  regs_189_io_reset; // @[RegFile.scala 66:20:@44534.4]
  wire [63:0] regs_189_io_out; // @[RegFile.scala 66:20:@44534.4]
  wire  regs_189_io_enable; // @[RegFile.scala 66:20:@44534.4]
  wire  regs_190_clock; // @[RegFile.scala 66:20:@44548.4]
  wire  regs_190_reset; // @[RegFile.scala 66:20:@44548.4]
  wire [63:0] regs_190_io_in; // @[RegFile.scala 66:20:@44548.4]
  wire  regs_190_io_reset; // @[RegFile.scala 66:20:@44548.4]
  wire [63:0] regs_190_io_out; // @[RegFile.scala 66:20:@44548.4]
  wire  regs_190_io_enable; // @[RegFile.scala 66:20:@44548.4]
  wire  regs_191_clock; // @[RegFile.scala 66:20:@44562.4]
  wire  regs_191_reset; // @[RegFile.scala 66:20:@44562.4]
  wire [63:0] regs_191_io_in; // @[RegFile.scala 66:20:@44562.4]
  wire  regs_191_io_reset; // @[RegFile.scala 66:20:@44562.4]
  wire [63:0] regs_191_io_out; // @[RegFile.scala 66:20:@44562.4]
  wire  regs_191_io_enable; // @[RegFile.scala 66:20:@44562.4]
  wire  regs_192_clock; // @[RegFile.scala 66:20:@44576.4]
  wire  regs_192_reset; // @[RegFile.scala 66:20:@44576.4]
  wire [63:0] regs_192_io_in; // @[RegFile.scala 66:20:@44576.4]
  wire  regs_192_io_reset; // @[RegFile.scala 66:20:@44576.4]
  wire [63:0] regs_192_io_out; // @[RegFile.scala 66:20:@44576.4]
  wire  regs_192_io_enable; // @[RegFile.scala 66:20:@44576.4]
  wire  regs_193_clock; // @[RegFile.scala 66:20:@44590.4]
  wire  regs_193_reset; // @[RegFile.scala 66:20:@44590.4]
  wire [63:0] regs_193_io_in; // @[RegFile.scala 66:20:@44590.4]
  wire  regs_193_io_reset; // @[RegFile.scala 66:20:@44590.4]
  wire [63:0] regs_193_io_out; // @[RegFile.scala 66:20:@44590.4]
  wire  regs_193_io_enable; // @[RegFile.scala 66:20:@44590.4]
  wire  regs_194_clock; // @[RegFile.scala 66:20:@44604.4]
  wire  regs_194_reset; // @[RegFile.scala 66:20:@44604.4]
  wire [63:0] regs_194_io_in; // @[RegFile.scala 66:20:@44604.4]
  wire  regs_194_io_reset; // @[RegFile.scala 66:20:@44604.4]
  wire [63:0] regs_194_io_out; // @[RegFile.scala 66:20:@44604.4]
  wire  regs_194_io_enable; // @[RegFile.scala 66:20:@44604.4]
  wire  regs_195_clock; // @[RegFile.scala 66:20:@44618.4]
  wire  regs_195_reset; // @[RegFile.scala 66:20:@44618.4]
  wire [63:0] regs_195_io_in; // @[RegFile.scala 66:20:@44618.4]
  wire  regs_195_io_reset; // @[RegFile.scala 66:20:@44618.4]
  wire [63:0] regs_195_io_out; // @[RegFile.scala 66:20:@44618.4]
  wire  regs_195_io_enable; // @[RegFile.scala 66:20:@44618.4]
  wire  regs_196_clock; // @[RegFile.scala 66:20:@44632.4]
  wire  regs_196_reset; // @[RegFile.scala 66:20:@44632.4]
  wire [63:0] regs_196_io_in; // @[RegFile.scala 66:20:@44632.4]
  wire  regs_196_io_reset; // @[RegFile.scala 66:20:@44632.4]
  wire [63:0] regs_196_io_out; // @[RegFile.scala 66:20:@44632.4]
  wire  regs_196_io_enable; // @[RegFile.scala 66:20:@44632.4]
  wire  regs_197_clock; // @[RegFile.scala 66:20:@44646.4]
  wire  regs_197_reset; // @[RegFile.scala 66:20:@44646.4]
  wire [63:0] regs_197_io_in; // @[RegFile.scala 66:20:@44646.4]
  wire  regs_197_io_reset; // @[RegFile.scala 66:20:@44646.4]
  wire [63:0] regs_197_io_out; // @[RegFile.scala 66:20:@44646.4]
  wire  regs_197_io_enable; // @[RegFile.scala 66:20:@44646.4]
  wire  regs_198_clock; // @[RegFile.scala 66:20:@44660.4]
  wire  regs_198_reset; // @[RegFile.scala 66:20:@44660.4]
  wire [63:0] regs_198_io_in; // @[RegFile.scala 66:20:@44660.4]
  wire  regs_198_io_reset; // @[RegFile.scala 66:20:@44660.4]
  wire [63:0] regs_198_io_out; // @[RegFile.scala 66:20:@44660.4]
  wire  regs_198_io_enable; // @[RegFile.scala 66:20:@44660.4]
  wire  regs_199_clock; // @[RegFile.scala 66:20:@44674.4]
  wire  regs_199_reset; // @[RegFile.scala 66:20:@44674.4]
  wire [63:0] regs_199_io_in; // @[RegFile.scala 66:20:@44674.4]
  wire  regs_199_io_reset; // @[RegFile.scala 66:20:@44674.4]
  wire [63:0] regs_199_io_out; // @[RegFile.scala 66:20:@44674.4]
  wire  regs_199_io_enable; // @[RegFile.scala 66:20:@44674.4]
  wire  regs_200_clock; // @[RegFile.scala 66:20:@44688.4]
  wire  regs_200_reset; // @[RegFile.scala 66:20:@44688.4]
  wire [63:0] regs_200_io_in; // @[RegFile.scala 66:20:@44688.4]
  wire  regs_200_io_reset; // @[RegFile.scala 66:20:@44688.4]
  wire [63:0] regs_200_io_out; // @[RegFile.scala 66:20:@44688.4]
  wire  regs_200_io_enable; // @[RegFile.scala 66:20:@44688.4]
  wire  regs_201_clock; // @[RegFile.scala 66:20:@44702.4]
  wire  regs_201_reset; // @[RegFile.scala 66:20:@44702.4]
  wire [63:0] regs_201_io_in; // @[RegFile.scala 66:20:@44702.4]
  wire  regs_201_io_reset; // @[RegFile.scala 66:20:@44702.4]
  wire [63:0] regs_201_io_out; // @[RegFile.scala 66:20:@44702.4]
  wire  regs_201_io_enable; // @[RegFile.scala 66:20:@44702.4]
  wire  regs_202_clock; // @[RegFile.scala 66:20:@44716.4]
  wire  regs_202_reset; // @[RegFile.scala 66:20:@44716.4]
  wire [63:0] regs_202_io_in; // @[RegFile.scala 66:20:@44716.4]
  wire  regs_202_io_reset; // @[RegFile.scala 66:20:@44716.4]
  wire [63:0] regs_202_io_out; // @[RegFile.scala 66:20:@44716.4]
  wire  regs_202_io_enable; // @[RegFile.scala 66:20:@44716.4]
  wire  regs_203_clock; // @[RegFile.scala 66:20:@44730.4]
  wire  regs_203_reset; // @[RegFile.scala 66:20:@44730.4]
  wire [63:0] regs_203_io_in; // @[RegFile.scala 66:20:@44730.4]
  wire  regs_203_io_reset; // @[RegFile.scala 66:20:@44730.4]
  wire [63:0] regs_203_io_out; // @[RegFile.scala 66:20:@44730.4]
  wire  regs_203_io_enable; // @[RegFile.scala 66:20:@44730.4]
  wire  regs_204_clock; // @[RegFile.scala 66:20:@44744.4]
  wire  regs_204_reset; // @[RegFile.scala 66:20:@44744.4]
  wire [63:0] regs_204_io_in; // @[RegFile.scala 66:20:@44744.4]
  wire  regs_204_io_reset; // @[RegFile.scala 66:20:@44744.4]
  wire [63:0] regs_204_io_out; // @[RegFile.scala 66:20:@44744.4]
  wire  regs_204_io_enable; // @[RegFile.scala 66:20:@44744.4]
  wire  regs_205_clock; // @[RegFile.scala 66:20:@44758.4]
  wire  regs_205_reset; // @[RegFile.scala 66:20:@44758.4]
  wire [63:0] regs_205_io_in; // @[RegFile.scala 66:20:@44758.4]
  wire  regs_205_io_reset; // @[RegFile.scala 66:20:@44758.4]
  wire [63:0] regs_205_io_out; // @[RegFile.scala 66:20:@44758.4]
  wire  regs_205_io_enable; // @[RegFile.scala 66:20:@44758.4]
  wire  regs_206_clock; // @[RegFile.scala 66:20:@44772.4]
  wire  regs_206_reset; // @[RegFile.scala 66:20:@44772.4]
  wire [63:0] regs_206_io_in; // @[RegFile.scala 66:20:@44772.4]
  wire  regs_206_io_reset; // @[RegFile.scala 66:20:@44772.4]
  wire [63:0] regs_206_io_out; // @[RegFile.scala 66:20:@44772.4]
  wire  regs_206_io_enable; // @[RegFile.scala 66:20:@44772.4]
  wire  regs_207_clock; // @[RegFile.scala 66:20:@44786.4]
  wire  regs_207_reset; // @[RegFile.scala 66:20:@44786.4]
  wire [63:0] regs_207_io_in; // @[RegFile.scala 66:20:@44786.4]
  wire  regs_207_io_reset; // @[RegFile.scala 66:20:@44786.4]
  wire [63:0] regs_207_io_out; // @[RegFile.scala 66:20:@44786.4]
  wire  regs_207_io_enable; // @[RegFile.scala 66:20:@44786.4]
  wire  regs_208_clock; // @[RegFile.scala 66:20:@44800.4]
  wire  regs_208_reset; // @[RegFile.scala 66:20:@44800.4]
  wire [63:0] regs_208_io_in; // @[RegFile.scala 66:20:@44800.4]
  wire  regs_208_io_reset; // @[RegFile.scala 66:20:@44800.4]
  wire [63:0] regs_208_io_out; // @[RegFile.scala 66:20:@44800.4]
  wire  regs_208_io_enable; // @[RegFile.scala 66:20:@44800.4]
  wire  regs_209_clock; // @[RegFile.scala 66:20:@44814.4]
  wire  regs_209_reset; // @[RegFile.scala 66:20:@44814.4]
  wire [63:0] regs_209_io_in; // @[RegFile.scala 66:20:@44814.4]
  wire  regs_209_io_reset; // @[RegFile.scala 66:20:@44814.4]
  wire [63:0] regs_209_io_out; // @[RegFile.scala 66:20:@44814.4]
  wire  regs_209_io_enable; // @[RegFile.scala 66:20:@44814.4]
  wire  regs_210_clock; // @[RegFile.scala 66:20:@44828.4]
  wire  regs_210_reset; // @[RegFile.scala 66:20:@44828.4]
  wire [63:0] regs_210_io_in; // @[RegFile.scala 66:20:@44828.4]
  wire  regs_210_io_reset; // @[RegFile.scala 66:20:@44828.4]
  wire [63:0] regs_210_io_out; // @[RegFile.scala 66:20:@44828.4]
  wire  regs_210_io_enable; // @[RegFile.scala 66:20:@44828.4]
  wire  regs_211_clock; // @[RegFile.scala 66:20:@44842.4]
  wire  regs_211_reset; // @[RegFile.scala 66:20:@44842.4]
  wire [63:0] regs_211_io_in; // @[RegFile.scala 66:20:@44842.4]
  wire  regs_211_io_reset; // @[RegFile.scala 66:20:@44842.4]
  wire [63:0] regs_211_io_out; // @[RegFile.scala 66:20:@44842.4]
  wire  regs_211_io_enable; // @[RegFile.scala 66:20:@44842.4]
  wire  regs_212_clock; // @[RegFile.scala 66:20:@44856.4]
  wire  regs_212_reset; // @[RegFile.scala 66:20:@44856.4]
  wire [63:0] regs_212_io_in; // @[RegFile.scala 66:20:@44856.4]
  wire  regs_212_io_reset; // @[RegFile.scala 66:20:@44856.4]
  wire [63:0] regs_212_io_out; // @[RegFile.scala 66:20:@44856.4]
  wire  regs_212_io_enable; // @[RegFile.scala 66:20:@44856.4]
  wire  regs_213_clock; // @[RegFile.scala 66:20:@44870.4]
  wire  regs_213_reset; // @[RegFile.scala 66:20:@44870.4]
  wire [63:0] regs_213_io_in; // @[RegFile.scala 66:20:@44870.4]
  wire  regs_213_io_reset; // @[RegFile.scala 66:20:@44870.4]
  wire [63:0] regs_213_io_out; // @[RegFile.scala 66:20:@44870.4]
  wire  regs_213_io_enable; // @[RegFile.scala 66:20:@44870.4]
  wire  regs_214_clock; // @[RegFile.scala 66:20:@44884.4]
  wire  regs_214_reset; // @[RegFile.scala 66:20:@44884.4]
  wire [63:0] regs_214_io_in; // @[RegFile.scala 66:20:@44884.4]
  wire  regs_214_io_reset; // @[RegFile.scala 66:20:@44884.4]
  wire [63:0] regs_214_io_out; // @[RegFile.scala 66:20:@44884.4]
  wire  regs_214_io_enable; // @[RegFile.scala 66:20:@44884.4]
  wire  regs_215_clock; // @[RegFile.scala 66:20:@44898.4]
  wire  regs_215_reset; // @[RegFile.scala 66:20:@44898.4]
  wire [63:0] regs_215_io_in; // @[RegFile.scala 66:20:@44898.4]
  wire  regs_215_io_reset; // @[RegFile.scala 66:20:@44898.4]
  wire [63:0] regs_215_io_out; // @[RegFile.scala 66:20:@44898.4]
  wire  regs_215_io_enable; // @[RegFile.scala 66:20:@44898.4]
  wire  regs_216_clock; // @[RegFile.scala 66:20:@44912.4]
  wire  regs_216_reset; // @[RegFile.scala 66:20:@44912.4]
  wire [63:0] regs_216_io_in; // @[RegFile.scala 66:20:@44912.4]
  wire  regs_216_io_reset; // @[RegFile.scala 66:20:@44912.4]
  wire [63:0] regs_216_io_out; // @[RegFile.scala 66:20:@44912.4]
  wire  regs_216_io_enable; // @[RegFile.scala 66:20:@44912.4]
  wire  regs_217_clock; // @[RegFile.scala 66:20:@44926.4]
  wire  regs_217_reset; // @[RegFile.scala 66:20:@44926.4]
  wire [63:0] regs_217_io_in; // @[RegFile.scala 66:20:@44926.4]
  wire  regs_217_io_reset; // @[RegFile.scala 66:20:@44926.4]
  wire [63:0] regs_217_io_out; // @[RegFile.scala 66:20:@44926.4]
  wire  regs_217_io_enable; // @[RegFile.scala 66:20:@44926.4]
  wire  regs_218_clock; // @[RegFile.scala 66:20:@44940.4]
  wire  regs_218_reset; // @[RegFile.scala 66:20:@44940.4]
  wire [63:0] regs_218_io_in; // @[RegFile.scala 66:20:@44940.4]
  wire  regs_218_io_reset; // @[RegFile.scala 66:20:@44940.4]
  wire [63:0] regs_218_io_out; // @[RegFile.scala 66:20:@44940.4]
  wire  regs_218_io_enable; // @[RegFile.scala 66:20:@44940.4]
  wire  regs_219_clock; // @[RegFile.scala 66:20:@44954.4]
  wire  regs_219_reset; // @[RegFile.scala 66:20:@44954.4]
  wire [63:0] regs_219_io_in; // @[RegFile.scala 66:20:@44954.4]
  wire  regs_219_io_reset; // @[RegFile.scala 66:20:@44954.4]
  wire [63:0] regs_219_io_out; // @[RegFile.scala 66:20:@44954.4]
  wire  regs_219_io_enable; // @[RegFile.scala 66:20:@44954.4]
  wire  regs_220_clock; // @[RegFile.scala 66:20:@44968.4]
  wire  regs_220_reset; // @[RegFile.scala 66:20:@44968.4]
  wire [63:0] regs_220_io_in; // @[RegFile.scala 66:20:@44968.4]
  wire  regs_220_io_reset; // @[RegFile.scala 66:20:@44968.4]
  wire [63:0] regs_220_io_out; // @[RegFile.scala 66:20:@44968.4]
  wire  regs_220_io_enable; // @[RegFile.scala 66:20:@44968.4]
  wire  regs_221_clock; // @[RegFile.scala 66:20:@44982.4]
  wire  regs_221_reset; // @[RegFile.scala 66:20:@44982.4]
  wire [63:0] regs_221_io_in; // @[RegFile.scala 66:20:@44982.4]
  wire  regs_221_io_reset; // @[RegFile.scala 66:20:@44982.4]
  wire [63:0] regs_221_io_out; // @[RegFile.scala 66:20:@44982.4]
  wire  regs_221_io_enable; // @[RegFile.scala 66:20:@44982.4]
  wire  regs_222_clock; // @[RegFile.scala 66:20:@44996.4]
  wire  regs_222_reset; // @[RegFile.scala 66:20:@44996.4]
  wire [63:0] regs_222_io_in; // @[RegFile.scala 66:20:@44996.4]
  wire  regs_222_io_reset; // @[RegFile.scala 66:20:@44996.4]
  wire [63:0] regs_222_io_out; // @[RegFile.scala 66:20:@44996.4]
  wire  regs_222_io_enable; // @[RegFile.scala 66:20:@44996.4]
  wire  regs_223_clock; // @[RegFile.scala 66:20:@45010.4]
  wire  regs_223_reset; // @[RegFile.scala 66:20:@45010.4]
  wire [63:0] regs_223_io_in; // @[RegFile.scala 66:20:@45010.4]
  wire  regs_223_io_reset; // @[RegFile.scala 66:20:@45010.4]
  wire [63:0] regs_223_io_out; // @[RegFile.scala 66:20:@45010.4]
  wire  regs_223_io_enable; // @[RegFile.scala 66:20:@45010.4]
  wire  regs_224_clock; // @[RegFile.scala 66:20:@45024.4]
  wire  regs_224_reset; // @[RegFile.scala 66:20:@45024.4]
  wire [63:0] regs_224_io_in; // @[RegFile.scala 66:20:@45024.4]
  wire  regs_224_io_reset; // @[RegFile.scala 66:20:@45024.4]
  wire [63:0] regs_224_io_out; // @[RegFile.scala 66:20:@45024.4]
  wire  regs_224_io_enable; // @[RegFile.scala 66:20:@45024.4]
  wire  regs_225_clock; // @[RegFile.scala 66:20:@45038.4]
  wire  regs_225_reset; // @[RegFile.scala 66:20:@45038.4]
  wire [63:0] regs_225_io_in; // @[RegFile.scala 66:20:@45038.4]
  wire  regs_225_io_reset; // @[RegFile.scala 66:20:@45038.4]
  wire [63:0] regs_225_io_out; // @[RegFile.scala 66:20:@45038.4]
  wire  regs_225_io_enable; // @[RegFile.scala 66:20:@45038.4]
  wire  regs_226_clock; // @[RegFile.scala 66:20:@45052.4]
  wire  regs_226_reset; // @[RegFile.scala 66:20:@45052.4]
  wire [63:0] regs_226_io_in; // @[RegFile.scala 66:20:@45052.4]
  wire  regs_226_io_reset; // @[RegFile.scala 66:20:@45052.4]
  wire [63:0] regs_226_io_out; // @[RegFile.scala 66:20:@45052.4]
  wire  regs_226_io_enable; // @[RegFile.scala 66:20:@45052.4]
  wire  regs_227_clock; // @[RegFile.scala 66:20:@45066.4]
  wire  regs_227_reset; // @[RegFile.scala 66:20:@45066.4]
  wire [63:0] regs_227_io_in; // @[RegFile.scala 66:20:@45066.4]
  wire  regs_227_io_reset; // @[RegFile.scala 66:20:@45066.4]
  wire [63:0] regs_227_io_out; // @[RegFile.scala 66:20:@45066.4]
  wire  regs_227_io_enable; // @[RegFile.scala 66:20:@45066.4]
  wire  regs_228_clock; // @[RegFile.scala 66:20:@45080.4]
  wire  regs_228_reset; // @[RegFile.scala 66:20:@45080.4]
  wire [63:0] regs_228_io_in; // @[RegFile.scala 66:20:@45080.4]
  wire  regs_228_io_reset; // @[RegFile.scala 66:20:@45080.4]
  wire [63:0] regs_228_io_out; // @[RegFile.scala 66:20:@45080.4]
  wire  regs_228_io_enable; // @[RegFile.scala 66:20:@45080.4]
  wire  regs_229_clock; // @[RegFile.scala 66:20:@45094.4]
  wire  regs_229_reset; // @[RegFile.scala 66:20:@45094.4]
  wire [63:0] regs_229_io_in; // @[RegFile.scala 66:20:@45094.4]
  wire  regs_229_io_reset; // @[RegFile.scala 66:20:@45094.4]
  wire [63:0] regs_229_io_out; // @[RegFile.scala 66:20:@45094.4]
  wire  regs_229_io_enable; // @[RegFile.scala 66:20:@45094.4]
  wire  regs_230_clock; // @[RegFile.scala 66:20:@45108.4]
  wire  regs_230_reset; // @[RegFile.scala 66:20:@45108.4]
  wire [63:0] regs_230_io_in; // @[RegFile.scala 66:20:@45108.4]
  wire  regs_230_io_reset; // @[RegFile.scala 66:20:@45108.4]
  wire [63:0] regs_230_io_out; // @[RegFile.scala 66:20:@45108.4]
  wire  regs_230_io_enable; // @[RegFile.scala 66:20:@45108.4]
  wire  regs_231_clock; // @[RegFile.scala 66:20:@45122.4]
  wire  regs_231_reset; // @[RegFile.scala 66:20:@45122.4]
  wire [63:0] regs_231_io_in; // @[RegFile.scala 66:20:@45122.4]
  wire  regs_231_io_reset; // @[RegFile.scala 66:20:@45122.4]
  wire [63:0] regs_231_io_out; // @[RegFile.scala 66:20:@45122.4]
  wire  regs_231_io_enable; // @[RegFile.scala 66:20:@45122.4]
  wire  regs_232_clock; // @[RegFile.scala 66:20:@45136.4]
  wire  regs_232_reset; // @[RegFile.scala 66:20:@45136.4]
  wire [63:0] regs_232_io_in; // @[RegFile.scala 66:20:@45136.4]
  wire  regs_232_io_reset; // @[RegFile.scala 66:20:@45136.4]
  wire [63:0] regs_232_io_out; // @[RegFile.scala 66:20:@45136.4]
  wire  regs_232_io_enable; // @[RegFile.scala 66:20:@45136.4]
  wire  regs_233_clock; // @[RegFile.scala 66:20:@45150.4]
  wire  regs_233_reset; // @[RegFile.scala 66:20:@45150.4]
  wire [63:0] regs_233_io_in; // @[RegFile.scala 66:20:@45150.4]
  wire  regs_233_io_reset; // @[RegFile.scala 66:20:@45150.4]
  wire [63:0] regs_233_io_out; // @[RegFile.scala 66:20:@45150.4]
  wire  regs_233_io_enable; // @[RegFile.scala 66:20:@45150.4]
  wire  regs_234_clock; // @[RegFile.scala 66:20:@45164.4]
  wire  regs_234_reset; // @[RegFile.scala 66:20:@45164.4]
  wire [63:0] regs_234_io_in; // @[RegFile.scala 66:20:@45164.4]
  wire  regs_234_io_reset; // @[RegFile.scala 66:20:@45164.4]
  wire [63:0] regs_234_io_out; // @[RegFile.scala 66:20:@45164.4]
  wire  regs_234_io_enable; // @[RegFile.scala 66:20:@45164.4]
  wire  regs_235_clock; // @[RegFile.scala 66:20:@45178.4]
  wire  regs_235_reset; // @[RegFile.scala 66:20:@45178.4]
  wire [63:0] regs_235_io_in; // @[RegFile.scala 66:20:@45178.4]
  wire  regs_235_io_reset; // @[RegFile.scala 66:20:@45178.4]
  wire [63:0] regs_235_io_out; // @[RegFile.scala 66:20:@45178.4]
  wire  regs_235_io_enable; // @[RegFile.scala 66:20:@45178.4]
  wire  regs_236_clock; // @[RegFile.scala 66:20:@45192.4]
  wire  regs_236_reset; // @[RegFile.scala 66:20:@45192.4]
  wire [63:0] regs_236_io_in; // @[RegFile.scala 66:20:@45192.4]
  wire  regs_236_io_reset; // @[RegFile.scala 66:20:@45192.4]
  wire [63:0] regs_236_io_out; // @[RegFile.scala 66:20:@45192.4]
  wire  regs_236_io_enable; // @[RegFile.scala 66:20:@45192.4]
  wire  regs_237_clock; // @[RegFile.scala 66:20:@45206.4]
  wire  regs_237_reset; // @[RegFile.scala 66:20:@45206.4]
  wire [63:0] regs_237_io_in; // @[RegFile.scala 66:20:@45206.4]
  wire  regs_237_io_reset; // @[RegFile.scala 66:20:@45206.4]
  wire [63:0] regs_237_io_out; // @[RegFile.scala 66:20:@45206.4]
  wire  regs_237_io_enable; // @[RegFile.scala 66:20:@45206.4]
  wire  regs_238_clock; // @[RegFile.scala 66:20:@45220.4]
  wire  regs_238_reset; // @[RegFile.scala 66:20:@45220.4]
  wire [63:0] regs_238_io_in; // @[RegFile.scala 66:20:@45220.4]
  wire  regs_238_io_reset; // @[RegFile.scala 66:20:@45220.4]
  wire [63:0] regs_238_io_out; // @[RegFile.scala 66:20:@45220.4]
  wire  regs_238_io_enable; // @[RegFile.scala 66:20:@45220.4]
  wire  regs_239_clock; // @[RegFile.scala 66:20:@45234.4]
  wire  regs_239_reset; // @[RegFile.scala 66:20:@45234.4]
  wire [63:0] regs_239_io_in; // @[RegFile.scala 66:20:@45234.4]
  wire  regs_239_io_reset; // @[RegFile.scala 66:20:@45234.4]
  wire [63:0] regs_239_io_out; // @[RegFile.scala 66:20:@45234.4]
  wire  regs_239_io_enable; // @[RegFile.scala 66:20:@45234.4]
  wire  regs_240_clock; // @[RegFile.scala 66:20:@45248.4]
  wire  regs_240_reset; // @[RegFile.scala 66:20:@45248.4]
  wire [63:0] regs_240_io_in; // @[RegFile.scala 66:20:@45248.4]
  wire  regs_240_io_reset; // @[RegFile.scala 66:20:@45248.4]
  wire [63:0] regs_240_io_out; // @[RegFile.scala 66:20:@45248.4]
  wire  regs_240_io_enable; // @[RegFile.scala 66:20:@45248.4]
  wire  regs_241_clock; // @[RegFile.scala 66:20:@45262.4]
  wire  regs_241_reset; // @[RegFile.scala 66:20:@45262.4]
  wire [63:0] regs_241_io_in; // @[RegFile.scala 66:20:@45262.4]
  wire  regs_241_io_reset; // @[RegFile.scala 66:20:@45262.4]
  wire [63:0] regs_241_io_out; // @[RegFile.scala 66:20:@45262.4]
  wire  regs_241_io_enable; // @[RegFile.scala 66:20:@45262.4]
  wire  regs_242_clock; // @[RegFile.scala 66:20:@45276.4]
  wire  regs_242_reset; // @[RegFile.scala 66:20:@45276.4]
  wire [63:0] regs_242_io_in; // @[RegFile.scala 66:20:@45276.4]
  wire  regs_242_io_reset; // @[RegFile.scala 66:20:@45276.4]
  wire [63:0] regs_242_io_out; // @[RegFile.scala 66:20:@45276.4]
  wire  regs_242_io_enable; // @[RegFile.scala 66:20:@45276.4]
  wire  regs_243_clock; // @[RegFile.scala 66:20:@45290.4]
  wire  regs_243_reset; // @[RegFile.scala 66:20:@45290.4]
  wire [63:0] regs_243_io_in; // @[RegFile.scala 66:20:@45290.4]
  wire  regs_243_io_reset; // @[RegFile.scala 66:20:@45290.4]
  wire [63:0] regs_243_io_out; // @[RegFile.scala 66:20:@45290.4]
  wire  regs_243_io_enable; // @[RegFile.scala 66:20:@45290.4]
  wire  regs_244_clock; // @[RegFile.scala 66:20:@45304.4]
  wire  regs_244_reset; // @[RegFile.scala 66:20:@45304.4]
  wire [63:0] regs_244_io_in; // @[RegFile.scala 66:20:@45304.4]
  wire  regs_244_io_reset; // @[RegFile.scala 66:20:@45304.4]
  wire [63:0] regs_244_io_out; // @[RegFile.scala 66:20:@45304.4]
  wire  regs_244_io_enable; // @[RegFile.scala 66:20:@45304.4]
  wire  regs_245_clock; // @[RegFile.scala 66:20:@45318.4]
  wire  regs_245_reset; // @[RegFile.scala 66:20:@45318.4]
  wire [63:0] regs_245_io_in; // @[RegFile.scala 66:20:@45318.4]
  wire  regs_245_io_reset; // @[RegFile.scala 66:20:@45318.4]
  wire [63:0] regs_245_io_out; // @[RegFile.scala 66:20:@45318.4]
  wire  regs_245_io_enable; // @[RegFile.scala 66:20:@45318.4]
  wire  regs_246_clock; // @[RegFile.scala 66:20:@45332.4]
  wire  regs_246_reset; // @[RegFile.scala 66:20:@45332.4]
  wire [63:0] regs_246_io_in; // @[RegFile.scala 66:20:@45332.4]
  wire  regs_246_io_reset; // @[RegFile.scala 66:20:@45332.4]
  wire [63:0] regs_246_io_out; // @[RegFile.scala 66:20:@45332.4]
  wire  regs_246_io_enable; // @[RegFile.scala 66:20:@45332.4]
  wire  regs_247_clock; // @[RegFile.scala 66:20:@45346.4]
  wire  regs_247_reset; // @[RegFile.scala 66:20:@45346.4]
  wire [63:0] regs_247_io_in; // @[RegFile.scala 66:20:@45346.4]
  wire  regs_247_io_reset; // @[RegFile.scala 66:20:@45346.4]
  wire [63:0] regs_247_io_out; // @[RegFile.scala 66:20:@45346.4]
  wire  regs_247_io_enable; // @[RegFile.scala 66:20:@45346.4]
  wire  regs_248_clock; // @[RegFile.scala 66:20:@45360.4]
  wire  regs_248_reset; // @[RegFile.scala 66:20:@45360.4]
  wire [63:0] regs_248_io_in; // @[RegFile.scala 66:20:@45360.4]
  wire  regs_248_io_reset; // @[RegFile.scala 66:20:@45360.4]
  wire [63:0] regs_248_io_out; // @[RegFile.scala 66:20:@45360.4]
  wire  regs_248_io_enable; // @[RegFile.scala 66:20:@45360.4]
  wire  regs_249_clock; // @[RegFile.scala 66:20:@45374.4]
  wire  regs_249_reset; // @[RegFile.scala 66:20:@45374.4]
  wire [63:0] regs_249_io_in; // @[RegFile.scala 66:20:@45374.4]
  wire  regs_249_io_reset; // @[RegFile.scala 66:20:@45374.4]
  wire [63:0] regs_249_io_out; // @[RegFile.scala 66:20:@45374.4]
  wire  regs_249_io_enable; // @[RegFile.scala 66:20:@45374.4]
  wire  regs_250_clock; // @[RegFile.scala 66:20:@45388.4]
  wire  regs_250_reset; // @[RegFile.scala 66:20:@45388.4]
  wire [63:0] regs_250_io_in; // @[RegFile.scala 66:20:@45388.4]
  wire  regs_250_io_reset; // @[RegFile.scala 66:20:@45388.4]
  wire [63:0] regs_250_io_out; // @[RegFile.scala 66:20:@45388.4]
  wire  regs_250_io_enable; // @[RegFile.scala 66:20:@45388.4]
  wire  regs_251_clock; // @[RegFile.scala 66:20:@45402.4]
  wire  regs_251_reset; // @[RegFile.scala 66:20:@45402.4]
  wire [63:0] regs_251_io_in; // @[RegFile.scala 66:20:@45402.4]
  wire  regs_251_io_reset; // @[RegFile.scala 66:20:@45402.4]
  wire [63:0] regs_251_io_out; // @[RegFile.scala 66:20:@45402.4]
  wire  regs_251_io_enable; // @[RegFile.scala 66:20:@45402.4]
  wire  regs_252_clock; // @[RegFile.scala 66:20:@45416.4]
  wire  regs_252_reset; // @[RegFile.scala 66:20:@45416.4]
  wire [63:0] regs_252_io_in; // @[RegFile.scala 66:20:@45416.4]
  wire  regs_252_io_reset; // @[RegFile.scala 66:20:@45416.4]
  wire [63:0] regs_252_io_out; // @[RegFile.scala 66:20:@45416.4]
  wire  regs_252_io_enable; // @[RegFile.scala 66:20:@45416.4]
  wire  regs_253_clock; // @[RegFile.scala 66:20:@45430.4]
  wire  regs_253_reset; // @[RegFile.scala 66:20:@45430.4]
  wire [63:0] regs_253_io_in; // @[RegFile.scala 66:20:@45430.4]
  wire  regs_253_io_reset; // @[RegFile.scala 66:20:@45430.4]
  wire [63:0] regs_253_io_out; // @[RegFile.scala 66:20:@45430.4]
  wire  regs_253_io_enable; // @[RegFile.scala 66:20:@45430.4]
  wire  regs_254_clock; // @[RegFile.scala 66:20:@45444.4]
  wire  regs_254_reset; // @[RegFile.scala 66:20:@45444.4]
  wire [63:0] regs_254_io_in; // @[RegFile.scala 66:20:@45444.4]
  wire  regs_254_io_reset; // @[RegFile.scala 66:20:@45444.4]
  wire [63:0] regs_254_io_out; // @[RegFile.scala 66:20:@45444.4]
  wire  regs_254_io_enable; // @[RegFile.scala 66:20:@45444.4]
  wire  regs_255_clock; // @[RegFile.scala 66:20:@45458.4]
  wire  regs_255_reset; // @[RegFile.scala 66:20:@45458.4]
  wire [63:0] regs_255_io_in; // @[RegFile.scala 66:20:@45458.4]
  wire  regs_255_io_reset; // @[RegFile.scala 66:20:@45458.4]
  wire [63:0] regs_255_io_out; // @[RegFile.scala 66:20:@45458.4]
  wire  regs_255_io_enable; // @[RegFile.scala 66:20:@45458.4]
  wire  regs_256_clock; // @[RegFile.scala 66:20:@45472.4]
  wire  regs_256_reset; // @[RegFile.scala 66:20:@45472.4]
  wire [63:0] regs_256_io_in; // @[RegFile.scala 66:20:@45472.4]
  wire  regs_256_io_reset; // @[RegFile.scala 66:20:@45472.4]
  wire [63:0] regs_256_io_out; // @[RegFile.scala 66:20:@45472.4]
  wire  regs_256_io_enable; // @[RegFile.scala 66:20:@45472.4]
  wire  regs_257_clock; // @[RegFile.scala 66:20:@45486.4]
  wire  regs_257_reset; // @[RegFile.scala 66:20:@45486.4]
  wire [63:0] regs_257_io_in; // @[RegFile.scala 66:20:@45486.4]
  wire  regs_257_io_reset; // @[RegFile.scala 66:20:@45486.4]
  wire [63:0] regs_257_io_out; // @[RegFile.scala 66:20:@45486.4]
  wire  regs_257_io_enable; // @[RegFile.scala 66:20:@45486.4]
  wire  regs_258_clock; // @[RegFile.scala 66:20:@45500.4]
  wire  regs_258_reset; // @[RegFile.scala 66:20:@45500.4]
  wire [63:0] regs_258_io_in; // @[RegFile.scala 66:20:@45500.4]
  wire  regs_258_io_reset; // @[RegFile.scala 66:20:@45500.4]
  wire [63:0] regs_258_io_out; // @[RegFile.scala 66:20:@45500.4]
  wire  regs_258_io_enable; // @[RegFile.scala 66:20:@45500.4]
  wire  regs_259_clock; // @[RegFile.scala 66:20:@45514.4]
  wire  regs_259_reset; // @[RegFile.scala 66:20:@45514.4]
  wire [63:0] regs_259_io_in; // @[RegFile.scala 66:20:@45514.4]
  wire  regs_259_io_reset; // @[RegFile.scala 66:20:@45514.4]
  wire [63:0] regs_259_io_out; // @[RegFile.scala 66:20:@45514.4]
  wire  regs_259_io_enable; // @[RegFile.scala 66:20:@45514.4]
  wire  regs_260_clock; // @[RegFile.scala 66:20:@45528.4]
  wire  regs_260_reset; // @[RegFile.scala 66:20:@45528.4]
  wire [63:0] regs_260_io_in; // @[RegFile.scala 66:20:@45528.4]
  wire  regs_260_io_reset; // @[RegFile.scala 66:20:@45528.4]
  wire [63:0] regs_260_io_out; // @[RegFile.scala 66:20:@45528.4]
  wire  regs_260_io_enable; // @[RegFile.scala 66:20:@45528.4]
  wire  regs_261_clock; // @[RegFile.scala 66:20:@45542.4]
  wire  regs_261_reset; // @[RegFile.scala 66:20:@45542.4]
  wire [63:0] regs_261_io_in; // @[RegFile.scala 66:20:@45542.4]
  wire  regs_261_io_reset; // @[RegFile.scala 66:20:@45542.4]
  wire [63:0] regs_261_io_out; // @[RegFile.scala 66:20:@45542.4]
  wire  regs_261_io_enable; // @[RegFile.scala 66:20:@45542.4]
  wire  regs_262_clock; // @[RegFile.scala 66:20:@45556.4]
  wire  regs_262_reset; // @[RegFile.scala 66:20:@45556.4]
  wire [63:0] regs_262_io_in; // @[RegFile.scala 66:20:@45556.4]
  wire  regs_262_io_reset; // @[RegFile.scala 66:20:@45556.4]
  wire [63:0] regs_262_io_out; // @[RegFile.scala 66:20:@45556.4]
  wire  regs_262_io_enable; // @[RegFile.scala 66:20:@45556.4]
  wire  regs_263_clock; // @[RegFile.scala 66:20:@45570.4]
  wire  regs_263_reset; // @[RegFile.scala 66:20:@45570.4]
  wire [63:0] regs_263_io_in; // @[RegFile.scala 66:20:@45570.4]
  wire  regs_263_io_reset; // @[RegFile.scala 66:20:@45570.4]
  wire [63:0] regs_263_io_out; // @[RegFile.scala 66:20:@45570.4]
  wire  regs_263_io_enable; // @[RegFile.scala 66:20:@45570.4]
  wire  regs_264_clock; // @[RegFile.scala 66:20:@45584.4]
  wire  regs_264_reset; // @[RegFile.scala 66:20:@45584.4]
  wire [63:0] regs_264_io_in; // @[RegFile.scala 66:20:@45584.4]
  wire  regs_264_io_reset; // @[RegFile.scala 66:20:@45584.4]
  wire [63:0] regs_264_io_out; // @[RegFile.scala 66:20:@45584.4]
  wire  regs_264_io_enable; // @[RegFile.scala 66:20:@45584.4]
  wire  regs_265_clock; // @[RegFile.scala 66:20:@45598.4]
  wire  regs_265_reset; // @[RegFile.scala 66:20:@45598.4]
  wire [63:0] regs_265_io_in; // @[RegFile.scala 66:20:@45598.4]
  wire  regs_265_io_reset; // @[RegFile.scala 66:20:@45598.4]
  wire [63:0] regs_265_io_out; // @[RegFile.scala 66:20:@45598.4]
  wire  regs_265_io_enable; // @[RegFile.scala 66:20:@45598.4]
  wire  regs_266_clock; // @[RegFile.scala 66:20:@45612.4]
  wire  regs_266_reset; // @[RegFile.scala 66:20:@45612.4]
  wire [63:0] regs_266_io_in; // @[RegFile.scala 66:20:@45612.4]
  wire  regs_266_io_reset; // @[RegFile.scala 66:20:@45612.4]
  wire [63:0] regs_266_io_out; // @[RegFile.scala 66:20:@45612.4]
  wire  regs_266_io_enable; // @[RegFile.scala 66:20:@45612.4]
  wire  regs_267_clock; // @[RegFile.scala 66:20:@45626.4]
  wire  regs_267_reset; // @[RegFile.scala 66:20:@45626.4]
  wire [63:0] regs_267_io_in; // @[RegFile.scala 66:20:@45626.4]
  wire  regs_267_io_reset; // @[RegFile.scala 66:20:@45626.4]
  wire [63:0] regs_267_io_out; // @[RegFile.scala 66:20:@45626.4]
  wire  regs_267_io_enable; // @[RegFile.scala 66:20:@45626.4]
  wire  regs_268_clock; // @[RegFile.scala 66:20:@45640.4]
  wire  regs_268_reset; // @[RegFile.scala 66:20:@45640.4]
  wire [63:0] regs_268_io_in; // @[RegFile.scala 66:20:@45640.4]
  wire  regs_268_io_reset; // @[RegFile.scala 66:20:@45640.4]
  wire [63:0] regs_268_io_out; // @[RegFile.scala 66:20:@45640.4]
  wire  regs_268_io_enable; // @[RegFile.scala 66:20:@45640.4]
  wire  regs_269_clock; // @[RegFile.scala 66:20:@45654.4]
  wire  regs_269_reset; // @[RegFile.scala 66:20:@45654.4]
  wire [63:0] regs_269_io_in; // @[RegFile.scala 66:20:@45654.4]
  wire  regs_269_io_reset; // @[RegFile.scala 66:20:@45654.4]
  wire [63:0] regs_269_io_out; // @[RegFile.scala 66:20:@45654.4]
  wire  regs_269_io_enable; // @[RegFile.scala 66:20:@45654.4]
  wire  regs_270_clock; // @[RegFile.scala 66:20:@45668.4]
  wire  regs_270_reset; // @[RegFile.scala 66:20:@45668.4]
  wire [63:0] regs_270_io_in; // @[RegFile.scala 66:20:@45668.4]
  wire  regs_270_io_reset; // @[RegFile.scala 66:20:@45668.4]
  wire [63:0] regs_270_io_out; // @[RegFile.scala 66:20:@45668.4]
  wire  regs_270_io_enable; // @[RegFile.scala 66:20:@45668.4]
  wire  regs_271_clock; // @[RegFile.scala 66:20:@45682.4]
  wire  regs_271_reset; // @[RegFile.scala 66:20:@45682.4]
  wire [63:0] regs_271_io_in; // @[RegFile.scala 66:20:@45682.4]
  wire  regs_271_io_reset; // @[RegFile.scala 66:20:@45682.4]
  wire [63:0] regs_271_io_out; // @[RegFile.scala 66:20:@45682.4]
  wire  regs_271_io_enable; // @[RegFile.scala 66:20:@45682.4]
  wire  regs_272_clock; // @[RegFile.scala 66:20:@45696.4]
  wire  regs_272_reset; // @[RegFile.scala 66:20:@45696.4]
  wire [63:0] regs_272_io_in; // @[RegFile.scala 66:20:@45696.4]
  wire  regs_272_io_reset; // @[RegFile.scala 66:20:@45696.4]
  wire [63:0] regs_272_io_out; // @[RegFile.scala 66:20:@45696.4]
  wire  regs_272_io_enable; // @[RegFile.scala 66:20:@45696.4]
  wire  regs_273_clock; // @[RegFile.scala 66:20:@45710.4]
  wire  regs_273_reset; // @[RegFile.scala 66:20:@45710.4]
  wire [63:0] regs_273_io_in; // @[RegFile.scala 66:20:@45710.4]
  wire  regs_273_io_reset; // @[RegFile.scala 66:20:@45710.4]
  wire [63:0] regs_273_io_out; // @[RegFile.scala 66:20:@45710.4]
  wire  regs_273_io_enable; // @[RegFile.scala 66:20:@45710.4]
  wire  regs_274_clock; // @[RegFile.scala 66:20:@45724.4]
  wire  regs_274_reset; // @[RegFile.scala 66:20:@45724.4]
  wire [63:0] regs_274_io_in; // @[RegFile.scala 66:20:@45724.4]
  wire  regs_274_io_reset; // @[RegFile.scala 66:20:@45724.4]
  wire [63:0] regs_274_io_out; // @[RegFile.scala 66:20:@45724.4]
  wire  regs_274_io_enable; // @[RegFile.scala 66:20:@45724.4]
  wire  regs_275_clock; // @[RegFile.scala 66:20:@45738.4]
  wire  regs_275_reset; // @[RegFile.scala 66:20:@45738.4]
  wire [63:0] regs_275_io_in; // @[RegFile.scala 66:20:@45738.4]
  wire  regs_275_io_reset; // @[RegFile.scala 66:20:@45738.4]
  wire [63:0] regs_275_io_out; // @[RegFile.scala 66:20:@45738.4]
  wire  regs_275_io_enable; // @[RegFile.scala 66:20:@45738.4]
  wire  regs_276_clock; // @[RegFile.scala 66:20:@45752.4]
  wire  regs_276_reset; // @[RegFile.scala 66:20:@45752.4]
  wire [63:0] regs_276_io_in; // @[RegFile.scala 66:20:@45752.4]
  wire  regs_276_io_reset; // @[RegFile.scala 66:20:@45752.4]
  wire [63:0] regs_276_io_out; // @[RegFile.scala 66:20:@45752.4]
  wire  regs_276_io_enable; // @[RegFile.scala 66:20:@45752.4]
  wire  regs_277_clock; // @[RegFile.scala 66:20:@45766.4]
  wire  regs_277_reset; // @[RegFile.scala 66:20:@45766.4]
  wire [63:0] regs_277_io_in; // @[RegFile.scala 66:20:@45766.4]
  wire  regs_277_io_reset; // @[RegFile.scala 66:20:@45766.4]
  wire [63:0] regs_277_io_out; // @[RegFile.scala 66:20:@45766.4]
  wire  regs_277_io_enable; // @[RegFile.scala 66:20:@45766.4]
  wire  regs_278_clock; // @[RegFile.scala 66:20:@45780.4]
  wire  regs_278_reset; // @[RegFile.scala 66:20:@45780.4]
  wire [63:0] regs_278_io_in; // @[RegFile.scala 66:20:@45780.4]
  wire  regs_278_io_reset; // @[RegFile.scala 66:20:@45780.4]
  wire [63:0] regs_278_io_out; // @[RegFile.scala 66:20:@45780.4]
  wire  regs_278_io_enable; // @[RegFile.scala 66:20:@45780.4]
  wire  regs_279_clock; // @[RegFile.scala 66:20:@45794.4]
  wire  regs_279_reset; // @[RegFile.scala 66:20:@45794.4]
  wire [63:0] regs_279_io_in; // @[RegFile.scala 66:20:@45794.4]
  wire  regs_279_io_reset; // @[RegFile.scala 66:20:@45794.4]
  wire [63:0] regs_279_io_out; // @[RegFile.scala 66:20:@45794.4]
  wire  regs_279_io_enable; // @[RegFile.scala 66:20:@45794.4]
  wire  regs_280_clock; // @[RegFile.scala 66:20:@45808.4]
  wire  regs_280_reset; // @[RegFile.scala 66:20:@45808.4]
  wire [63:0] regs_280_io_in; // @[RegFile.scala 66:20:@45808.4]
  wire  regs_280_io_reset; // @[RegFile.scala 66:20:@45808.4]
  wire [63:0] regs_280_io_out; // @[RegFile.scala 66:20:@45808.4]
  wire  regs_280_io_enable; // @[RegFile.scala 66:20:@45808.4]
  wire  regs_281_clock; // @[RegFile.scala 66:20:@45822.4]
  wire  regs_281_reset; // @[RegFile.scala 66:20:@45822.4]
  wire [63:0] regs_281_io_in; // @[RegFile.scala 66:20:@45822.4]
  wire  regs_281_io_reset; // @[RegFile.scala 66:20:@45822.4]
  wire [63:0] regs_281_io_out; // @[RegFile.scala 66:20:@45822.4]
  wire  regs_281_io_enable; // @[RegFile.scala 66:20:@45822.4]
  wire  regs_282_clock; // @[RegFile.scala 66:20:@45836.4]
  wire  regs_282_reset; // @[RegFile.scala 66:20:@45836.4]
  wire [63:0] regs_282_io_in; // @[RegFile.scala 66:20:@45836.4]
  wire  regs_282_io_reset; // @[RegFile.scala 66:20:@45836.4]
  wire [63:0] regs_282_io_out; // @[RegFile.scala 66:20:@45836.4]
  wire  regs_282_io_enable; // @[RegFile.scala 66:20:@45836.4]
  wire  regs_283_clock; // @[RegFile.scala 66:20:@45850.4]
  wire  regs_283_reset; // @[RegFile.scala 66:20:@45850.4]
  wire [63:0] regs_283_io_in; // @[RegFile.scala 66:20:@45850.4]
  wire  regs_283_io_reset; // @[RegFile.scala 66:20:@45850.4]
  wire [63:0] regs_283_io_out; // @[RegFile.scala 66:20:@45850.4]
  wire  regs_283_io_enable; // @[RegFile.scala 66:20:@45850.4]
  wire  regs_284_clock; // @[RegFile.scala 66:20:@45864.4]
  wire  regs_284_reset; // @[RegFile.scala 66:20:@45864.4]
  wire [63:0] regs_284_io_in; // @[RegFile.scala 66:20:@45864.4]
  wire  regs_284_io_reset; // @[RegFile.scala 66:20:@45864.4]
  wire [63:0] regs_284_io_out; // @[RegFile.scala 66:20:@45864.4]
  wire  regs_284_io_enable; // @[RegFile.scala 66:20:@45864.4]
  wire  regs_285_clock; // @[RegFile.scala 66:20:@45878.4]
  wire  regs_285_reset; // @[RegFile.scala 66:20:@45878.4]
  wire [63:0] regs_285_io_in; // @[RegFile.scala 66:20:@45878.4]
  wire  regs_285_io_reset; // @[RegFile.scala 66:20:@45878.4]
  wire [63:0] regs_285_io_out; // @[RegFile.scala 66:20:@45878.4]
  wire  regs_285_io_enable; // @[RegFile.scala 66:20:@45878.4]
  wire  regs_286_clock; // @[RegFile.scala 66:20:@45892.4]
  wire  regs_286_reset; // @[RegFile.scala 66:20:@45892.4]
  wire [63:0] regs_286_io_in; // @[RegFile.scala 66:20:@45892.4]
  wire  regs_286_io_reset; // @[RegFile.scala 66:20:@45892.4]
  wire [63:0] regs_286_io_out; // @[RegFile.scala 66:20:@45892.4]
  wire  regs_286_io_enable; // @[RegFile.scala 66:20:@45892.4]
  wire  regs_287_clock; // @[RegFile.scala 66:20:@45906.4]
  wire  regs_287_reset; // @[RegFile.scala 66:20:@45906.4]
  wire [63:0] regs_287_io_in; // @[RegFile.scala 66:20:@45906.4]
  wire  regs_287_io_reset; // @[RegFile.scala 66:20:@45906.4]
  wire [63:0] regs_287_io_out; // @[RegFile.scala 66:20:@45906.4]
  wire  regs_287_io_enable; // @[RegFile.scala 66:20:@45906.4]
  wire  regs_288_clock; // @[RegFile.scala 66:20:@45920.4]
  wire  regs_288_reset; // @[RegFile.scala 66:20:@45920.4]
  wire [63:0] regs_288_io_in; // @[RegFile.scala 66:20:@45920.4]
  wire  regs_288_io_reset; // @[RegFile.scala 66:20:@45920.4]
  wire [63:0] regs_288_io_out; // @[RegFile.scala 66:20:@45920.4]
  wire  regs_288_io_enable; // @[RegFile.scala 66:20:@45920.4]
  wire  regs_289_clock; // @[RegFile.scala 66:20:@45934.4]
  wire  regs_289_reset; // @[RegFile.scala 66:20:@45934.4]
  wire [63:0] regs_289_io_in; // @[RegFile.scala 66:20:@45934.4]
  wire  regs_289_io_reset; // @[RegFile.scala 66:20:@45934.4]
  wire [63:0] regs_289_io_out; // @[RegFile.scala 66:20:@45934.4]
  wire  regs_289_io_enable; // @[RegFile.scala 66:20:@45934.4]
  wire  regs_290_clock; // @[RegFile.scala 66:20:@45948.4]
  wire  regs_290_reset; // @[RegFile.scala 66:20:@45948.4]
  wire [63:0] regs_290_io_in; // @[RegFile.scala 66:20:@45948.4]
  wire  regs_290_io_reset; // @[RegFile.scala 66:20:@45948.4]
  wire [63:0] regs_290_io_out; // @[RegFile.scala 66:20:@45948.4]
  wire  regs_290_io_enable; // @[RegFile.scala 66:20:@45948.4]
  wire  regs_291_clock; // @[RegFile.scala 66:20:@45962.4]
  wire  regs_291_reset; // @[RegFile.scala 66:20:@45962.4]
  wire [63:0] regs_291_io_in; // @[RegFile.scala 66:20:@45962.4]
  wire  regs_291_io_reset; // @[RegFile.scala 66:20:@45962.4]
  wire [63:0] regs_291_io_out; // @[RegFile.scala 66:20:@45962.4]
  wire  regs_291_io_enable; // @[RegFile.scala 66:20:@45962.4]
  wire  regs_292_clock; // @[RegFile.scala 66:20:@45976.4]
  wire  regs_292_reset; // @[RegFile.scala 66:20:@45976.4]
  wire [63:0] regs_292_io_in; // @[RegFile.scala 66:20:@45976.4]
  wire  regs_292_io_reset; // @[RegFile.scala 66:20:@45976.4]
  wire [63:0] regs_292_io_out; // @[RegFile.scala 66:20:@45976.4]
  wire  regs_292_io_enable; // @[RegFile.scala 66:20:@45976.4]
  wire  regs_293_clock; // @[RegFile.scala 66:20:@45990.4]
  wire  regs_293_reset; // @[RegFile.scala 66:20:@45990.4]
  wire [63:0] regs_293_io_in; // @[RegFile.scala 66:20:@45990.4]
  wire  regs_293_io_reset; // @[RegFile.scala 66:20:@45990.4]
  wire [63:0] regs_293_io_out; // @[RegFile.scala 66:20:@45990.4]
  wire  regs_293_io_enable; // @[RegFile.scala 66:20:@45990.4]
  wire  regs_294_clock; // @[RegFile.scala 66:20:@46004.4]
  wire  regs_294_reset; // @[RegFile.scala 66:20:@46004.4]
  wire [63:0] regs_294_io_in; // @[RegFile.scala 66:20:@46004.4]
  wire  regs_294_io_reset; // @[RegFile.scala 66:20:@46004.4]
  wire [63:0] regs_294_io_out; // @[RegFile.scala 66:20:@46004.4]
  wire  regs_294_io_enable; // @[RegFile.scala 66:20:@46004.4]
  wire  regs_295_clock; // @[RegFile.scala 66:20:@46018.4]
  wire  regs_295_reset; // @[RegFile.scala 66:20:@46018.4]
  wire [63:0] regs_295_io_in; // @[RegFile.scala 66:20:@46018.4]
  wire  regs_295_io_reset; // @[RegFile.scala 66:20:@46018.4]
  wire [63:0] regs_295_io_out; // @[RegFile.scala 66:20:@46018.4]
  wire  regs_295_io_enable; // @[RegFile.scala 66:20:@46018.4]
  wire  regs_296_clock; // @[RegFile.scala 66:20:@46032.4]
  wire  regs_296_reset; // @[RegFile.scala 66:20:@46032.4]
  wire [63:0] regs_296_io_in; // @[RegFile.scala 66:20:@46032.4]
  wire  regs_296_io_reset; // @[RegFile.scala 66:20:@46032.4]
  wire [63:0] regs_296_io_out; // @[RegFile.scala 66:20:@46032.4]
  wire  regs_296_io_enable; // @[RegFile.scala 66:20:@46032.4]
  wire  regs_297_clock; // @[RegFile.scala 66:20:@46046.4]
  wire  regs_297_reset; // @[RegFile.scala 66:20:@46046.4]
  wire [63:0] regs_297_io_in; // @[RegFile.scala 66:20:@46046.4]
  wire  regs_297_io_reset; // @[RegFile.scala 66:20:@46046.4]
  wire [63:0] regs_297_io_out; // @[RegFile.scala 66:20:@46046.4]
  wire  regs_297_io_enable; // @[RegFile.scala 66:20:@46046.4]
  wire  regs_298_clock; // @[RegFile.scala 66:20:@46060.4]
  wire  regs_298_reset; // @[RegFile.scala 66:20:@46060.4]
  wire [63:0] regs_298_io_in; // @[RegFile.scala 66:20:@46060.4]
  wire  regs_298_io_reset; // @[RegFile.scala 66:20:@46060.4]
  wire [63:0] regs_298_io_out; // @[RegFile.scala 66:20:@46060.4]
  wire  regs_298_io_enable; // @[RegFile.scala 66:20:@46060.4]
  wire  regs_299_clock; // @[RegFile.scala 66:20:@46074.4]
  wire  regs_299_reset; // @[RegFile.scala 66:20:@46074.4]
  wire [63:0] regs_299_io_in; // @[RegFile.scala 66:20:@46074.4]
  wire  regs_299_io_reset; // @[RegFile.scala 66:20:@46074.4]
  wire [63:0] regs_299_io_out; // @[RegFile.scala 66:20:@46074.4]
  wire  regs_299_io_enable; // @[RegFile.scala 66:20:@46074.4]
  wire  regs_300_clock; // @[RegFile.scala 66:20:@46088.4]
  wire  regs_300_reset; // @[RegFile.scala 66:20:@46088.4]
  wire [63:0] regs_300_io_in; // @[RegFile.scala 66:20:@46088.4]
  wire  regs_300_io_reset; // @[RegFile.scala 66:20:@46088.4]
  wire [63:0] regs_300_io_out; // @[RegFile.scala 66:20:@46088.4]
  wire  regs_300_io_enable; // @[RegFile.scala 66:20:@46088.4]
  wire  regs_301_clock; // @[RegFile.scala 66:20:@46102.4]
  wire  regs_301_reset; // @[RegFile.scala 66:20:@46102.4]
  wire [63:0] regs_301_io_in; // @[RegFile.scala 66:20:@46102.4]
  wire  regs_301_io_reset; // @[RegFile.scala 66:20:@46102.4]
  wire [63:0] regs_301_io_out; // @[RegFile.scala 66:20:@46102.4]
  wire  regs_301_io_enable; // @[RegFile.scala 66:20:@46102.4]
  wire  regs_302_clock; // @[RegFile.scala 66:20:@46116.4]
  wire  regs_302_reset; // @[RegFile.scala 66:20:@46116.4]
  wire [63:0] regs_302_io_in; // @[RegFile.scala 66:20:@46116.4]
  wire  regs_302_io_reset; // @[RegFile.scala 66:20:@46116.4]
  wire [63:0] regs_302_io_out; // @[RegFile.scala 66:20:@46116.4]
  wire  regs_302_io_enable; // @[RegFile.scala 66:20:@46116.4]
  wire  regs_303_clock; // @[RegFile.scala 66:20:@46130.4]
  wire  regs_303_reset; // @[RegFile.scala 66:20:@46130.4]
  wire [63:0] regs_303_io_in; // @[RegFile.scala 66:20:@46130.4]
  wire  regs_303_io_reset; // @[RegFile.scala 66:20:@46130.4]
  wire [63:0] regs_303_io_out; // @[RegFile.scala 66:20:@46130.4]
  wire  regs_303_io_enable; // @[RegFile.scala 66:20:@46130.4]
  wire  regs_304_clock; // @[RegFile.scala 66:20:@46144.4]
  wire  regs_304_reset; // @[RegFile.scala 66:20:@46144.4]
  wire [63:0] regs_304_io_in; // @[RegFile.scala 66:20:@46144.4]
  wire  regs_304_io_reset; // @[RegFile.scala 66:20:@46144.4]
  wire [63:0] regs_304_io_out; // @[RegFile.scala 66:20:@46144.4]
  wire  regs_304_io_enable; // @[RegFile.scala 66:20:@46144.4]
  wire  regs_305_clock; // @[RegFile.scala 66:20:@46158.4]
  wire  regs_305_reset; // @[RegFile.scala 66:20:@46158.4]
  wire [63:0] regs_305_io_in; // @[RegFile.scala 66:20:@46158.4]
  wire  regs_305_io_reset; // @[RegFile.scala 66:20:@46158.4]
  wire [63:0] regs_305_io_out; // @[RegFile.scala 66:20:@46158.4]
  wire  regs_305_io_enable; // @[RegFile.scala 66:20:@46158.4]
  wire  regs_306_clock; // @[RegFile.scala 66:20:@46172.4]
  wire  regs_306_reset; // @[RegFile.scala 66:20:@46172.4]
  wire [63:0] regs_306_io_in; // @[RegFile.scala 66:20:@46172.4]
  wire  regs_306_io_reset; // @[RegFile.scala 66:20:@46172.4]
  wire [63:0] regs_306_io_out; // @[RegFile.scala 66:20:@46172.4]
  wire  regs_306_io_enable; // @[RegFile.scala 66:20:@46172.4]
  wire  regs_307_clock; // @[RegFile.scala 66:20:@46186.4]
  wire  regs_307_reset; // @[RegFile.scala 66:20:@46186.4]
  wire [63:0] regs_307_io_in; // @[RegFile.scala 66:20:@46186.4]
  wire  regs_307_io_reset; // @[RegFile.scala 66:20:@46186.4]
  wire [63:0] regs_307_io_out; // @[RegFile.scala 66:20:@46186.4]
  wire  regs_307_io_enable; // @[RegFile.scala 66:20:@46186.4]
  wire  regs_308_clock; // @[RegFile.scala 66:20:@46200.4]
  wire  regs_308_reset; // @[RegFile.scala 66:20:@46200.4]
  wire [63:0] regs_308_io_in; // @[RegFile.scala 66:20:@46200.4]
  wire  regs_308_io_reset; // @[RegFile.scala 66:20:@46200.4]
  wire [63:0] regs_308_io_out; // @[RegFile.scala 66:20:@46200.4]
  wire  regs_308_io_enable; // @[RegFile.scala 66:20:@46200.4]
  wire  regs_309_clock; // @[RegFile.scala 66:20:@46214.4]
  wire  regs_309_reset; // @[RegFile.scala 66:20:@46214.4]
  wire [63:0] regs_309_io_in; // @[RegFile.scala 66:20:@46214.4]
  wire  regs_309_io_reset; // @[RegFile.scala 66:20:@46214.4]
  wire [63:0] regs_309_io_out; // @[RegFile.scala 66:20:@46214.4]
  wire  regs_309_io_enable; // @[RegFile.scala 66:20:@46214.4]
  wire  regs_310_clock; // @[RegFile.scala 66:20:@46228.4]
  wire  regs_310_reset; // @[RegFile.scala 66:20:@46228.4]
  wire [63:0] regs_310_io_in; // @[RegFile.scala 66:20:@46228.4]
  wire  regs_310_io_reset; // @[RegFile.scala 66:20:@46228.4]
  wire [63:0] regs_310_io_out; // @[RegFile.scala 66:20:@46228.4]
  wire  regs_310_io_enable; // @[RegFile.scala 66:20:@46228.4]
  wire  regs_311_clock; // @[RegFile.scala 66:20:@46242.4]
  wire  regs_311_reset; // @[RegFile.scala 66:20:@46242.4]
  wire [63:0] regs_311_io_in; // @[RegFile.scala 66:20:@46242.4]
  wire  regs_311_io_reset; // @[RegFile.scala 66:20:@46242.4]
  wire [63:0] regs_311_io_out; // @[RegFile.scala 66:20:@46242.4]
  wire  regs_311_io_enable; // @[RegFile.scala 66:20:@46242.4]
  wire  regs_312_clock; // @[RegFile.scala 66:20:@46256.4]
  wire  regs_312_reset; // @[RegFile.scala 66:20:@46256.4]
  wire [63:0] regs_312_io_in; // @[RegFile.scala 66:20:@46256.4]
  wire  regs_312_io_reset; // @[RegFile.scala 66:20:@46256.4]
  wire [63:0] regs_312_io_out; // @[RegFile.scala 66:20:@46256.4]
  wire  regs_312_io_enable; // @[RegFile.scala 66:20:@46256.4]
  wire  regs_313_clock; // @[RegFile.scala 66:20:@46270.4]
  wire  regs_313_reset; // @[RegFile.scala 66:20:@46270.4]
  wire [63:0] regs_313_io_in; // @[RegFile.scala 66:20:@46270.4]
  wire  regs_313_io_reset; // @[RegFile.scala 66:20:@46270.4]
  wire [63:0] regs_313_io_out; // @[RegFile.scala 66:20:@46270.4]
  wire  regs_313_io_enable; // @[RegFile.scala 66:20:@46270.4]
  wire  regs_314_clock; // @[RegFile.scala 66:20:@46284.4]
  wire  regs_314_reset; // @[RegFile.scala 66:20:@46284.4]
  wire [63:0] regs_314_io_in; // @[RegFile.scala 66:20:@46284.4]
  wire  regs_314_io_reset; // @[RegFile.scala 66:20:@46284.4]
  wire [63:0] regs_314_io_out; // @[RegFile.scala 66:20:@46284.4]
  wire  regs_314_io_enable; // @[RegFile.scala 66:20:@46284.4]
  wire  regs_315_clock; // @[RegFile.scala 66:20:@46298.4]
  wire  regs_315_reset; // @[RegFile.scala 66:20:@46298.4]
  wire [63:0] regs_315_io_in; // @[RegFile.scala 66:20:@46298.4]
  wire  regs_315_io_reset; // @[RegFile.scala 66:20:@46298.4]
  wire [63:0] regs_315_io_out; // @[RegFile.scala 66:20:@46298.4]
  wire  regs_315_io_enable; // @[RegFile.scala 66:20:@46298.4]
  wire  regs_316_clock; // @[RegFile.scala 66:20:@46312.4]
  wire  regs_316_reset; // @[RegFile.scala 66:20:@46312.4]
  wire [63:0] regs_316_io_in; // @[RegFile.scala 66:20:@46312.4]
  wire  regs_316_io_reset; // @[RegFile.scala 66:20:@46312.4]
  wire [63:0] regs_316_io_out; // @[RegFile.scala 66:20:@46312.4]
  wire  regs_316_io_enable; // @[RegFile.scala 66:20:@46312.4]
  wire  regs_317_clock; // @[RegFile.scala 66:20:@46326.4]
  wire  regs_317_reset; // @[RegFile.scala 66:20:@46326.4]
  wire [63:0] regs_317_io_in; // @[RegFile.scala 66:20:@46326.4]
  wire  regs_317_io_reset; // @[RegFile.scala 66:20:@46326.4]
  wire [63:0] regs_317_io_out; // @[RegFile.scala 66:20:@46326.4]
  wire  regs_317_io_enable; // @[RegFile.scala 66:20:@46326.4]
  wire  regs_318_clock; // @[RegFile.scala 66:20:@46340.4]
  wire  regs_318_reset; // @[RegFile.scala 66:20:@46340.4]
  wire [63:0] regs_318_io_in; // @[RegFile.scala 66:20:@46340.4]
  wire  regs_318_io_reset; // @[RegFile.scala 66:20:@46340.4]
  wire [63:0] regs_318_io_out; // @[RegFile.scala 66:20:@46340.4]
  wire  regs_318_io_enable; // @[RegFile.scala 66:20:@46340.4]
  wire  regs_319_clock; // @[RegFile.scala 66:20:@46354.4]
  wire  regs_319_reset; // @[RegFile.scala 66:20:@46354.4]
  wire [63:0] regs_319_io_in; // @[RegFile.scala 66:20:@46354.4]
  wire  regs_319_io_reset; // @[RegFile.scala 66:20:@46354.4]
  wire [63:0] regs_319_io_out; // @[RegFile.scala 66:20:@46354.4]
  wire  regs_319_io_enable; // @[RegFile.scala 66:20:@46354.4]
  wire  regs_320_clock; // @[RegFile.scala 66:20:@46368.4]
  wire  regs_320_reset; // @[RegFile.scala 66:20:@46368.4]
  wire [63:0] regs_320_io_in; // @[RegFile.scala 66:20:@46368.4]
  wire  regs_320_io_reset; // @[RegFile.scala 66:20:@46368.4]
  wire [63:0] regs_320_io_out; // @[RegFile.scala 66:20:@46368.4]
  wire  regs_320_io_enable; // @[RegFile.scala 66:20:@46368.4]
  wire  regs_321_clock; // @[RegFile.scala 66:20:@46382.4]
  wire  regs_321_reset; // @[RegFile.scala 66:20:@46382.4]
  wire [63:0] regs_321_io_in; // @[RegFile.scala 66:20:@46382.4]
  wire  regs_321_io_reset; // @[RegFile.scala 66:20:@46382.4]
  wire [63:0] regs_321_io_out; // @[RegFile.scala 66:20:@46382.4]
  wire  regs_321_io_enable; // @[RegFile.scala 66:20:@46382.4]
  wire  regs_322_clock; // @[RegFile.scala 66:20:@46396.4]
  wire  regs_322_reset; // @[RegFile.scala 66:20:@46396.4]
  wire [63:0] regs_322_io_in; // @[RegFile.scala 66:20:@46396.4]
  wire  regs_322_io_reset; // @[RegFile.scala 66:20:@46396.4]
  wire [63:0] regs_322_io_out; // @[RegFile.scala 66:20:@46396.4]
  wire  regs_322_io_enable; // @[RegFile.scala 66:20:@46396.4]
  wire  regs_323_clock; // @[RegFile.scala 66:20:@46410.4]
  wire  regs_323_reset; // @[RegFile.scala 66:20:@46410.4]
  wire [63:0] regs_323_io_in; // @[RegFile.scala 66:20:@46410.4]
  wire  regs_323_io_reset; // @[RegFile.scala 66:20:@46410.4]
  wire [63:0] regs_323_io_out; // @[RegFile.scala 66:20:@46410.4]
  wire  regs_323_io_enable; // @[RegFile.scala 66:20:@46410.4]
  wire  regs_324_clock; // @[RegFile.scala 66:20:@46424.4]
  wire  regs_324_reset; // @[RegFile.scala 66:20:@46424.4]
  wire [63:0] regs_324_io_in; // @[RegFile.scala 66:20:@46424.4]
  wire  regs_324_io_reset; // @[RegFile.scala 66:20:@46424.4]
  wire [63:0] regs_324_io_out; // @[RegFile.scala 66:20:@46424.4]
  wire  regs_324_io_enable; // @[RegFile.scala 66:20:@46424.4]
  wire  regs_325_clock; // @[RegFile.scala 66:20:@46438.4]
  wire  regs_325_reset; // @[RegFile.scala 66:20:@46438.4]
  wire [63:0] regs_325_io_in; // @[RegFile.scala 66:20:@46438.4]
  wire  regs_325_io_reset; // @[RegFile.scala 66:20:@46438.4]
  wire [63:0] regs_325_io_out; // @[RegFile.scala 66:20:@46438.4]
  wire  regs_325_io_enable; // @[RegFile.scala 66:20:@46438.4]
  wire  regs_326_clock; // @[RegFile.scala 66:20:@46452.4]
  wire  regs_326_reset; // @[RegFile.scala 66:20:@46452.4]
  wire [63:0] regs_326_io_in; // @[RegFile.scala 66:20:@46452.4]
  wire  regs_326_io_reset; // @[RegFile.scala 66:20:@46452.4]
  wire [63:0] regs_326_io_out; // @[RegFile.scala 66:20:@46452.4]
  wire  regs_326_io_enable; // @[RegFile.scala 66:20:@46452.4]
  wire  regs_327_clock; // @[RegFile.scala 66:20:@46466.4]
  wire  regs_327_reset; // @[RegFile.scala 66:20:@46466.4]
  wire [63:0] regs_327_io_in; // @[RegFile.scala 66:20:@46466.4]
  wire  regs_327_io_reset; // @[RegFile.scala 66:20:@46466.4]
  wire [63:0] regs_327_io_out; // @[RegFile.scala 66:20:@46466.4]
  wire  regs_327_io_enable; // @[RegFile.scala 66:20:@46466.4]
  wire  regs_328_clock; // @[RegFile.scala 66:20:@46480.4]
  wire  regs_328_reset; // @[RegFile.scala 66:20:@46480.4]
  wire [63:0] regs_328_io_in; // @[RegFile.scala 66:20:@46480.4]
  wire  regs_328_io_reset; // @[RegFile.scala 66:20:@46480.4]
  wire [63:0] regs_328_io_out; // @[RegFile.scala 66:20:@46480.4]
  wire  regs_328_io_enable; // @[RegFile.scala 66:20:@46480.4]
  wire  regs_329_clock; // @[RegFile.scala 66:20:@46494.4]
  wire  regs_329_reset; // @[RegFile.scala 66:20:@46494.4]
  wire [63:0] regs_329_io_in; // @[RegFile.scala 66:20:@46494.4]
  wire  regs_329_io_reset; // @[RegFile.scala 66:20:@46494.4]
  wire [63:0] regs_329_io_out; // @[RegFile.scala 66:20:@46494.4]
  wire  regs_329_io_enable; // @[RegFile.scala 66:20:@46494.4]
  wire  regs_330_clock; // @[RegFile.scala 66:20:@46508.4]
  wire  regs_330_reset; // @[RegFile.scala 66:20:@46508.4]
  wire [63:0] regs_330_io_in; // @[RegFile.scala 66:20:@46508.4]
  wire  regs_330_io_reset; // @[RegFile.scala 66:20:@46508.4]
  wire [63:0] regs_330_io_out; // @[RegFile.scala 66:20:@46508.4]
  wire  regs_330_io_enable; // @[RegFile.scala 66:20:@46508.4]
  wire  regs_331_clock; // @[RegFile.scala 66:20:@46522.4]
  wire  regs_331_reset; // @[RegFile.scala 66:20:@46522.4]
  wire [63:0] regs_331_io_in; // @[RegFile.scala 66:20:@46522.4]
  wire  regs_331_io_reset; // @[RegFile.scala 66:20:@46522.4]
  wire [63:0] regs_331_io_out; // @[RegFile.scala 66:20:@46522.4]
  wire  regs_331_io_enable; // @[RegFile.scala 66:20:@46522.4]
  wire  regs_332_clock; // @[RegFile.scala 66:20:@46536.4]
  wire  regs_332_reset; // @[RegFile.scala 66:20:@46536.4]
  wire [63:0] regs_332_io_in; // @[RegFile.scala 66:20:@46536.4]
  wire  regs_332_io_reset; // @[RegFile.scala 66:20:@46536.4]
  wire [63:0] regs_332_io_out; // @[RegFile.scala 66:20:@46536.4]
  wire  regs_332_io_enable; // @[RegFile.scala 66:20:@46536.4]
  wire  regs_333_clock; // @[RegFile.scala 66:20:@46550.4]
  wire  regs_333_reset; // @[RegFile.scala 66:20:@46550.4]
  wire [63:0] regs_333_io_in; // @[RegFile.scala 66:20:@46550.4]
  wire  regs_333_io_reset; // @[RegFile.scala 66:20:@46550.4]
  wire [63:0] regs_333_io_out; // @[RegFile.scala 66:20:@46550.4]
  wire  regs_333_io_enable; // @[RegFile.scala 66:20:@46550.4]
  wire  regs_334_clock; // @[RegFile.scala 66:20:@46564.4]
  wire  regs_334_reset; // @[RegFile.scala 66:20:@46564.4]
  wire [63:0] regs_334_io_in; // @[RegFile.scala 66:20:@46564.4]
  wire  regs_334_io_reset; // @[RegFile.scala 66:20:@46564.4]
  wire [63:0] regs_334_io_out; // @[RegFile.scala 66:20:@46564.4]
  wire  regs_334_io_enable; // @[RegFile.scala 66:20:@46564.4]
  wire  regs_335_clock; // @[RegFile.scala 66:20:@46578.4]
  wire  regs_335_reset; // @[RegFile.scala 66:20:@46578.4]
  wire [63:0] regs_335_io_in; // @[RegFile.scala 66:20:@46578.4]
  wire  regs_335_io_reset; // @[RegFile.scala 66:20:@46578.4]
  wire [63:0] regs_335_io_out; // @[RegFile.scala 66:20:@46578.4]
  wire  regs_335_io_enable; // @[RegFile.scala 66:20:@46578.4]
  wire  regs_336_clock; // @[RegFile.scala 66:20:@46592.4]
  wire  regs_336_reset; // @[RegFile.scala 66:20:@46592.4]
  wire [63:0] regs_336_io_in; // @[RegFile.scala 66:20:@46592.4]
  wire  regs_336_io_reset; // @[RegFile.scala 66:20:@46592.4]
  wire [63:0] regs_336_io_out; // @[RegFile.scala 66:20:@46592.4]
  wire  regs_336_io_enable; // @[RegFile.scala 66:20:@46592.4]
  wire  regs_337_clock; // @[RegFile.scala 66:20:@46606.4]
  wire  regs_337_reset; // @[RegFile.scala 66:20:@46606.4]
  wire [63:0] regs_337_io_in; // @[RegFile.scala 66:20:@46606.4]
  wire  regs_337_io_reset; // @[RegFile.scala 66:20:@46606.4]
  wire [63:0] regs_337_io_out; // @[RegFile.scala 66:20:@46606.4]
  wire  regs_337_io_enable; // @[RegFile.scala 66:20:@46606.4]
  wire  regs_338_clock; // @[RegFile.scala 66:20:@46620.4]
  wire  regs_338_reset; // @[RegFile.scala 66:20:@46620.4]
  wire [63:0] regs_338_io_in; // @[RegFile.scala 66:20:@46620.4]
  wire  regs_338_io_reset; // @[RegFile.scala 66:20:@46620.4]
  wire [63:0] regs_338_io_out; // @[RegFile.scala 66:20:@46620.4]
  wire  regs_338_io_enable; // @[RegFile.scala 66:20:@46620.4]
  wire  regs_339_clock; // @[RegFile.scala 66:20:@46634.4]
  wire  regs_339_reset; // @[RegFile.scala 66:20:@46634.4]
  wire [63:0] regs_339_io_in; // @[RegFile.scala 66:20:@46634.4]
  wire  regs_339_io_reset; // @[RegFile.scala 66:20:@46634.4]
  wire [63:0] regs_339_io_out; // @[RegFile.scala 66:20:@46634.4]
  wire  regs_339_io_enable; // @[RegFile.scala 66:20:@46634.4]
  wire  regs_340_clock; // @[RegFile.scala 66:20:@46648.4]
  wire  regs_340_reset; // @[RegFile.scala 66:20:@46648.4]
  wire [63:0] regs_340_io_in; // @[RegFile.scala 66:20:@46648.4]
  wire  regs_340_io_reset; // @[RegFile.scala 66:20:@46648.4]
  wire [63:0] regs_340_io_out; // @[RegFile.scala 66:20:@46648.4]
  wire  regs_340_io_enable; // @[RegFile.scala 66:20:@46648.4]
  wire  regs_341_clock; // @[RegFile.scala 66:20:@46662.4]
  wire  regs_341_reset; // @[RegFile.scala 66:20:@46662.4]
  wire [63:0] regs_341_io_in; // @[RegFile.scala 66:20:@46662.4]
  wire  regs_341_io_reset; // @[RegFile.scala 66:20:@46662.4]
  wire [63:0] regs_341_io_out; // @[RegFile.scala 66:20:@46662.4]
  wire  regs_341_io_enable; // @[RegFile.scala 66:20:@46662.4]
  wire  regs_342_clock; // @[RegFile.scala 66:20:@46676.4]
  wire  regs_342_reset; // @[RegFile.scala 66:20:@46676.4]
  wire [63:0] regs_342_io_in; // @[RegFile.scala 66:20:@46676.4]
  wire  regs_342_io_reset; // @[RegFile.scala 66:20:@46676.4]
  wire [63:0] regs_342_io_out; // @[RegFile.scala 66:20:@46676.4]
  wire  regs_342_io_enable; // @[RegFile.scala 66:20:@46676.4]
  wire  regs_343_clock; // @[RegFile.scala 66:20:@46690.4]
  wire  regs_343_reset; // @[RegFile.scala 66:20:@46690.4]
  wire [63:0] regs_343_io_in; // @[RegFile.scala 66:20:@46690.4]
  wire  regs_343_io_reset; // @[RegFile.scala 66:20:@46690.4]
  wire [63:0] regs_343_io_out; // @[RegFile.scala 66:20:@46690.4]
  wire  regs_343_io_enable; // @[RegFile.scala 66:20:@46690.4]
  wire  regs_344_clock; // @[RegFile.scala 66:20:@46704.4]
  wire  regs_344_reset; // @[RegFile.scala 66:20:@46704.4]
  wire [63:0] regs_344_io_in; // @[RegFile.scala 66:20:@46704.4]
  wire  regs_344_io_reset; // @[RegFile.scala 66:20:@46704.4]
  wire [63:0] regs_344_io_out; // @[RegFile.scala 66:20:@46704.4]
  wire  regs_344_io_enable; // @[RegFile.scala 66:20:@46704.4]
  wire  regs_345_clock; // @[RegFile.scala 66:20:@46718.4]
  wire  regs_345_reset; // @[RegFile.scala 66:20:@46718.4]
  wire [63:0] regs_345_io_in; // @[RegFile.scala 66:20:@46718.4]
  wire  regs_345_io_reset; // @[RegFile.scala 66:20:@46718.4]
  wire [63:0] regs_345_io_out; // @[RegFile.scala 66:20:@46718.4]
  wire  regs_345_io_enable; // @[RegFile.scala 66:20:@46718.4]
  wire  regs_346_clock; // @[RegFile.scala 66:20:@46732.4]
  wire  regs_346_reset; // @[RegFile.scala 66:20:@46732.4]
  wire [63:0] regs_346_io_in; // @[RegFile.scala 66:20:@46732.4]
  wire  regs_346_io_reset; // @[RegFile.scala 66:20:@46732.4]
  wire [63:0] regs_346_io_out; // @[RegFile.scala 66:20:@46732.4]
  wire  regs_346_io_enable; // @[RegFile.scala 66:20:@46732.4]
  wire  regs_347_clock; // @[RegFile.scala 66:20:@46746.4]
  wire  regs_347_reset; // @[RegFile.scala 66:20:@46746.4]
  wire [63:0] regs_347_io_in; // @[RegFile.scala 66:20:@46746.4]
  wire  regs_347_io_reset; // @[RegFile.scala 66:20:@46746.4]
  wire [63:0] regs_347_io_out; // @[RegFile.scala 66:20:@46746.4]
  wire  regs_347_io_enable; // @[RegFile.scala 66:20:@46746.4]
  wire  regs_348_clock; // @[RegFile.scala 66:20:@46760.4]
  wire  regs_348_reset; // @[RegFile.scala 66:20:@46760.4]
  wire [63:0] regs_348_io_in; // @[RegFile.scala 66:20:@46760.4]
  wire  regs_348_io_reset; // @[RegFile.scala 66:20:@46760.4]
  wire [63:0] regs_348_io_out; // @[RegFile.scala 66:20:@46760.4]
  wire  regs_348_io_enable; // @[RegFile.scala 66:20:@46760.4]
  wire  regs_349_clock; // @[RegFile.scala 66:20:@46774.4]
  wire  regs_349_reset; // @[RegFile.scala 66:20:@46774.4]
  wire [63:0] regs_349_io_in; // @[RegFile.scala 66:20:@46774.4]
  wire  regs_349_io_reset; // @[RegFile.scala 66:20:@46774.4]
  wire [63:0] regs_349_io_out; // @[RegFile.scala 66:20:@46774.4]
  wire  regs_349_io_enable; // @[RegFile.scala 66:20:@46774.4]
  wire  regs_350_clock; // @[RegFile.scala 66:20:@46788.4]
  wire  regs_350_reset; // @[RegFile.scala 66:20:@46788.4]
  wire [63:0] regs_350_io_in; // @[RegFile.scala 66:20:@46788.4]
  wire  regs_350_io_reset; // @[RegFile.scala 66:20:@46788.4]
  wire [63:0] regs_350_io_out; // @[RegFile.scala 66:20:@46788.4]
  wire  regs_350_io_enable; // @[RegFile.scala 66:20:@46788.4]
  wire  regs_351_clock; // @[RegFile.scala 66:20:@46802.4]
  wire  regs_351_reset; // @[RegFile.scala 66:20:@46802.4]
  wire [63:0] regs_351_io_in; // @[RegFile.scala 66:20:@46802.4]
  wire  regs_351_io_reset; // @[RegFile.scala 66:20:@46802.4]
  wire [63:0] regs_351_io_out; // @[RegFile.scala 66:20:@46802.4]
  wire  regs_351_io_enable; // @[RegFile.scala 66:20:@46802.4]
  wire  regs_352_clock; // @[RegFile.scala 66:20:@46816.4]
  wire  regs_352_reset; // @[RegFile.scala 66:20:@46816.4]
  wire [63:0] regs_352_io_in; // @[RegFile.scala 66:20:@46816.4]
  wire  regs_352_io_reset; // @[RegFile.scala 66:20:@46816.4]
  wire [63:0] regs_352_io_out; // @[RegFile.scala 66:20:@46816.4]
  wire  regs_352_io_enable; // @[RegFile.scala 66:20:@46816.4]
  wire  regs_353_clock; // @[RegFile.scala 66:20:@46830.4]
  wire  regs_353_reset; // @[RegFile.scala 66:20:@46830.4]
  wire [63:0] regs_353_io_in; // @[RegFile.scala 66:20:@46830.4]
  wire  regs_353_io_reset; // @[RegFile.scala 66:20:@46830.4]
  wire [63:0] regs_353_io_out; // @[RegFile.scala 66:20:@46830.4]
  wire  regs_353_io_enable; // @[RegFile.scala 66:20:@46830.4]
  wire  regs_354_clock; // @[RegFile.scala 66:20:@46844.4]
  wire  regs_354_reset; // @[RegFile.scala 66:20:@46844.4]
  wire [63:0] regs_354_io_in; // @[RegFile.scala 66:20:@46844.4]
  wire  regs_354_io_reset; // @[RegFile.scala 66:20:@46844.4]
  wire [63:0] regs_354_io_out; // @[RegFile.scala 66:20:@46844.4]
  wire  regs_354_io_enable; // @[RegFile.scala 66:20:@46844.4]
  wire  regs_355_clock; // @[RegFile.scala 66:20:@46858.4]
  wire  regs_355_reset; // @[RegFile.scala 66:20:@46858.4]
  wire [63:0] regs_355_io_in; // @[RegFile.scala 66:20:@46858.4]
  wire  regs_355_io_reset; // @[RegFile.scala 66:20:@46858.4]
  wire [63:0] regs_355_io_out; // @[RegFile.scala 66:20:@46858.4]
  wire  regs_355_io_enable; // @[RegFile.scala 66:20:@46858.4]
  wire  regs_356_clock; // @[RegFile.scala 66:20:@46872.4]
  wire  regs_356_reset; // @[RegFile.scala 66:20:@46872.4]
  wire [63:0] regs_356_io_in; // @[RegFile.scala 66:20:@46872.4]
  wire  regs_356_io_reset; // @[RegFile.scala 66:20:@46872.4]
  wire [63:0] regs_356_io_out; // @[RegFile.scala 66:20:@46872.4]
  wire  regs_356_io_enable; // @[RegFile.scala 66:20:@46872.4]
  wire  regs_357_clock; // @[RegFile.scala 66:20:@46886.4]
  wire  regs_357_reset; // @[RegFile.scala 66:20:@46886.4]
  wire [63:0] regs_357_io_in; // @[RegFile.scala 66:20:@46886.4]
  wire  regs_357_io_reset; // @[RegFile.scala 66:20:@46886.4]
  wire [63:0] regs_357_io_out; // @[RegFile.scala 66:20:@46886.4]
  wire  regs_357_io_enable; // @[RegFile.scala 66:20:@46886.4]
  wire  regs_358_clock; // @[RegFile.scala 66:20:@46900.4]
  wire  regs_358_reset; // @[RegFile.scala 66:20:@46900.4]
  wire [63:0] regs_358_io_in; // @[RegFile.scala 66:20:@46900.4]
  wire  regs_358_io_reset; // @[RegFile.scala 66:20:@46900.4]
  wire [63:0] regs_358_io_out; // @[RegFile.scala 66:20:@46900.4]
  wire  regs_358_io_enable; // @[RegFile.scala 66:20:@46900.4]
  wire  regs_359_clock; // @[RegFile.scala 66:20:@46914.4]
  wire  regs_359_reset; // @[RegFile.scala 66:20:@46914.4]
  wire [63:0] regs_359_io_in; // @[RegFile.scala 66:20:@46914.4]
  wire  regs_359_io_reset; // @[RegFile.scala 66:20:@46914.4]
  wire [63:0] regs_359_io_out; // @[RegFile.scala 66:20:@46914.4]
  wire  regs_359_io_enable; // @[RegFile.scala 66:20:@46914.4]
  wire  regs_360_clock; // @[RegFile.scala 66:20:@46928.4]
  wire  regs_360_reset; // @[RegFile.scala 66:20:@46928.4]
  wire [63:0] regs_360_io_in; // @[RegFile.scala 66:20:@46928.4]
  wire  regs_360_io_reset; // @[RegFile.scala 66:20:@46928.4]
  wire [63:0] regs_360_io_out; // @[RegFile.scala 66:20:@46928.4]
  wire  regs_360_io_enable; // @[RegFile.scala 66:20:@46928.4]
  wire  regs_361_clock; // @[RegFile.scala 66:20:@46942.4]
  wire  regs_361_reset; // @[RegFile.scala 66:20:@46942.4]
  wire [63:0] regs_361_io_in; // @[RegFile.scala 66:20:@46942.4]
  wire  regs_361_io_reset; // @[RegFile.scala 66:20:@46942.4]
  wire [63:0] regs_361_io_out; // @[RegFile.scala 66:20:@46942.4]
  wire  regs_361_io_enable; // @[RegFile.scala 66:20:@46942.4]
  wire  regs_362_clock; // @[RegFile.scala 66:20:@46956.4]
  wire  regs_362_reset; // @[RegFile.scala 66:20:@46956.4]
  wire [63:0] regs_362_io_in; // @[RegFile.scala 66:20:@46956.4]
  wire  regs_362_io_reset; // @[RegFile.scala 66:20:@46956.4]
  wire [63:0] regs_362_io_out; // @[RegFile.scala 66:20:@46956.4]
  wire  regs_362_io_enable; // @[RegFile.scala 66:20:@46956.4]
  wire  regs_363_clock; // @[RegFile.scala 66:20:@46970.4]
  wire  regs_363_reset; // @[RegFile.scala 66:20:@46970.4]
  wire [63:0] regs_363_io_in; // @[RegFile.scala 66:20:@46970.4]
  wire  regs_363_io_reset; // @[RegFile.scala 66:20:@46970.4]
  wire [63:0] regs_363_io_out; // @[RegFile.scala 66:20:@46970.4]
  wire  regs_363_io_enable; // @[RegFile.scala 66:20:@46970.4]
  wire  regs_364_clock; // @[RegFile.scala 66:20:@46984.4]
  wire  regs_364_reset; // @[RegFile.scala 66:20:@46984.4]
  wire [63:0] regs_364_io_in; // @[RegFile.scala 66:20:@46984.4]
  wire  regs_364_io_reset; // @[RegFile.scala 66:20:@46984.4]
  wire [63:0] regs_364_io_out; // @[RegFile.scala 66:20:@46984.4]
  wire  regs_364_io_enable; // @[RegFile.scala 66:20:@46984.4]
  wire  regs_365_clock; // @[RegFile.scala 66:20:@46998.4]
  wire  regs_365_reset; // @[RegFile.scala 66:20:@46998.4]
  wire [63:0] regs_365_io_in; // @[RegFile.scala 66:20:@46998.4]
  wire  regs_365_io_reset; // @[RegFile.scala 66:20:@46998.4]
  wire [63:0] regs_365_io_out; // @[RegFile.scala 66:20:@46998.4]
  wire  regs_365_io_enable; // @[RegFile.scala 66:20:@46998.4]
  wire  regs_366_clock; // @[RegFile.scala 66:20:@47012.4]
  wire  regs_366_reset; // @[RegFile.scala 66:20:@47012.4]
  wire [63:0] regs_366_io_in; // @[RegFile.scala 66:20:@47012.4]
  wire  regs_366_io_reset; // @[RegFile.scala 66:20:@47012.4]
  wire [63:0] regs_366_io_out; // @[RegFile.scala 66:20:@47012.4]
  wire  regs_366_io_enable; // @[RegFile.scala 66:20:@47012.4]
  wire  regs_367_clock; // @[RegFile.scala 66:20:@47026.4]
  wire  regs_367_reset; // @[RegFile.scala 66:20:@47026.4]
  wire [63:0] regs_367_io_in; // @[RegFile.scala 66:20:@47026.4]
  wire  regs_367_io_reset; // @[RegFile.scala 66:20:@47026.4]
  wire [63:0] regs_367_io_out; // @[RegFile.scala 66:20:@47026.4]
  wire  regs_367_io_enable; // @[RegFile.scala 66:20:@47026.4]
  wire  regs_368_clock; // @[RegFile.scala 66:20:@47040.4]
  wire  regs_368_reset; // @[RegFile.scala 66:20:@47040.4]
  wire [63:0] regs_368_io_in; // @[RegFile.scala 66:20:@47040.4]
  wire  regs_368_io_reset; // @[RegFile.scala 66:20:@47040.4]
  wire [63:0] regs_368_io_out; // @[RegFile.scala 66:20:@47040.4]
  wire  regs_368_io_enable; // @[RegFile.scala 66:20:@47040.4]
  wire  regs_369_clock; // @[RegFile.scala 66:20:@47054.4]
  wire  regs_369_reset; // @[RegFile.scala 66:20:@47054.4]
  wire [63:0] regs_369_io_in; // @[RegFile.scala 66:20:@47054.4]
  wire  regs_369_io_reset; // @[RegFile.scala 66:20:@47054.4]
  wire [63:0] regs_369_io_out; // @[RegFile.scala 66:20:@47054.4]
  wire  regs_369_io_enable; // @[RegFile.scala 66:20:@47054.4]
  wire  regs_370_clock; // @[RegFile.scala 66:20:@47068.4]
  wire  regs_370_reset; // @[RegFile.scala 66:20:@47068.4]
  wire [63:0] regs_370_io_in; // @[RegFile.scala 66:20:@47068.4]
  wire  regs_370_io_reset; // @[RegFile.scala 66:20:@47068.4]
  wire [63:0] regs_370_io_out; // @[RegFile.scala 66:20:@47068.4]
  wire  regs_370_io_enable; // @[RegFile.scala 66:20:@47068.4]
  wire  regs_371_clock; // @[RegFile.scala 66:20:@47082.4]
  wire  regs_371_reset; // @[RegFile.scala 66:20:@47082.4]
  wire [63:0] regs_371_io_in; // @[RegFile.scala 66:20:@47082.4]
  wire  regs_371_io_reset; // @[RegFile.scala 66:20:@47082.4]
  wire [63:0] regs_371_io_out; // @[RegFile.scala 66:20:@47082.4]
  wire  regs_371_io_enable; // @[RegFile.scala 66:20:@47082.4]
  wire  regs_372_clock; // @[RegFile.scala 66:20:@47096.4]
  wire  regs_372_reset; // @[RegFile.scala 66:20:@47096.4]
  wire [63:0] regs_372_io_in; // @[RegFile.scala 66:20:@47096.4]
  wire  regs_372_io_reset; // @[RegFile.scala 66:20:@47096.4]
  wire [63:0] regs_372_io_out; // @[RegFile.scala 66:20:@47096.4]
  wire  regs_372_io_enable; // @[RegFile.scala 66:20:@47096.4]
  wire  regs_373_clock; // @[RegFile.scala 66:20:@47110.4]
  wire  regs_373_reset; // @[RegFile.scala 66:20:@47110.4]
  wire [63:0] regs_373_io_in; // @[RegFile.scala 66:20:@47110.4]
  wire  regs_373_io_reset; // @[RegFile.scala 66:20:@47110.4]
  wire [63:0] regs_373_io_out; // @[RegFile.scala 66:20:@47110.4]
  wire  regs_373_io_enable; // @[RegFile.scala 66:20:@47110.4]
  wire  regs_374_clock; // @[RegFile.scala 66:20:@47124.4]
  wire  regs_374_reset; // @[RegFile.scala 66:20:@47124.4]
  wire [63:0] regs_374_io_in; // @[RegFile.scala 66:20:@47124.4]
  wire  regs_374_io_reset; // @[RegFile.scala 66:20:@47124.4]
  wire [63:0] regs_374_io_out; // @[RegFile.scala 66:20:@47124.4]
  wire  regs_374_io_enable; // @[RegFile.scala 66:20:@47124.4]
  wire  regs_375_clock; // @[RegFile.scala 66:20:@47138.4]
  wire  regs_375_reset; // @[RegFile.scala 66:20:@47138.4]
  wire [63:0] regs_375_io_in; // @[RegFile.scala 66:20:@47138.4]
  wire  regs_375_io_reset; // @[RegFile.scala 66:20:@47138.4]
  wire [63:0] regs_375_io_out; // @[RegFile.scala 66:20:@47138.4]
  wire  regs_375_io_enable; // @[RegFile.scala 66:20:@47138.4]
  wire  regs_376_clock; // @[RegFile.scala 66:20:@47152.4]
  wire  regs_376_reset; // @[RegFile.scala 66:20:@47152.4]
  wire [63:0] regs_376_io_in; // @[RegFile.scala 66:20:@47152.4]
  wire  regs_376_io_reset; // @[RegFile.scala 66:20:@47152.4]
  wire [63:0] regs_376_io_out; // @[RegFile.scala 66:20:@47152.4]
  wire  regs_376_io_enable; // @[RegFile.scala 66:20:@47152.4]
  wire  regs_377_clock; // @[RegFile.scala 66:20:@47166.4]
  wire  regs_377_reset; // @[RegFile.scala 66:20:@47166.4]
  wire [63:0] regs_377_io_in; // @[RegFile.scala 66:20:@47166.4]
  wire  regs_377_io_reset; // @[RegFile.scala 66:20:@47166.4]
  wire [63:0] regs_377_io_out; // @[RegFile.scala 66:20:@47166.4]
  wire  regs_377_io_enable; // @[RegFile.scala 66:20:@47166.4]
  wire  regs_378_clock; // @[RegFile.scala 66:20:@47180.4]
  wire  regs_378_reset; // @[RegFile.scala 66:20:@47180.4]
  wire [63:0] regs_378_io_in; // @[RegFile.scala 66:20:@47180.4]
  wire  regs_378_io_reset; // @[RegFile.scala 66:20:@47180.4]
  wire [63:0] regs_378_io_out; // @[RegFile.scala 66:20:@47180.4]
  wire  regs_378_io_enable; // @[RegFile.scala 66:20:@47180.4]
  wire  regs_379_clock; // @[RegFile.scala 66:20:@47194.4]
  wire  regs_379_reset; // @[RegFile.scala 66:20:@47194.4]
  wire [63:0] regs_379_io_in; // @[RegFile.scala 66:20:@47194.4]
  wire  regs_379_io_reset; // @[RegFile.scala 66:20:@47194.4]
  wire [63:0] regs_379_io_out; // @[RegFile.scala 66:20:@47194.4]
  wire  regs_379_io_enable; // @[RegFile.scala 66:20:@47194.4]
  wire  regs_380_clock; // @[RegFile.scala 66:20:@47208.4]
  wire  regs_380_reset; // @[RegFile.scala 66:20:@47208.4]
  wire [63:0] regs_380_io_in; // @[RegFile.scala 66:20:@47208.4]
  wire  regs_380_io_reset; // @[RegFile.scala 66:20:@47208.4]
  wire [63:0] regs_380_io_out; // @[RegFile.scala 66:20:@47208.4]
  wire  regs_380_io_enable; // @[RegFile.scala 66:20:@47208.4]
  wire  regs_381_clock; // @[RegFile.scala 66:20:@47222.4]
  wire  regs_381_reset; // @[RegFile.scala 66:20:@47222.4]
  wire [63:0] regs_381_io_in; // @[RegFile.scala 66:20:@47222.4]
  wire  regs_381_io_reset; // @[RegFile.scala 66:20:@47222.4]
  wire [63:0] regs_381_io_out; // @[RegFile.scala 66:20:@47222.4]
  wire  regs_381_io_enable; // @[RegFile.scala 66:20:@47222.4]
  wire  regs_382_clock; // @[RegFile.scala 66:20:@47236.4]
  wire  regs_382_reset; // @[RegFile.scala 66:20:@47236.4]
  wire [63:0] regs_382_io_in; // @[RegFile.scala 66:20:@47236.4]
  wire  regs_382_io_reset; // @[RegFile.scala 66:20:@47236.4]
  wire [63:0] regs_382_io_out; // @[RegFile.scala 66:20:@47236.4]
  wire  regs_382_io_enable; // @[RegFile.scala 66:20:@47236.4]
  wire  regs_383_clock; // @[RegFile.scala 66:20:@47250.4]
  wire  regs_383_reset; // @[RegFile.scala 66:20:@47250.4]
  wire [63:0] regs_383_io_in; // @[RegFile.scala 66:20:@47250.4]
  wire  regs_383_io_reset; // @[RegFile.scala 66:20:@47250.4]
  wire [63:0] regs_383_io_out; // @[RegFile.scala 66:20:@47250.4]
  wire  regs_383_io_enable; // @[RegFile.scala 66:20:@47250.4]
  wire  regs_384_clock; // @[RegFile.scala 66:20:@47264.4]
  wire  regs_384_reset; // @[RegFile.scala 66:20:@47264.4]
  wire [63:0] regs_384_io_in; // @[RegFile.scala 66:20:@47264.4]
  wire  regs_384_io_reset; // @[RegFile.scala 66:20:@47264.4]
  wire [63:0] regs_384_io_out; // @[RegFile.scala 66:20:@47264.4]
  wire  regs_384_io_enable; // @[RegFile.scala 66:20:@47264.4]
  wire  regs_385_clock; // @[RegFile.scala 66:20:@47278.4]
  wire  regs_385_reset; // @[RegFile.scala 66:20:@47278.4]
  wire [63:0] regs_385_io_in; // @[RegFile.scala 66:20:@47278.4]
  wire  regs_385_io_reset; // @[RegFile.scala 66:20:@47278.4]
  wire [63:0] regs_385_io_out; // @[RegFile.scala 66:20:@47278.4]
  wire  regs_385_io_enable; // @[RegFile.scala 66:20:@47278.4]
  wire  regs_386_clock; // @[RegFile.scala 66:20:@47292.4]
  wire  regs_386_reset; // @[RegFile.scala 66:20:@47292.4]
  wire [63:0] regs_386_io_in; // @[RegFile.scala 66:20:@47292.4]
  wire  regs_386_io_reset; // @[RegFile.scala 66:20:@47292.4]
  wire [63:0] regs_386_io_out; // @[RegFile.scala 66:20:@47292.4]
  wire  regs_386_io_enable; // @[RegFile.scala 66:20:@47292.4]
  wire  regs_387_clock; // @[RegFile.scala 66:20:@47306.4]
  wire  regs_387_reset; // @[RegFile.scala 66:20:@47306.4]
  wire [63:0] regs_387_io_in; // @[RegFile.scala 66:20:@47306.4]
  wire  regs_387_io_reset; // @[RegFile.scala 66:20:@47306.4]
  wire [63:0] regs_387_io_out; // @[RegFile.scala 66:20:@47306.4]
  wire  regs_387_io_enable; // @[RegFile.scala 66:20:@47306.4]
  wire  regs_388_clock; // @[RegFile.scala 66:20:@47320.4]
  wire  regs_388_reset; // @[RegFile.scala 66:20:@47320.4]
  wire [63:0] regs_388_io_in; // @[RegFile.scala 66:20:@47320.4]
  wire  regs_388_io_reset; // @[RegFile.scala 66:20:@47320.4]
  wire [63:0] regs_388_io_out; // @[RegFile.scala 66:20:@47320.4]
  wire  regs_388_io_enable; // @[RegFile.scala 66:20:@47320.4]
  wire  regs_389_clock; // @[RegFile.scala 66:20:@47334.4]
  wire  regs_389_reset; // @[RegFile.scala 66:20:@47334.4]
  wire [63:0] regs_389_io_in; // @[RegFile.scala 66:20:@47334.4]
  wire  regs_389_io_reset; // @[RegFile.scala 66:20:@47334.4]
  wire [63:0] regs_389_io_out; // @[RegFile.scala 66:20:@47334.4]
  wire  regs_389_io_enable; // @[RegFile.scala 66:20:@47334.4]
  wire  regs_390_clock; // @[RegFile.scala 66:20:@47348.4]
  wire  regs_390_reset; // @[RegFile.scala 66:20:@47348.4]
  wire [63:0] regs_390_io_in; // @[RegFile.scala 66:20:@47348.4]
  wire  regs_390_io_reset; // @[RegFile.scala 66:20:@47348.4]
  wire [63:0] regs_390_io_out; // @[RegFile.scala 66:20:@47348.4]
  wire  regs_390_io_enable; // @[RegFile.scala 66:20:@47348.4]
  wire  regs_391_clock; // @[RegFile.scala 66:20:@47362.4]
  wire  regs_391_reset; // @[RegFile.scala 66:20:@47362.4]
  wire [63:0] regs_391_io_in; // @[RegFile.scala 66:20:@47362.4]
  wire  regs_391_io_reset; // @[RegFile.scala 66:20:@47362.4]
  wire [63:0] regs_391_io_out; // @[RegFile.scala 66:20:@47362.4]
  wire  regs_391_io_enable; // @[RegFile.scala 66:20:@47362.4]
  wire  regs_392_clock; // @[RegFile.scala 66:20:@47376.4]
  wire  regs_392_reset; // @[RegFile.scala 66:20:@47376.4]
  wire [63:0] regs_392_io_in; // @[RegFile.scala 66:20:@47376.4]
  wire  regs_392_io_reset; // @[RegFile.scala 66:20:@47376.4]
  wire [63:0] regs_392_io_out; // @[RegFile.scala 66:20:@47376.4]
  wire  regs_392_io_enable; // @[RegFile.scala 66:20:@47376.4]
  wire  regs_393_clock; // @[RegFile.scala 66:20:@47390.4]
  wire  regs_393_reset; // @[RegFile.scala 66:20:@47390.4]
  wire [63:0] regs_393_io_in; // @[RegFile.scala 66:20:@47390.4]
  wire  regs_393_io_reset; // @[RegFile.scala 66:20:@47390.4]
  wire [63:0] regs_393_io_out; // @[RegFile.scala 66:20:@47390.4]
  wire  regs_393_io_enable; // @[RegFile.scala 66:20:@47390.4]
  wire  regs_394_clock; // @[RegFile.scala 66:20:@47404.4]
  wire  regs_394_reset; // @[RegFile.scala 66:20:@47404.4]
  wire [63:0] regs_394_io_in; // @[RegFile.scala 66:20:@47404.4]
  wire  regs_394_io_reset; // @[RegFile.scala 66:20:@47404.4]
  wire [63:0] regs_394_io_out; // @[RegFile.scala 66:20:@47404.4]
  wire  regs_394_io_enable; // @[RegFile.scala 66:20:@47404.4]
  wire  regs_395_clock; // @[RegFile.scala 66:20:@47418.4]
  wire  regs_395_reset; // @[RegFile.scala 66:20:@47418.4]
  wire [63:0] regs_395_io_in; // @[RegFile.scala 66:20:@47418.4]
  wire  regs_395_io_reset; // @[RegFile.scala 66:20:@47418.4]
  wire [63:0] regs_395_io_out; // @[RegFile.scala 66:20:@47418.4]
  wire  regs_395_io_enable; // @[RegFile.scala 66:20:@47418.4]
  wire  regs_396_clock; // @[RegFile.scala 66:20:@47432.4]
  wire  regs_396_reset; // @[RegFile.scala 66:20:@47432.4]
  wire [63:0] regs_396_io_in; // @[RegFile.scala 66:20:@47432.4]
  wire  regs_396_io_reset; // @[RegFile.scala 66:20:@47432.4]
  wire [63:0] regs_396_io_out; // @[RegFile.scala 66:20:@47432.4]
  wire  regs_396_io_enable; // @[RegFile.scala 66:20:@47432.4]
  wire  regs_397_clock; // @[RegFile.scala 66:20:@47446.4]
  wire  regs_397_reset; // @[RegFile.scala 66:20:@47446.4]
  wire [63:0] regs_397_io_in; // @[RegFile.scala 66:20:@47446.4]
  wire  regs_397_io_reset; // @[RegFile.scala 66:20:@47446.4]
  wire [63:0] regs_397_io_out; // @[RegFile.scala 66:20:@47446.4]
  wire  regs_397_io_enable; // @[RegFile.scala 66:20:@47446.4]
  wire  regs_398_clock; // @[RegFile.scala 66:20:@47460.4]
  wire  regs_398_reset; // @[RegFile.scala 66:20:@47460.4]
  wire [63:0] regs_398_io_in; // @[RegFile.scala 66:20:@47460.4]
  wire  regs_398_io_reset; // @[RegFile.scala 66:20:@47460.4]
  wire [63:0] regs_398_io_out; // @[RegFile.scala 66:20:@47460.4]
  wire  regs_398_io_enable; // @[RegFile.scala 66:20:@47460.4]
  wire  regs_399_clock; // @[RegFile.scala 66:20:@47474.4]
  wire  regs_399_reset; // @[RegFile.scala 66:20:@47474.4]
  wire [63:0] regs_399_io_in; // @[RegFile.scala 66:20:@47474.4]
  wire  regs_399_io_reset; // @[RegFile.scala 66:20:@47474.4]
  wire [63:0] regs_399_io_out; // @[RegFile.scala 66:20:@47474.4]
  wire  regs_399_io_enable; // @[RegFile.scala 66:20:@47474.4]
  wire  regs_400_clock; // @[RegFile.scala 66:20:@47488.4]
  wire  regs_400_reset; // @[RegFile.scala 66:20:@47488.4]
  wire [63:0] regs_400_io_in; // @[RegFile.scala 66:20:@47488.4]
  wire  regs_400_io_reset; // @[RegFile.scala 66:20:@47488.4]
  wire [63:0] regs_400_io_out; // @[RegFile.scala 66:20:@47488.4]
  wire  regs_400_io_enable; // @[RegFile.scala 66:20:@47488.4]
  wire  regs_401_clock; // @[RegFile.scala 66:20:@47502.4]
  wire  regs_401_reset; // @[RegFile.scala 66:20:@47502.4]
  wire [63:0] regs_401_io_in; // @[RegFile.scala 66:20:@47502.4]
  wire  regs_401_io_reset; // @[RegFile.scala 66:20:@47502.4]
  wire [63:0] regs_401_io_out; // @[RegFile.scala 66:20:@47502.4]
  wire  regs_401_io_enable; // @[RegFile.scala 66:20:@47502.4]
  wire  regs_402_clock; // @[RegFile.scala 66:20:@47516.4]
  wire  regs_402_reset; // @[RegFile.scala 66:20:@47516.4]
  wire [63:0] regs_402_io_in; // @[RegFile.scala 66:20:@47516.4]
  wire  regs_402_io_reset; // @[RegFile.scala 66:20:@47516.4]
  wire [63:0] regs_402_io_out; // @[RegFile.scala 66:20:@47516.4]
  wire  regs_402_io_enable; // @[RegFile.scala 66:20:@47516.4]
  wire  regs_403_clock; // @[RegFile.scala 66:20:@47530.4]
  wire  regs_403_reset; // @[RegFile.scala 66:20:@47530.4]
  wire [63:0] regs_403_io_in; // @[RegFile.scala 66:20:@47530.4]
  wire  regs_403_io_reset; // @[RegFile.scala 66:20:@47530.4]
  wire [63:0] regs_403_io_out; // @[RegFile.scala 66:20:@47530.4]
  wire  regs_403_io_enable; // @[RegFile.scala 66:20:@47530.4]
  wire  regs_404_clock; // @[RegFile.scala 66:20:@47544.4]
  wire  regs_404_reset; // @[RegFile.scala 66:20:@47544.4]
  wire [63:0] regs_404_io_in; // @[RegFile.scala 66:20:@47544.4]
  wire  regs_404_io_reset; // @[RegFile.scala 66:20:@47544.4]
  wire [63:0] regs_404_io_out; // @[RegFile.scala 66:20:@47544.4]
  wire  regs_404_io_enable; // @[RegFile.scala 66:20:@47544.4]
  wire  regs_405_clock; // @[RegFile.scala 66:20:@47558.4]
  wire  regs_405_reset; // @[RegFile.scala 66:20:@47558.4]
  wire [63:0] regs_405_io_in; // @[RegFile.scala 66:20:@47558.4]
  wire  regs_405_io_reset; // @[RegFile.scala 66:20:@47558.4]
  wire [63:0] regs_405_io_out; // @[RegFile.scala 66:20:@47558.4]
  wire  regs_405_io_enable; // @[RegFile.scala 66:20:@47558.4]
  wire  regs_406_clock; // @[RegFile.scala 66:20:@47572.4]
  wire  regs_406_reset; // @[RegFile.scala 66:20:@47572.4]
  wire [63:0] regs_406_io_in; // @[RegFile.scala 66:20:@47572.4]
  wire  regs_406_io_reset; // @[RegFile.scala 66:20:@47572.4]
  wire [63:0] regs_406_io_out; // @[RegFile.scala 66:20:@47572.4]
  wire  regs_406_io_enable; // @[RegFile.scala 66:20:@47572.4]
  wire  regs_407_clock; // @[RegFile.scala 66:20:@47586.4]
  wire  regs_407_reset; // @[RegFile.scala 66:20:@47586.4]
  wire [63:0] regs_407_io_in; // @[RegFile.scala 66:20:@47586.4]
  wire  regs_407_io_reset; // @[RegFile.scala 66:20:@47586.4]
  wire [63:0] regs_407_io_out; // @[RegFile.scala 66:20:@47586.4]
  wire  regs_407_io_enable; // @[RegFile.scala 66:20:@47586.4]
  wire  regs_408_clock; // @[RegFile.scala 66:20:@47600.4]
  wire  regs_408_reset; // @[RegFile.scala 66:20:@47600.4]
  wire [63:0] regs_408_io_in; // @[RegFile.scala 66:20:@47600.4]
  wire  regs_408_io_reset; // @[RegFile.scala 66:20:@47600.4]
  wire [63:0] regs_408_io_out; // @[RegFile.scala 66:20:@47600.4]
  wire  regs_408_io_enable; // @[RegFile.scala 66:20:@47600.4]
  wire  regs_409_clock; // @[RegFile.scala 66:20:@47614.4]
  wire  regs_409_reset; // @[RegFile.scala 66:20:@47614.4]
  wire [63:0] regs_409_io_in; // @[RegFile.scala 66:20:@47614.4]
  wire  regs_409_io_reset; // @[RegFile.scala 66:20:@47614.4]
  wire [63:0] regs_409_io_out; // @[RegFile.scala 66:20:@47614.4]
  wire  regs_409_io_enable; // @[RegFile.scala 66:20:@47614.4]
  wire  regs_410_clock; // @[RegFile.scala 66:20:@47628.4]
  wire  regs_410_reset; // @[RegFile.scala 66:20:@47628.4]
  wire [63:0] regs_410_io_in; // @[RegFile.scala 66:20:@47628.4]
  wire  regs_410_io_reset; // @[RegFile.scala 66:20:@47628.4]
  wire [63:0] regs_410_io_out; // @[RegFile.scala 66:20:@47628.4]
  wire  regs_410_io_enable; // @[RegFile.scala 66:20:@47628.4]
  wire  regs_411_clock; // @[RegFile.scala 66:20:@47642.4]
  wire  regs_411_reset; // @[RegFile.scala 66:20:@47642.4]
  wire [63:0] regs_411_io_in; // @[RegFile.scala 66:20:@47642.4]
  wire  regs_411_io_reset; // @[RegFile.scala 66:20:@47642.4]
  wire [63:0] regs_411_io_out; // @[RegFile.scala 66:20:@47642.4]
  wire  regs_411_io_enable; // @[RegFile.scala 66:20:@47642.4]
  wire  regs_412_clock; // @[RegFile.scala 66:20:@47656.4]
  wire  regs_412_reset; // @[RegFile.scala 66:20:@47656.4]
  wire [63:0] regs_412_io_in; // @[RegFile.scala 66:20:@47656.4]
  wire  regs_412_io_reset; // @[RegFile.scala 66:20:@47656.4]
  wire [63:0] regs_412_io_out; // @[RegFile.scala 66:20:@47656.4]
  wire  regs_412_io_enable; // @[RegFile.scala 66:20:@47656.4]
  wire  regs_413_clock; // @[RegFile.scala 66:20:@47670.4]
  wire  regs_413_reset; // @[RegFile.scala 66:20:@47670.4]
  wire [63:0] regs_413_io_in; // @[RegFile.scala 66:20:@47670.4]
  wire  regs_413_io_reset; // @[RegFile.scala 66:20:@47670.4]
  wire [63:0] regs_413_io_out; // @[RegFile.scala 66:20:@47670.4]
  wire  regs_413_io_enable; // @[RegFile.scala 66:20:@47670.4]
  wire  regs_414_clock; // @[RegFile.scala 66:20:@47684.4]
  wire  regs_414_reset; // @[RegFile.scala 66:20:@47684.4]
  wire [63:0] regs_414_io_in; // @[RegFile.scala 66:20:@47684.4]
  wire  regs_414_io_reset; // @[RegFile.scala 66:20:@47684.4]
  wire [63:0] regs_414_io_out; // @[RegFile.scala 66:20:@47684.4]
  wire  regs_414_io_enable; // @[RegFile.scala 66:20:@47684.4]
  wire  regs_415_clock; // @[RegFile.scala 66:20:@47698.4]
  wire  regs_415_reset; // @[RegFile.scala 66:20:@47698.4]
  wire [63:0] regs_415_io_in; // @[RegFile.scala 66:20:@47698.4]
  wire  regs_415_io_reset; // @[RegFile.scala 66:20:@47698.4]
  wire [63:0] regs_415_io_out; // @[RegFile.scala 66:20:@47698.4]
  wire  regs_415_io_enable; // @[RegFile.scala 66:20:@47698.4]
  wire  regs_416_clock; // @[RegFile.scala 66:20:@47712.4]
  wire  regs_416_reset; // @[RegFile.scala 66:20:@47712.4]
  wire [63:0] regs_416_io_in; // @[RegFile.scala 66:20:@47712.4]
  wire  regs_416_io_reset; // @[RegFile.scala 66:20:@47712.4]
  wire [63:0] regs_416_io_out; // @[RegFile.scala 66:20:@47712.4]
  wire  regs_416_io_enable; // @[RegFile.scala 66:20:@47712.4]
  wire  regs_417_clock; // @[RegFile.scala 66:20:@47726.4]
  wire  regs_417_reset; // @[RegFile.scala 66:20:@47726.4]
  wire [63:0] regs_417_io_in; // @[RegFile.scala 66:20:@47726.4]
  wire  regs_417_io_reset; // @[RegFile.scala 66:20:@47726.4]
  wire [63:0] regs_417_io_out; // @[RegFile.scala 66:20:@47726.4]
  wire  regs_417_io_enable; // @[RegFile.scala 66:20:@47726.4]
  wire  regs_418_clock; // @[RegFile.scala 66:20:@47740.4]
  wire  regs_418_reset; // @[RegFile.scala 66:20:@47740.4]
  wire [63:0] regs_418_io_in; // @[RegFile.scala 66:20:@47740.4]
  wire  regs_418_io_reset; // @[RegFile.scala 66:20:@47740.4]
  wire [63:0] regs_418_io_out; // @[RegFile.scala 66:20:@47740.4]
  wire  regs_418_io_enable; // @[RegFile.scala 66:20:@47740.4]
  wire  regs_419_clock; // @[RegFile.scala 66:20:@47754.4]
  wire  regs_419_reset; // @[RegFile.scala 66:20:@47754.4]
  wire [63:0] regs_419_io_in; // @[RegFile.scala 66:20:@47754.4]
  wire  regs_419_io_reset; // @[RegFile.scala 66:20:@47754.4]
  wire [63:0] regs_419_io_out; // @[RegFile.scala 66:20:@47754.4]
  wire  regs_419_io_enable; // @[RegFile.scala 66:20:@47754.4]
  wire  regs_420_clock; // @[RegFile.scala 66:20:@47768.4]
  wire  regs_420_reset; // @[RegFile.scala 66:20:@47768.4]
  wire [63:0] regs_420_io_in; // @[RegFile.scala 66:20:@47768.4]
  wire  regs_420_io_reset; // @[RegFile.scala 66:20:@47768.4]
  wire [63:0] regs_420_io_out; // @[RegFile.scala 66:20:@47768.4]
  wire  regs_420_io_enable; // @[RegFile.scala 66:20:@47768.4]
  wire  regs_421_clock; // @[RegFile.scala 66:20:@47782.4]
  wire  regs_421_reset; // @[RegFile.scala 66:20:@47782.4]
  wire [63:0] regs_421_io_in; // @[RegFile.scala 66:20:@47782.4]
  wire  regs_421_io_reset; // @[RegFile.scala 66:20:@47782.4]
  wire [63:0] regs_421_io_out; // @[RegFile.scala 66:20:@47782.4]
  wire  regs_421_io_enable; // @[RegFile.scala 66:20:@47782.4]
  wire  regs_422_clock; // @[RegFile.scala 66:20:@47796.4]
  wire  regs_422_reset; // @[RegFile.scala 66:20:@47796.4]
  wire [63:0] regs_422_io_in; // @[RegFile.scala 66:20:@47796.4]
  wire  regs_422_io_reset; // @[RegFile.scala 66:20:@47796.4]
  wire [63:0] regs_422_io_out; // @[RegFile.scala 66:20:@47796.4]
  wire  regs_422_io_enable; // @[RegFile.scala 66:20:@47796.4]
  wire  regs_423_clock; // @[RegFile.scala 66:20:@47810.4]
  wire  regs_423_reset; // @[RegFile.scala 66:20:@47810.4]
  wire [63:0] regs_423_io_in; // @[RegFile.scala 66:20:@47810.4]
  wire  regs_423_io_reset; // @[RegFile.scala 66:20:@47810.4]
  wire [63:0] regs_423_io_out; // @[RegFile.scala 66:20:@47810.4]
  wire  regs_423_io_enable; // @[RegFile.scala 66:20:@47810.4]
  wire  regs_424_clock; // @[RegFile.scala 66:20:@47824.4]
  wire  regs_424_reset; // @[RegFile.scala 66:20:@47824.4]
  wire [63:0] regs_424_io_in; // @[RegFile.scala 66:20:@47824.4]
  wire  regs_424_io_reset; // @[RegFile.scala 66:20:@47824.4]
  wire [63:0] regs_424_io_out; // @[RegFile.scala 66:20:@47824.4]
  wire  regs_424_io_enable; // @[RegFile.scala 66:20:@47824.4]
  wire  regs_425_clock; // @[RegFile.scala 66:20:@47838.4]
  wire  regs_425_reset; // @[RegFile.scala 66:20:@47838.4]
  wire [63:0] regs_425_io_in; // @[RegFile.scala 66:20:@47838.4]
  wire  regs_425_io_reset; // @[RegFile.scala 66:20:@47838.4]
  wire [63:0] regs_425_io_out; // @[RegFile.scala 66:20:@47838.4]
  wire  regs_425_io_enable; // @[RegFile.scala 66:20:@47838.4]
  wire  regs_426_clock; // @[RegFile.scala 66:20:@47852.4]
  wire  regs_426_reset; // @[RegFile.scala 66:20:@47852.4]
  wire [63:0] regs_426_io_in; // @[RegFile.scala 66:20:@47852.4]
  wire  regs_426_io_reset; // @[RegFile.scala 66:20:@47852.4]
  wire [63:0] regs_426_io_out; // @[RegFile.scala 66:20:@47852.4]
  wire  regs_426_io_enable; // @[RegFile.scala 66:20:@47852.4]
  wire  regs_427_clock; // @[RegFile.scala 66:20:@47866.4]
  wire  regs_427_reset; // @[RegFile.scala 66:20:@47866.4]
  wire [63:0] regs_427_io_in; // @[RegFile.scala 66:20:@47866.4]
  wire  regs_427_io_reset; // @[RegFile.scala 66:20:@47866.4]
  wire [63:0] regs_427_io_out; // @[RegFile.scala 66:20:@47866.4]
  wire  regs_427_io_enable; // @[RegFile.scala 66:20:@47866.4]
  wire  regs_428_clock; // @[RegFile.scala 66:20:@47880.4]
  wire  regs_428_reset; // @[RegFile.scala 66:20:@47880.4]
  wire [63:0] regs_428_io_in; // @[RegFile.scala 66:20:@47880.4]
  wire  regs_428_io_reset; // @[RegFile.scala 66:20:@47880.4]
  wire [63:0] regs_428_io_out; // @[RegFile.scala 66:20:@47880.4]
  wire  regs_428_io_enable; // @[RegFile.scala 66:20:@47880.4]
  wire  regs_429_clock; // @[RegFile.scala 66:20:@47894.4]
  wire  regs_429_reset; // @[RegFile.scala 66:20:@47894.4]
  wire [63:0] regs_429_io_in; // @[RegFile.scala 66:20:@47894.4]
  wire  regs_429_io_reset; // @[RegFile.scala 66:20:@47894.4]
  wire [63:0] regs_429_io_out; // @[RegFile.scala 66:20:@47894.4]
  wire  regs_429_io_enable; // @[RegFile.scala 66:20:@47894.4]
  wire  regs_430_clock; // @[RegFile.scala 66:20:@47908.4]
  wire  regs_430_reset; // @[RegFile.scala 66:20:@47908.4]
  wire [63:0] regs_430_io_in; // @[RegFile.scala 66:20:@47908.4]
  wire  regs_430_io_reset; // @[RegFile.scala 66:20:@47908.4]
  wire [63:0] regs_430_io_out; // @[RegFile.scala 66:20:@47908.4]
  wire  regs_430_io_enable; // @[RegFile.scala 66:20:@47908.4]
  wire  regs_431_clock; // @[RegFile.scala 66:20:@47922.4]
  wire  regs_431_reset; // @[RegFile.scala 66:20:@47922.4]
  wire [63:0] regs_431_io_in; // @[RegFile.scala 66:20:@47922.4]
  wire  regs_431_io_reset; // @[RegFile.scala 66:20:@47922.4]
  wire [63:0] regs_431_io_out; // @[RegFile.scala 66:20:@47922.4]
  wire  regs_431_io_enable; // @[RegFile.scala 66:20:@47922.4]
  wire  regs_432_clock; // @[RegFile.scala 66:20:@47936.4]
  wire  regs_432_reset; // @[RegFile.scala 66:20:@47936.4]
  wire [63:0] regs_432_io_in; // @[RegFile.scala 66:20:@47936.4]
  wire  regs_432_io_reset; // @[RegFile.scala 66:20:@47936.4]
  wire [63:0] regs_432_io_out; // @[RegFile.scala 66:20:@47936.4]
  wire  regs_432_io_enable; // @[RegFile.scala 66:20:@47936.4]
  wire  regs_433_clock; // @[RegFile.scala 66:20:@47950.4]
  wire  regs_433_reset; // @[RegFile.scala 66:20:@47950.4]
  wire [63:0] regs_433_io_in; // @[RegFile.scala 66:20:@47950.4]
  wire  regs_433_io_reset; // @[RegFile.scala 66:20:@47950.4]
  wire [63:0] regs_433_io_out; // @[RegFile.scala 66:20:@47950.4]
  wire  regs_433_io_enable; // @[RegFile.scala 66:20:@47950.4]
  wire  regs_434_clock; // @[RegFile.scala 66:20:@47964.4]
  wire  regs_434_reset; // @[RegFile.scala 66:20:@47964.4]
  wire [63:0] regs_434_io_in; // @[RegFile.scala 66:20:@47964.4]
  wire  regs_434_io_reset; // @[RegFile.scala 66:20:@47964.4]
  wire [63:0] regs_434_io_out; // @[RegFile.scala 66:20:@47964.4]
  wire  regs_434_io_enable; // @[RegFile.scala 66:20:@47964.4]
  wire  regs_435_clock; // @[RegFile.scala 66:20:@47978.4]
  wire  regs_435_reset; // @[RegFile.scala 66:20:@47978.4]
  wire [63:0] regs_435_io_in; // @[RegFile.scala 66:20:@47978.4]
  wire  regs_435_io_reset; // @[RegFile.scala 66:20:@47978.4]
  wire [63:0] regs_435_io_out; // @[RegFile.scala 66:20:@47978.4]
  wire  regs_435_io_enable; // @[RegFile.scala 66:20:@47978.4]
  wire  regs_436_clock; // @[RegFile.scala 66:20:@47992.4]
  wire  regs_436_reset; // @[RegFile.scala 66:20:@47992.4]
  wire [63:0] regs_436_io_in; // @[RegFile.scala 66:20:@47992.4]
  wire  regs_436_io_reset; // @[RegFile.scala 66:20:@47992.4]
  wire [63:0] regs_436_io_out; // @[RegFile.scala 66:20:@47992.4]
  wire  regs_436_io_enable; // @[RegFile.scala 66:20:@47992.4]
  wire  regs_437_clock; // @[RegFile.scala 66:20:@48006.4]
  wire  regs_437_reset; // @[RegFile.scala 66:20:@48006.4]
  wire [63:0] regs_437_io_in; // @[RegFile.scala 66:20:@48006.4]
  wire  regs_437_io_reset; // @[RegFile.scala 66:20:@48006.4]
  wire [63:0] regs_437_io_out; // @[RegFile.scala 66:20:@48006.4]
  wire  regs_437_io_enable; // @[RegFile.scala 66:20:@48006.4]
  wire  regs_438_clock; // @[RegFile.scala 66:20:@48020.4]
  wire  regs_438_reset; // @[RegFile.scala 66:20:@48020.4]
  wire [63:0] regs_438_io_in; // @[RegFile.scala 66:20:@48020.4]
  wire  regs_438_io_reset; // @[RegFile.scala 66:20:@48020.4]
  wire [63:0] regs_438_io_out; // @[RegFile.scala 66:20:@48020.4]
  wire  regs_438_io_enable; // @[RegFile.scala 66:20:@48020.4]
  wire  regs_439_clock; // @[RegFile.scala 66:20:@48034.4]
  wire  regs_439_reset; // @[RegFile.scala 66:20:@48034.4]
  wire [63:0] regs_439_io_in; // @[RegFile.scala 66:20:@48034.4]
  wire  regs_439_io_reset; // @[RegFile.scala 66:20:@48034.4]
  wire [63:0] regs_439_io_out; // @[RegFile.scala 66:20:@48034.4]
  wire  regs_439_io_enable; // @[RegFile.scala 66:20:@48034.4]
  wire  regs_440_clock; // @[RegFile.scala 66:20:@48048.4]
  wire  regs_440_reset; // @[RegFile.scala 66:20:@48048.4]
  wire [63:0] regs_440_io_in; // @[RegFile.scala 66:20:@48048.4]
  wire  regs_440_io_reset; // @[RegFile.scala 66:20:@48048.4]
  wire [63:0] regs_440_io_out; // @[RegFile.scala 66:20:@48048.4]
  wire  regs_440_io_enable; // @[RegFile.scala 66:20:@48048.4]
  wire  regs_441_clock; // @[RegFile.scala 66:20:@48062.4]
  wire  regs_441_reset; // @[RegFile.scala 66:20:@48062.4]
  wire [63:0] regs_441_io_in; // @[RegFile.scala 66:20:@48062.4]
  wire  regs_441_io_reset; // @[RegFile.scala 66:20:@48062.4]
  wire [63:0] regs_441_io_out; // @[RegFile.scala 66:20:@48062.4]
  wire  regs_441_io_enable; // @[RegFile.scala 66:20:@48062.4]
  wire  regs_442_clock; // @[RegFile.scala 66:20:@48076.4]
  wire  regs_442_reset; // @[RegFile.scala 66:20:@48076.4]
  wire [63:0] regs_442_io_in; // @[RegFile.scala 66:20:@48076.4]
  wire  regs_442_io_reset; // @[RegFile.scala 66:20:@48076.4]
  wire [63:0] regs_442_io_out; // @[RegFile.scala 66:20:@48076.4]
  wire  regs_442_io_enable; // @[RegFile.scala 66:20:@48076.4]
  wire  regs_443_clock; // @[RegFile.scala 66:20:@48090.4]
  wire  regs_443_reset; // @[RegFile.scala 66:20:@48090.4]
  wire [63:0] regs_443_io_in; // @[RegFile.scala 66:20:@48090.4]
  wire  regs_443_io_reset; // @[RegFile.scala 66:20:@48090.4]
  wire [63:0] regs_443_io_out; // @[RegFile.scala 66:20:@48090.4]
  wire  regs_443_io_enable; // @[RegFile.scala 66:20:@48090.4]
  wire  regs_444_clock; // @[RegFile.scala 66:20:@48104.4]
  wire  regs_444_reset; // @[RegFile.scala 66:20:@48104.4]
  wire [63:0] regs_444_io_in; // @[RegFile.scala 66:20:@48104.4]
  wire  regs_444_io_reset; // @[RegFile.scala 66:20:@48104.4]
  wire [63:0] regs_444_io_out; // @[RegFile.scala 66:20:@48104.4]
  wire  regs_444_io_enable; // @[RegFile.scala 66:20:@48104.4]
  wire  regs_445_clock; // @[RegFile.scala 66:20:@48118.4]
  wire  regs_445_reset; // @[RegFile.scala 66:20:@48118.4]
  wire [63:0] regs_445_io_in; // @[RegFile.scala 66:20:@48118.4]
  wire  regs_445_io_reset; // @[RegFile.scala 66:20:@48118.4]
  wire [63:0] regs_445_io_out; // @[RegFile.scala 66:20:@48118.4]
  wire  regs_445_io_enable; // @[RegFile.scala 66:20:@48118.4]
  wire  regs_446_clock; // @[RegFile.scala 66:20:@48132.4]
  wire  regs_446_reset; // @[RegFile.scala 66:20:@48132.4]
  wire [63:0] regs_446_io_in; // @[RegFile.scala 66:20:@48132.4]
  wire  regs_446_io_reset; // @[RegFile.scala 66:20:@48132.4]
  wire [63:0] regs_446_io_out; // @[RegFile.scala 66:20:@48132.4]
  wire  regs_446_io_enable; // @[RegFile.scala 66:20:@48132.4]
  wire  regs_447_clock; // @[RegFile.scala 66:20:@48146.4]
  wire  regs_447_reset; // @[RegFile.scala 66:20:@48146.4]
  wire [63:0] regs_447_io_in; // @[RegFile.scala 66:20:@48146.4]
  wire  regs_447_io_reset; // @[RegFile.scala 66:20:@48146.4]
  wire [63:0] regs_447_io_out; // @[RegFile.scala 66:20:@48146.4]
  wire  regs_447_io_enable; // @[RegFile.scala 66:20:@48146.4]
  wire  regs_448_clock; // @[RegFile.scala 66:20:@48160.4]
  wire  regs_448_reset; // @[RegFile.scala 66:20:@48160.4]
  wire [63:0] regs_448_io_in; // @[RegFile.scala 66:20:@48160.4]
  wire  regs_448_io_reset; // @[RegFile.scala 66:20:@48160.4]
  wire [63:0] regs_448_io_out; // @[RegFile.scala 66:20:@48160.4]
  wire  regs_448_io_enable; // @[RegFile.scala 66:20:@48160.4]
  wire  regs_449_clock; // @[RegFile.scala 66:20:@48174.4]
  wire  regs_449_reset; // @[RegFile.scala 66:20:@48174.4]
  wire [63:0] regs_449_io_in; // @[RegFile.scala 66:20:@48174.4]
  wire  regs_449_io_reset; // @[RegFile.scala 66:20:@48174.4]
  wire [63:0] regs_449_io_out; // @[RegFile.scala 66:20:@48174.4]
  wire  regs_449_io_enable; // @[RegFile.scala 66:20:@48174.4]
  wire  regs_450_clock; // @[RegFile.scala 66:20:@48188.4]
  wire  regs_450_reset; // @[RegFile.scala 66:20:@48188.4]
  wire [63:0] regs_450_io_in; // @[RegFile.scala 66:20:@48188.4]
  wire  regs_450_io_reset; // @[RegFile.scala 66:20:@48188.4]
  wire [63:0] regs_450_io_out; // @[RegFile.scala 66:20:@48188.4]
  wire  regs_450_io_enable; // @[RegFile.scala 66:20:@48188.4]
  wire  regs_451_clock; // @[RegFile.scala 66:20:@48202.4]
  wire  regs_451_reset; // @[RegFile.scala 66:20:@48202.4]
  wire [63:0] regs_451_io_in; // @[RegFile.scala 66:20:@48202.4]
  wire  regs_451_io_reset; // @[RegFile.scala 66:20:@48202.4]
  wire [63:0] regs_451_io_out; // @[RegFile.scala 66:20:@48202.4]
  wire  regs_451_io_enable; // @[RegFile.scala 66:20:@48202.4]
  wire  regs_452_clock; // @[RegFile.scala 66:20:@48216.4]
  wire  regs_452_reset; // @[RegFile.scala 66:20:@48216.4]
  wire [63:0] regs_452_io_in; // @[RegFile.scala 66:20:@48216.4]
  wire  regs_452_io_reset; // @[RegFile.scala 66:20:@48216.4]
  wire [63:0] regs_452_io_out; // @[RegFile.scala 66:20:@48216.4]
  wire  regs_452_io_enable; // @[RegFile.scala 66:20:@48216.4]
  wire  regs_453_clock; // @[RegFile.scala 66:20:@48230.4]
  wire  regs_453_reset; // @[RegFile.scala 66:20:@48230.4]
  wire [63:0] regs_453_io_in; // @[RegFile.scala 66:20:@48230.4]
  wire  regs_453_io_reset; // @[RegFile.scala 66:20:@48230.4]
  wire [63:0] regs_453_io_out; // @[RegFile.scala 66:20:@48230.4]
  wire  regs_453_io_enable; // @[RegFile.scala 66:20:@48230.4]
  wire  regs_454_clock; // @[RegFile.scala 66:20:@48244.4]
  wire  regs_454_reset; // @[RegFile.scala 66:20:@48244.4]
  wire [63:0] regs_454_io_in; // @[RegFile.scala 66:20:@48244.4]
  wire  regs_454_io_reset; // @[RegFile.scala 66:20:@48244.4]
  wire [63:0] regs_454_io_out; // @[RegFile.scala 66:20:@48244.4]
  wire  regs_454_io_enable; // @[RegFile.scala 66:20:@48244.4]
  wire  regs_455_clock; // @[RegFile.scala 66:20:@48258.4]
  wire  regs_455_reset; // @[RegFile.scala 66:20:@48258.4]
  wire [63:0] regs_455_io_in; // @[RegFile.scala 66:20:@48258.4]
  wire  regs_455_io_reset; // @[RegFile.scala 66:20:@48258.4]
  wire [63:0] regs_455_io_out; // @[RegFile.scala 66:20:@48258.4]
  wire  regs_455_io_enable; // @[RegFile.scala 66:20:@48258.4]
  wire  regs_456_clock; // @[RegFile.scala 66:20:@48272.4]
  wire  regs_456_reset; // @[RegFile.scala 66:20:@48272.4]
  wire [63:0] regs_456_io_in; // @[RegFile.scala 66:20:@48272.4]
  wire  regs_456_io_reset; // @[RegFile.scala 66:20:@48272.4]
  wire [63:0] regs_456_io_out; // @[RegFile.scala 66:20:@48272.4]
  wire  regs_456_io_enable; // @[RegFile.scala 66:20:@48272.4]
  wire  regs_457_clock; // @[RegFile.scala 66:20:@48286.4]
  wire  regs_457_reset; // @[RegFile.scala 66:20:@48286.4]
  wire [63:0] regs_457_io_in; // @[RegFile.scala 66:20:@48286.4]
  wire  regs_457_io_reset; // @[RegFile.scala 66:20:@48286.4]
  wire [63:0] regs_457_io_out; // @[RegFile.scala 66:20:@48286.4]
  wire  regs_457_io_enable; // @[RegFile.scala 66:20:@48286.4]
  wire  regs_458_clock; // @[RegFile.scala 66:20:@48300.4]
  wire  regs_458_reset; // @[RegFile.scala 66:20:@48300.4]
  wire [63:0] regs_458_io_in; // @[RegFile.scala 66:20:@48300.4]
  wire  regs_458_io_reset; // @[RegFile.scala 66:20:@48300.4]
  wire [63:0] regs_458_io_out; // @[RegFile.scala 66:20:@48300.4]
  wire  regs_458_io_enable; // @[RegFile.scala 66:20:@48300.4]
  wire  regs_459_clock; // @[RegFile.scala 66:20:@48314.4]
  wire  regs_459_reset; // @[RegFile.scala 66:20:@48314.4]
  wire [63:0] regs_459_io_in; // @[RegFile.scala 66:20:@48314.4]
  wire  regs_459_io_reset; // @[RegFile.scala 66:20:@48314.4]
  wire [63:0] regs_459_io_out; // @[RegFile.scala 66:20:@48314.4]
  wire  regs_459_io_enable; // @[RegFile.scala 66:20:@48314.4]
  wire  regs_460_clock; // @[RegFile.scala 66:20:@48328.4]
  wire  regs_460_reset; // @[RegFile.scala 66:20:@48328.4]
  wire [63:0] regs_460_io_in; // @[RegFile.scala 66:20:@48328.4]
  wire  regs_460_io_reset; // @[RegFile.scala 66:20:@48328.4]
  wire [63:0] regs_460_io_out; // @[RegFile.scala 66:20:@48328.4]
  wire  regs_460_io_enable; // @[RegFile.scala 66:20:@48328.4]
  wire  regs_461_clock; // @[RegFile.scala 66:20:@48342.4]
  wire  regs_461_reset; // @[RegFile.scala 66:20:@48342.4]
  wire [63:0] regs_461_io_in; // @[RegFile.scala 66:20:@48342.4]
  wire  regs_461_io_reset; // @[RegFile.scala 66:20:@48342.4]
  wire [63:0] regs_461_io_out; // @[RegFile.scala 66:20:@48342.4]
  wire  regs_461_io_enable; // @[RegFile.scala 66:20:@48342.4]
  wire  regs_462_clock; // @[RegFile.scala 66:20:@48356.4]
  wire  regs_462_reset; // @[RegFile.scala 66:20:@48356.4]
  wire [63:0] regs_462_io_in; // @[RegFile.scala 66:20:@48356.4]
  wire  regs_462_io_reset; // @[RegFile.scala 66:20:@48356.4]
  wire [63:0] regs_462_io_out; // @[RegFile.scala 66:20:@48356.4]
  wire  regs_462_io_enable; // @[RegFile.scala 66:20:@48356.4]
  wire  regs_463_clock; // @[RegFile.scala 66:20:@48370.4]
  wire  regs_463_reset; // @[RegFile.scala 66:20:@48370.4]
  wire [63:0] regs_463_io_in; // @[RegFile.scala 66:20:@48370.4]
  wire  regs_463_io_reset; // @[RegFile.scala 66:20:@48370.4]
  wire [63:0] regs_463_io_out; // @[RegFile.scala 66:20:@48370.4]
  wire  regs_463_io_enable; // @[RegFile.scala 66:20:@48370.4]
  wire  regs_464_clock; // @[RegFile.scala 66:20:@48384.4]
  wire  regs_464_reset; // @[RegFile.scala 66:20:@48384.4]
  wire [63:0] regs_464_io_in; // @[RegFile.scala 66:20:@48384.4]
  wire  regs_464_io_reset; // @[RegFile.scala 66:20:@48384.4]
  wire [63:0] regs_464_io_out; // @[RegFile.scala 66:20:@48384.4]
  wire  regs_464_io_enable; // @[RegFile.scala 66:20:@48384.4]
  wire  regs_465_clock; // @[RegFile.scala 66:20:@48398.4]
  wire  regs_465_reset; // @[RegFile.scala 66:20:@48398.4]
  wire [63:0] regs_465_io_in; // @[RegFile.scala 66:20:@48398.4]
  wire  regs_465_io_reset; // @[RegFile.scala 66:20:@48398.4]
  wire [63:0] regs_465_io_out; // @[RegFile.scala 66:20:@48398.4]
  wire  regs_465_io_enable; // @[RegFile.scala 66:20:@48398.4]
  wire  regs_466_clock; // @[RegFile.scala 66:20:@48412.4]
  wire  regs_466_reset; // @[RegFile.scala 66:20:@48412.4]
  wire [63:0] regs_466_io_in; // @[RegFile.scala 66:20:@48412.4]
  wire  regs_466_io_reset; // @[RegFile.scala 66:20:@48412.4]
  wire [63:0] regs_466_io_out; // @[RegFile.scala 66:20:@48412.4]
  wire  regs_466_io_enable; // @[RegFile.scala 66:20:@48412.4]
  wire  regs_467_clock; // @[RegFile.scala 66:20:@48426.4]
  wire  regs_467_reset; // @[RegFile.scala 66:20:@48426.4]
  wire [63:0] regs_467_io_in; // @[RegFile.scala 66:20:@48426.4]
  wire  regs_467_io_reset; // @[RegFile.scala 66:20:@48426.4]
  wire [63:0] regs_467_io_out; // @[RegFile.scala 66:20:@48426.4]
  wire  regs_467_io_enable; // @[RegFile.scala 66:20:@48426.4]
  wire  regs_468_clock; // @[RegFile.scala 66:20:@48440.4]
  wire  regs_468_reset; // @[RegFile.scala 66:20:@48440.4]
  wire [63:0] regs_468_io_in; // @[RegFile.scala 66:20:@48440.4]
  wire  regs_468_io_reset; // @[RegFile.scala 66:20:@48440.4]
  wire [63:0] regs_468_io_out; // @[RegFile.scala 66:20:@48440.4]
  wire  regs_468_io_enable; // @[RegFile.scala 66:20:@48440.4]
  wire  regs_469_clock; // @[RegFile.scala 66:20:@48454.4]
  wire  regs_469_reset; // @[RegFile.scala 66:20:@48454.4]
  wire [63:0] regs_469_io_in; // @[RegFile.scala 66:20:@48454.4]
  wire  regs_469_io_reset; // @[RegFile.scala 66:20:@48454.4]
  wire [63:0] regs_469_io_out; // @[RegFile.scala 66:20:@48454.4]
  wire  regs_469_io_enable; // @[RegFile.scala 66:20:@48454.4]
  wire  regs_470_clock; // @[RegFile.scala 66:20:@48468.4]
  wire  regs_470_reset; // @[RegFile.scala 66:20:@48468.4]
  wire [63:0] regs_470_io_in; // @[RegFile.scala 66:20:@48468.4]
  wire  regs_470_io_reset; // @[RegFile.scala 66:20:@48468.4]
  wire [63:0] regs_470_io_out; // @[RegFile.scala 66:20:@48468.4]
  wire  regs_470_io_enable; // @[RegFile.scala 66:20:@48468.4]
  wire  regs_471_clock; // @[RegFile.scala 66:20:@48482.4]
  wire  regs_471_reset; // @[RegFile.scala 66:20:@48482.4]
  wire [63:0] regs_471_io_in; // @[RegFile.scala 66:20:@48482.4]
  wire  regs_471_io_reset; // @[RegFile.scala 66:20:@48482.4]
  wire [63:0] regs_471_io_out; // @[RegFile.scala 66:20:@48482.4]
  wire  regs_471_io_enable; // @[RegFile.scala 66:20:@48482.4]
  wire  regs_472_clock; // @[RegFile.scala 66:20:@48496.4]
  wire  regs_472_reset; // @[RegFile.scala 66:20:@48496.4]
  wire [63:0] regs_472_io_in; // @[RegFile.scala 66:20:@48496.4]
  wire  regs_472_io_reset; // @[RegFile.scala 66:20:@48496.4]
  wire [63:0] regs_472_io_out; // @[RegFile.scala 66:20:@48496.4]
  wire  regs_472_io_enable; // @[RegFile.scala 66:20:@48496.4]
  wire  regs_473_clock; // @[RegFile.scala 66:20:@48510.4]
  wire  regs_473_reset; // @[RegFile.scala 66:20:@48510.4]
  wire [63:0] regs_473_io_in; // @[RegFile.scala 66:20:@48510.4]
  wire  regs_473_io_reset; // @[RegFile.scala 66:20:@48510.4]
  wire [63:0] regs_473_io_out; // @[RegFile.scala 66:20:@48510.4]
  wire  regs_473_io_enable; // @[RegFile.scala 66:20:@48510.4]
  wire  regs_474_clock; // @[RegFile.scala 66:20:@48524.4]
  wire  regs_474_reset; // @[RegFile.scala 66:20:@48524.4]
  wire [63:0] regs_474_io_in; // @[RegFile.scala 66:20:@48524.4]
  wire  regs_474_io_reset; // @[RegFile.scala 66:20:@48524.4]
  wire [63:0] regs_474_io_out; // @[RegFile.scala 66:20:@48524.4]
  wire  regs_474_io_enable; // @[RegFile.scala 66:20:@48524.4]
  wire  regs_475_clock; // @[RegFile.scala 66:20:@48538.4]
  wire  regs_475_reset; // @[RegFile.scala 66:20:@48538.4]
  wire [63:0] regs_475_io_in; // @[RegFile.scala 66:20:@48538.4]
  wire  regs_475_io_reset; // @[RegFile.scala 66:20:@48538.4]
  wire [63:0] regs_475_io_out; // @[RegFile.scala 66:20:@48538.4]
  wire  regs_475_io_enable; // @[RegFile.scala 66:20:@48538.4]
  wire  regs_476_clock; // @[RegFile.scala 66:20:@48552.4]
  wire  regs_476_reset; // @[RegFile.scala 66:20:@48552.4]
  wire [63:0] regs_476_io_in; // @[RegFile.scala 66:20:@48552.4]
  wire  regs_476_io_reset; // @[RegFile.scala 66:20:@48552.4]
  wire [63:0] regs_476_io_out; // @[RegFile.scala 66:20:@48552.4]
  wire  regs_476_io_enable; // @[RegFile.scala 66:20:@48552.4]
  wire  regs_477_clock; // @[RegFile.scala 66:20:@48566.4]
  wire  regs_477_reset; // @[RegFile.scala 66:20:@48566.4]
  wire [63:0] regs_477_io_in; // @[RegFile.scala 66:20:@48566.4]
  wire  regs_477_io_reset; // @[RegFile.scala 66:20:@48566.4]
  wire [63:0] regs_477_io_out; // @[RegFile.scala 66:20:@48566.4]
  wire  regs_477_io_enable; // @[RegFile.scala 66:20:@48566.4]
  wire  regs_478_clock; // @[RegFile.scala 66:20:@48580.4]
  wire  regs_478_reset; // @[RegFile.scala 66:20:@48580.4]
  wire [63:0] regs_478_io_in; // @[RegFile.scala 66:20:@48580.4]
  wire  regs_478_io_reset; // @[RegFile.scala 66:20:@48580.4]
  wire [63:0] regs_478_io_out; // @[RegFile.scala 66:20:@48580.4]
  wire  regs_478_io_enable; // @[RegFile.scala 66:20:@48580.4]
  wire  regs_479_clock; // @[RegFile.scala 66:20:@48594.4]
  wire  regs_479_reset; // @[RegFile.scala 66:20:@48594.4]
  wire [63:0] regs_479_io_in; // @[RegFile.scala 66:20:@48594.4]
  wire  regs_479_io_reset; // @[RegFile.scala 66:20:@48594.4]
  wire [63:0] regs_479_io_out; // @[RegFile.scala 66:20:@48594.4]
  wire  regs_479_io_enable; // @[RegFile.scala 66:20:@48594.4]
  wire  regs_480_clock; // @[RegFile.scala 66:20:@48608.4]
  wire  regs_480_reset; // @[RegFile.scala 66:20:@48608.4]
  wire [63:0] regs_480_io_in; // @[RegFile.scala 66:20:@48608.4]
  wire  regs_480_io_reset; // @[RegFile.scala 66:20:@48608.4]
  wire [63:0] regs_480_io_out; // @[RegFile.scala 66:20:@48608.4]
  wire  regs_480_io_enable; // @[RegFile.scala 66:20:@48608.4]
  wire  regs_481_clock; // @[RegFile.scala 66:20:@48622.4]
  wire  regs_481_reset; // @[RegFile.scala 66:20:@48622.4]
  wire [63:0] regs_481_io_in; // @[RegFile.scala 66:20:@48622.4]
  wire  regs_481_io_reset; // @[RegFile.scala 66:20:@48622.4]
  wire [63:0] regs_481_io_out; // @[RegFile.scala 66:20:@48622.4]
  wire  regs_481_io_enable; // @[RegFile.scala 66:20:@48622.4]
  wire  regs_482_clock; // @[RegFile.scala 66:20:@48636.4]
  wire  regs_482_reset; // @[RegFile.scala 66:20:@48636.4]
  wire [63:0] regs_482_io_in; // @[RegFile.scala 66:20:@48636.4]
  wire  regs_482_io_reset; // @[RegFile.scala 66:20:@48636.4]
  wire [63:0] regs_482_io_out; // @[RegFile.scala 66:20:@48636.4]
  wire  regs_482_io_enable; // @[RegFile.scala 66:20:@48636.4]
  wire  regs_483_clock; // @[RegFile.scala 66:20:@48650.4]
  wire  regs_483_reset; // @[RegFile.scala 66:20:@48650.4]
  wire [63:0] regs_483_io_in; // @[RegFile.scala 66:20:@48650.4]
  wire  regs_483_io_reset; // @[RegFile.scala 66:20:@48650.4]
  wire [63:0] regs_483_io_out; // @[RegFile.scala 66:20:@48650.4]
  wire  regs_483_io_enable; // @[RegFile.scala 66:20:@48650.4]
  wire  regs_484_clock; // @[RegFile.scala 66:20:@48664.4]
  wire  regs_484_reset; // @[RegFile.scala 66:20:@48664.4]
  wire [63:0] regs_484_io_in; // @[RegFile.scala 66:20:@48664.4]
  wire  regs_484_io_reset; // @[RegFile.scala 66:20:@48664.4]
  wire [63:0] regs_484_io_out; // @[RegFile.scala 66:20:@48664.4]
  wire  regs_484_io_enable; // @[RegFile.scala 66:20:@48664.4]
  wire  regs_485_clock; // @[RegFile.scala 66:20:@48678.4]
  wire  regs_485_reset; // @[RegFile.scala 66:20:@48678.4]
  wire [63:0] regs_485_io_in; // @[RegFile.scala 66:20:@48678.4]
  wire  regs_485_io_reset; // @[RegFile.scala 66:20:@48678.4]
  wire [63:0] regs_485_io_out; // @[RegFile.scala 66:20:@48678.4]
  wire  regs_485_io_enable; // @[RegFile.scala 66:20:@48678.4]
  wire  regs_486_clock; // @[RegFile.scala 66:20:@48692.4]
  wire  regs_486_reset; // @[RegFile.scala 66:20:@48692.4]
  wire [63:0] regs_486_io_in; // @[RegFile.scala 66:20:@48692.4]
  wire  regs_486_io_reset; // @[RegFile.scala 66:20:@48692.4]
  wire [63:0] regs_486_io_out; // @[RegFile.scala 66:20:@48692.4]
  wire  regs_486_io_enable; // @[RegFile.scala 66:20:@48692.4]
  wire  regs_487_clock; // @[RegFile.scala 66:20:@48706.4]
  wire  regs_487_reset; // @[RegFile.scala 66:20:@48706.4]
  wire [63:0] regs_487_io_in; // @[RegFile.scala 66:20:@48706.4]
  wire  regs_487_io_reset; // @[RegFile.scala 66:20:@48706.4]
  wire [63:0] regs_487_io_out; // @[RegFile.scala 66:20:@48706.4]
  wire  regs_487_io_enable; // @[RegFile.scala 66:20:@48706.4]
  wire  regs_488_clock; // @[RegFile.scala 66:20:@48720.4]
  wire  regs_488_reset; // @[RegFile.scala 66:20:@48720.4]
  wire [63:0] regs_488_io_in; // @[RegFile.scala 66:20:@48720.4]
  wire  regs_488_io_reset; // @[RegFile.scala 66:20:@48720.4]
  wire [63:0] regs_488_io_out; // @[RegFile.scala 66:20:@48720.4]
  wire  regs_488_io_enable; // @[RegFile.scala 66:20:@48720.4]
  wire  regs_489_clock; // @[RegFile.scala 66:20:@48734.4]
  wire  regs_489_reset; // @[RegFile.scala 66:20:@48734.4]
  wire [63:0] regs_489_io_in; // @[RegFile.scala 66:20:@48734.4]
  wire  regs_489_io_reset; // @[RegFile.scala 66:20:@48734.4]
  wire [63:0] regs_489_io_out; // @[RegFile.scala 66:20:@48734.4]
  wire  regs_489_io_enable; // @[RegFile.scala 66:20:@48734.4]
  wire  regs_490_clock; // @[RegFile.scala 66:20:@48748.4]
  wire  regs_490_reset; // @[RegFile.scala 66:20:@48748.4]
  wire [63:0] regs_490_io_in; // @[RegFile.scala 66:20:@48748.4]
  wire  regs_490_io_reset; // @[RegFile.scala 66:20:@48748.4]
  wire [63:0] regs_490_io_out; // @[RegFile.scala 66:20:@48748.4]
  wire  regs_490_io_enable; // @[RegFile.scala 66:20:@48748.4]
  wire  regs_491_clock; // @[RegFile.scala 66:20:@48762.4]
  wire  regs_491_reset; // @[RegFile.scala 66:20:@48762.4]
  wire [63:0] regs_491_io_in; // @[RegFile.scala 66:20:@48762.4]
  wire  regs_491_io_reset; // @[RegFile.scala 66:20:@48762.4]
  wire [63:0] regs_491_io_out; // @[RegFile.scala 66:20:@48762.4]
  wire  regs_491_io_enable; // @[RegFile.scala 66:20:@48762.4]
  wire  regs_492_clock; // @[RegFile.scala 66:20:@48776.4]
  wire  regs_492_reset; // @[RegFile.scala 66:20:@48776.4]
  wire [63:0] regs_492_io_in; // @[RegFile.scala 66:20:@48776.4]
  wire  regs_492_io_reset; // @[RegFile.scala 66:20:@48776.4]
  wire [63:0] regs_492_io_out; // @[RegFile.scala 66:20:@48776.4]
  wire  regs_492_io_enable; // @[RegFile.scala 66:20:@48776.4]
  wire  regs_493_clock; // @[RegFile.scala 66:20:@48790.4]
  wire  regs_493_reset; // @[RegFile.scala 66:20:@48790.4]
  wire [63:0] regs_493_io_in; // @[RegFile.scala 66:20:@48790.4]
  wire  regs_493_io_reset; // @[RegFile.scala 66:20:@48790.4]
  wire [63:0] regs_493_io_out; // @[RegFile.scala 66:20:@48790.4]
  wire  regs_493_io_enable; // @[RegFile.scala 66:20:@48790.4]
  wire  regs_494_clock; // @[RegFile.scala 66:20:@48804.4]
  wire  regs_494_reset; // @[RegFile.scala 66:20:@48804.4]
  wire [63:0] regs_494_io_in; // @[RegFile.scala 66:20:@48804.4]
  wire  regs_494_io_reset; // @[RegFile.scala 66:20:@48804.4]
  wire [63:0] regs_494_io_out; // @[RegFile.scala 66:20:@48804.4]
  wire  regs_494_io_enable; // @[RegFile.scala 66:20:@48804.4]
  wire  regs_495_clock; // @[RegFile.scala 66:20:@48818.4]
  wire  regs_495_reset; // @[RegFile.scala 66:20:@48818.4]
  wire [63:0] regs_495_io_in; // @[RegFile.scala 66:20:@48818.4]
  wire  regs_495_io_reset; // @[RegFile.scala 66:20:@48818.4]
  wire [63:0] regs_495_io_out; // @[RegFile.scala 66:20:@48818.4]
  wire  regs_495_io_enable; // @[RegFile.scala 66:20:@48818.4]
  wire  regs_496_clock; // @[RegFile.scala 66:20:@48832.4]
  wire  regs_496_reset; // @[RegFile.scala 66:20:@48832.4]
  wire [63:0] regs_496_io_in; // @[RegFile.scala 66:20:@48832.4]
  wire  regs_496_io_reset; // @[RegFile.scala 66:20:@48832.4]
  wire [63:0] regs_496_io_out; // @[RegFile.scala 66:20:@48832.4]
  wire  regs_496_io_enable; // @[RegFile.scala 66:20:@48832.4]
  wire  regs_497_clock; // @[RegFile.scala 66:20:@48846.4]
  wire  regs_497_reset; // @[RegFile.scala 66:20:@48846.4]
  wire [63:0] regs_497_io_in; // @[RegFile.scala 66:20:@48846.4]
  wire  regs_497_io_reset; // @[RegFile.scala 66:20:@48846.4]
  wire [63:0] regs_497_io_out; // @[RegFile.scala 66:20:@48846.4]
  wire  regs_497_io_enable; // @[RegFile.scala 66:20:@48846.4]
  wire  regs_498_clock; // @[RegFile.scala 66:20:@48860.4]
  wire  regs_498_reset; // @[RegFile.scala 66:20:@48860.4]
  wire [63:0] regs_498_io_in; // @[RegFile.scala 66:20:@48860.4]
  wire  regs_498_io_reset; // @[RegFile.scala 66:20:@48860.4]
  wire [63:0] regs_498_io_out; // @[RegFile.scala 66:20:@48860.4]
  wire  regs_498_io_enable; // @[RegFile.scala 66:20:@48860.4]
  wire  regs_499_clock; // @[RegFile.scala 66:20:@48874.4]
  wire  regs_499_reset; // @[RegFile.scala 66:20:@48874.4]
  wire [63:0] regs_499_io_in; // @[RegFile.scala 66:20:@48874.4]
  wire  regs_499_io_reset; // @[RegFile.scala 66:20:@48874.4]
  wire [63:0] regs_499_io_out; // @[RegFile.scala 66:20:@48874.4]
  wire  regs_499_io_enable; // @[RegFile.scala 66:20:@48874.4]
  wire  regs_500_clock; // @[RegFile.scala 66:20:@48888.4]
  wire  regs_500_reset; // @[RegFile.scala 66:20:@48888.4]
  wire [63:0] regs_500_io_in; // @[RegFile.scala 66:20:@48888.4]
  wire  regs_500_io_reset; // @[RegFile.scala 66:20:@48888.4]
  wire [63:0] regs_500_io_out; // @[RegFile.scala 66:20:@48888.4]
  wire  regs_500_io_enable; // @[RegFile.scala 66:20:@48888.4]
  wire  regs_501_clock; // @[RegFile.scala 66:20:@48902.4]
  wire  regs_501_reset; // @[RegFile.scala 66:20:@48902.4]
  wire [63:0] regs_501_io_in; // @[RegFile.scala 66:20:@48902.4]
  wire  regs_501_io_reset; // @[RegFile.scala 66:20:@48902.4]
  wire [63:0] regs_501_io_out; // @[RegFile.scala 66:20:@48902.4]
  wire  regs_501_io_enable; // @[RegFile.scala 66:20:@48902.4]
  wire  regs_502_clock; // @[RegFile.scala 66:20:@48916.4]
  wire  regs_502_reset; // @[RegFile.scala 66:20:@48916.4]
  wire [63:0] regs_502_io_in; // @[RegFile.scala 66:20:@48916.4]
  wire  regs_502_io_reset; // @[RegFile.scala 66:20:@48916.4]
  wire [63:0] regs_502_io_out; // @[RegFile.scala 66:20:@48916.4]
  wire  regs_502_io_enable; // @[RegFile.scala 66:20:@48916.4]
  wire  regs_503_clock; // @[RegFile.scala 66:20:@48930.4]
  wire  regs_503_reset; // @[RegFile.scala 66:20:@48930.4]
  wire [63:0] regs_503_io_in; // @[RegFile.scala 66:20:@48930.4]
  wire  regs_503_io_reset; // @[RegFile.scala 66:20:@48930.4]
  wire [63:0] regs_503_io_out; // @[RegFile.scala 66:20:@48930.4]
  wire  regs_503_io_enable; // @[RegFile.scala 66:20:@48930.4]
  wire  regs_504_clock; // @[RegFile.scala 66:20:@48944.4]
  wire  regs_504_reset; // @[RegFile.scala 66:20:@48944.4]
  wire [63:0] regs_504_io_in; // @[RegFile.scala 66:20:@48944.4]
  wire  regs_504_io_reset; // @[RegFile.scala 66:20:@48944.4]
  wire [63:0] regs_504_io_out; // @[RegFile.scala 66:20:@48944.4]
  wire  regs_504_io_enable; // @[RegFile.scala 66:20:@48944.4]
  wire  regs_505_clock; // @[RegFile.scala 66:20:@48958.4]
  wire  regs_505_reset; // @[RegFile.scala 66:20:@48958.4]
  wire [63:0] regs_505_io_in; // @[RegFile.scala 66:20:@48958.4]
  wire  regs_505_io_reset; // @[RegFile.scala 66:20:@48958.4]
  wire [63:0] regs_505_io_out; // @[RegFile.scala 66:20:@48958.4]
  wire  regs_505_io_enable; // @[RegFile.scala 66:20:@48958.4]
  wire  regs_506_clock; // @[RegFile.scala 66:20:@48972.4]
  wire  regs_506_reset; // @[RegFile.scala 66:20:@48972.4]
  wire [63:0] regs_506_io_in; // @[RegFile.scala 66:20:@48972.4]
  wire  regs_506_io_reset; // @[RegFile.scala 66:20:@48972.4]
  wire [63:0] regs_506_io_out; // @[RegFile.scala 66:20:@48972.4]
  wire  regs_506_io_enable; // @[RegFile.scala 66:20:@48972.4]
  wire  regs_507_clock; // @[RegFile.scala 66:20:@48986.4]
  wire  regs_507_reset; // @[RegFile.scala 66:20:@48986.4]
  wire [63:0] regs_507_io_in; // @[RegFile.scala 66:20:@48986.4]
  wire  regs_507_io_reset; // @[RegFile.scala 66:20:@48986.4]
  wire [63:0] regs_507_io_out; // @[RegFile.scala 66:20:@48986.4]
  wire  regs_507_io_enable; // @[RegFile.scala 66:20:@48986.4]
  wire  regs_508_clock; // @[RegFile.scala 66:20:@49000.4]
  wire  regs_508_reset; // @[RegFile.scala 66:20:@49000.4]
  wire [63:0] regs_508_io_in; // @[RegFile.scala 66:20:@49000.4]
  wire  regs_508_io_reset; // @[RegFile.scala 66:20:@49000.4]
  wire [63:0] regs_508_io_out; // @[RegFile.scala 66:20:@49000.4]
  wire  regs_508_io_enable; // @[RegFile.scala 66:20:@49000.4]
  wire  regs_509_clock; // @[RegFile.scala 66:20:@49014.4]
  wire  regs_509_reset; // @[RegFile.scala 66:20:@49014.4]
  wire [63:0] regs_509_io_in; // @[RegFile.scala 66:20:@49014.4]
  wire  regs_509_io_reset; // @[RegFile.scala 66:20:@49014.4]
  wire [63:0] regs_509_io_out; // @[RegFile.scala 66:20:@49014.4]
  wire  regs_509_io_enable; // @[RegFile.scala 66:20:@49014.4]
  wire  regs_510_clock; // @[RegFile.scala 66:20:@49028.4]
  wire  regs_510_reset; // @[RegFile.scala 66:20:@49028.4]
  wire [63:0] regs_510_io_in; // @[RegFile.scala 66:20:@49028.4]
  wire  regs_510_io_reset; // @[RegFile.scala 66:20:@49028.4]
  wire [63:0] regs_510_io_out; // @[RegFile.scala 66:20:@49028.4]
  wire  regs_510_io_enable; // @[RegFile.scala 66:20:@49028.4]
  wire  regs_511_clock; // @[RegFile.scala 66:20:@49042.4]
  wire  regs_511_reset; // @[RegFile.scala 66:20:@49042.4]
  wire [63:0] regs_511_io_in; // @[RegFile.scala 66:20:@49042.4]
  wire  regs_511_io_reset; // @[RegFile.scala 66:20:@49042.4]
  wire [63:0] regs_511_io_out; // @[RegFile.scala 66:20:@49042.4]
  wire  regs_511_io_enable; // @[RegFile.scala 66:20:@49042.4]
  wire  regs_512_clock; // @[RegFile.scala 66:20:@49056.4]
  wire  regs_512_reset; // @[RegFile.scala 66:20:@49056.4]
  wire [63:0] regs_512_io_in; // @[RegFile.scala 66:20:@49056.4]
  wire  regs_512_io_reset; // @[RegFile.scala 66:20:@49056.4]
  wire [63:0] regs_512_io_out; // @[RegFile.scala 66:20:@49056.4]
  wire  regs_512_io_enable; // @[RegFile.scala 66:20:@49056.4]
  wire  regs_513_clock; // @[RegFile.scala 66:20:@49070.4]
  wire  regs_513_reset; // @[RegFile.scala 66:20:@49070.4]
  wire [63:0] regs_513_io_in; // @[RegFile.scala 66:20:@49070.4]
  wire  regs_513_io_reset; // @[RegFile.scala 66:20:@49070.4]
  wire [63:0] regs_513_io_out; // @[RegFile.scala 66:20:@49070.4]
  wire  regs_513_io_enable; // @[RegFile.scala 66:20:@49070.4]
  wire  regs_514_clock; // @[RegFile.scala 66:20:@49084.4]
  wire  regs_514_reset; // @[RegFile.scala 66:20:@49084.4]
  wire [63:0] regs_514_io_in; // @[RegFile.scala 66:20:@49084.4]
  wire  regs_514_io_reset; // @[RegFile.scala 66:20:@49084.4]
  wire [63:0] regs_514_io_out; // @[RegFile.scala 66:20:@49084.4]
  wire  regs_514_io_enable; // @[RegFile.scala 66:20:@49084.4]
  wire  regs_515_clock; // @[RegFile.scala 66:20:@49098.4]
  wire  regs_515_reset; // @[RegFile.scala 66:20:@49098.4]
  wire [63:0] regs_515_io_in; // @[RegFile.scala 66:20:@49098.4]
  wire  regs_515_io_reset; // @[RegFile.scala 66:20:@49098.4]
  wire [63:0] regs_515_io_out; // @[RegFile.scala 66:20:@49098.4]
  wire  regs_515_io_enable; // @[RegFile.scala 66:20:@49098.4]
  wire  regs_516_clock; // @[RegFile.scala 66:20:@49112.4]
  wire  regs_516_reset; // @[RegFile.scala 66:20:@49112.4]
  wire [63:0] regs_516_io_in; // @[RegFile.scala 66:20:@49112.4]
  wire  regs_516_io_reset; // @[RegFile.scala 66:20:@49112.4]
  wire [63:0] regs_516_io_out; // @[RegFile.scala 66:20:@49112.4]
  wire  regs_516_io_enable; // @[RegFile.scala 66:20:@49112.4]
  wire  regs_517_clock; // @[RegFile.scala 66:20:@49126.4]
  wire  regs_517_reset; // @[RegFile.scala 66:20:@49126.4]
  wire [63:0] regs_517_io_in; // @[RegFile.scala 66:20:@49126.4]
  wire  regs_517_io_reset; // @[RegFile.scala 66:20:@49126.4]
  wire [63:0] regs_517_io_out; // @[RegFile.scala 66:20:@49126.4]
  wire  regs_517_io_enable; // @[RegFile.scala 66:20:@49126.4]
  wire  regs_518_clock; // @[RegFile.scala 66:20:@49140.4]
  wire  regs_518_reset; // @[RegFile.scala 66:20:@49140.4]
  wire [63:0] regs_518_io_in; // @[RegFile.scala 66:20:@49140.4]
  wire  regs_518_io_reset; // @[RegFile.scala 66:20:@49140.4]
  wire [63:0] regs_518_io_out; // @[RegFile.scala 66:20:@49140.4]
  wire  regs_518_io_enable; // @[RegFile.scala 66:20:@49140.4]
  wire  regs_519_clock; // @[RegFile.scala 66:20:@49154.4]
  wire  regs_519_reset; // @[RegFile.scala 66:20:@49154.4]
  wire [63:0] regs_519_io_in; // @[RegFile.scala 66:20:@49154.4]
  wire  regs_519_io_reset; // @[RegFile.scala 66:20:@49154.4]
  wire [63:0] regs_519_io_out; // @[RegFile.scala 66:20:@49154.4]
  wire  regs_519_io_enable; // @[RegFile.scala 66:20:@49154.4]
  wire  regs_520_clock; // @[RegFile.scala 66:20:@49168.4]
  wire  regs_520_reset; // @[RegFile.scala 66:20:@49168.4]
  wire [63:0] regs_520_io_in; // @[RegFile.scala 66:20:@49168.4]
  wire  regs_520_io_reset; // @[RegFile.scala 66:20:@49168.4]
  wire [63:0] regs_520_io_out; // @[RegFile.scala 66:20:@49168.4]
  wire  regs_520_io_enable; // @[RegFile.scala 66:20:@49168.4]
  wire  regs_521_clock; // @[RegFile.scala 66:20:@49182.4]
  wire  regs_521_reset; // @[RegFile.scala 66:20:@49182.4]
  wire [63:0] regs_521_io_in; // @[RegFile.scala 66:20:@49182.4]
  wire  regs_521_io_reset; // @[RegFile.scala 66:20:@49182.4]
  wire [63:0] regs_521_io_out; // @[RegFile.scala 66:20:@49182.4]
  wire  regs_521_io_enable; // @[RegFile.scala 66:20:@49182.4]
  wire [63:0] rport_io_ins_0; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_1; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_2; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_3; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_4; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_5; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_6; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_7; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_8; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_9; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_10; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_11; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_12; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_13; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_14; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_15; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_16; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_17; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_18; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_19; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_20; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_21; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_22; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_23; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_24; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_25; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_26; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_27; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_28; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_29; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_30; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_31; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_32; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_33; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_34; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_35; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_36; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_37; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_38; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_39; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_40; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_41; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_42; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_43; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_44; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_45; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_46; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_47; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_48; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_49; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_50; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_51; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_52; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_53; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_54; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_55; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_56; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_57; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_58; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_59; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_60; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_61; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_62; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_63; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_64; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_65; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_66; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_67; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_68; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_69; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_70; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_71; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_72; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_73; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_74; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_75; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_76; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_77; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_78; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_79; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_80; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_81; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_82; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_83; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_84; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_85; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_86; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_87; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_88; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_89; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_90; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_91; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_92; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_93; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_94; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_95; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_96; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_97; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_98; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_99; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_100; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_101; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_102; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_103; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_104; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_105; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_106; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_107; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_108; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_109; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_110; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_111; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_112; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_113; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_114; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_115; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_116; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_117; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_118; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_119; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_120; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_121; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_122; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_123; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_124; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_125; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_126; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_127; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_128; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_129; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_130; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_131; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_132; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_133; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_134; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_135; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_136; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_137; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_138; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_139; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_140; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_141; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_142; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_143; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_144; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_145; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_146; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_147; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_148; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_149; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_150; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_151; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_152; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_153; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_154; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_155; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_156; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_157; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_158; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_159; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_160; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_161; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_162; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_163; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_164; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_165; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_166; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_167; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_168; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_169; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_170; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_171; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_172; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_173; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_174; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_175; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_176; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_177; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_178; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_179; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_180; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_181; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_182; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_183; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_184; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_185; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_186; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_187; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_188; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_189; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_190; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_191; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_192; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_193; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_194; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_195; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_196; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_197; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_198; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_199; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_200; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_201; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_202; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_203; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_204; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_205; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_206; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_207; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_208; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_209; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_210; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_211; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_212; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_213; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_214; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_215; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_216; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_217; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_218; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_219; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_220; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_221; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_222; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_223; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_224; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_225; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_226; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_227; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_228; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_229; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_230; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_231; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_232; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_233; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_234; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_235; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_236; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_237; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_238; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_239; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_240; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_241; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_242; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_243; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_244; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_245; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_246; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_247; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_248; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_249; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_250; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_251; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_252; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_253; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_254; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_255; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_256; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_257; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_258; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_259; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_260; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_261; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_262; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_263; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_264; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_265; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_266; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_267; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_268; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_269; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_270; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_271; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_272; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_273; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_274; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_275; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_276; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_277; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_278; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_279; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_280; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_281; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_282; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_283; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_284; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_285; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_286; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_287; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_288; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_289; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_290; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_291; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_292; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_293; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_294; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_295; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_296; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_297; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_298; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_299; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_300; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_301; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_302; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_303; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_304; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_305; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_306; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_307; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_308; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_309; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_310; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_311; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_312; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_313; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_314; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_315; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_316; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_317; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_318; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_319; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_320; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_321; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_322; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_323; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_324; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_325; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_326; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_327; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_328; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_329; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_330; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_331; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_332; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_333; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_334; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_335; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_336; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_337; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_338; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_339; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_340; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_341; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_342; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_343; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_344; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_345; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_346; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_347; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_348; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_349; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_350; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_351; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_352; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_353; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_354; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_355; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_356; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_357; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_358; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_359; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_360; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_361; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_362; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_363; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_364; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_365; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_366; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_367; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_368; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_369; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_370; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_371; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_372; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_373; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_374; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_375; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_376; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_377; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_378; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_379; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_380; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_381; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_382; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_383; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_384; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_385; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_386; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_387; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_388; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_389; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_390; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_391; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_392; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_393; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_394; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_395; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_396; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_397; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_398; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_399; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_400; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_401; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_402; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_403; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_404; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_405; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_406; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_407; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_408; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_409; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_410; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_411; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_412; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_413; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_414; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_415; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_416; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_417; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_418; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_419; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_420; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_421; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_422; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_423; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_424; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_425; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_426; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_427; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_428; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_429; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_430; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_431; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_432; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_433; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_434; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_435; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_436; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_437; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_438; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_439; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_440; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_441; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_442; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_443; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_444; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_445; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_446; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_447; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_448; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_449; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_450; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_451; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_452; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_453; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_454; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_455; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_456; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_457; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_458; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_459; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_460; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_461; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_462; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_463; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_464; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_465; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_466; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_467; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_468; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_469; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_470; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_471; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_472; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_473; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_474; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_475; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_476; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_477; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_478; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_479; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_480; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_481; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_482; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_483; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_484; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_485; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_486; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_487; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_488; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_489; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_490; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_491; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_492; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_493; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_494; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_495; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_496; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_497; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_498; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_499; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_500; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_501; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_502; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_503; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_504; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_505; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_506; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_507; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_508; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_509; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_510; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_511; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_512; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_513; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_514; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_515; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_516; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_517; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_518; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_519; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_520; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_ins_521; // @[RegFile.scala 95:21:@49196.4]
  wire [9:0] rport_io_sel; // @[RegFile.scala 95:21:@49196.4]
  wire [63:0] rport_io_out; // @[RegFile.scala 95:21:@49196.4]
  wire  _T_3190; // @[RegFile.scala 80:42:@41890.4]
  wire  _T_3196; // @[RegFile.scala 68:46:@41902.4]
  wire  _T_3197; // @[RegFile.scala 68:34:@41903.4]
  wire  _T_3210; // @[RegFile.scala 80:42:@41921.4]
  wire  _T_3216; // @[RegFile.scala 74:80:@41933.4]
  wire  _T_3217; // @[RegFile.scala 74:68:@41934.4]
  wire  _T_3223; // @[RegFile.scala 74:80:@41947.4]
  wire  _T_3224; // @[RegFile.scala 74:68:@41948.4]
  wire  _T_3230; // @[RegFile.scala 74:80:@41961.4]
  wire  _T_3231; // @[RegFile.scala 74:68:@41962.4]
  wire  _T_3237; // @[RegFile.scala 74:80:@41975.4]
  wire  _T_3238; // @[RegFile.scala 74:68:@41976.4]
  wire  _T_3244; // @[RegFile.scala 74:80:@41989.4]
  wire  _T_3245; // @[RegFile.scala 74:68:@41990.4]
  wire  _T_3251; // @[RegFile.scala 74:80:@42003.4]
  wire  _T_3252; // @[RegFile.scala 74:68:@42004.4]
  wire  _T_3258; // @[RegFile.scala 74:80:@42017.4]
  wire  _T_3259; // @[RegFile.scala 74:68:@42018.4]
  wire  _T_3265; // @[RegFile.scala 74:80:@42031.4]
  wire  _T_3266; // @[RegFile.scala 74:68:@42032.4]
  wire  _T_3272; // @[RegFile.scala 74:80:@42045.4]
  wire  _T_3273; // @[RegFile.scala 74:68:@42046.4]
  wire  _T_3279; // @[RegFile.scala 74:80:@42059.4]
  wire  _T_3280; // @[RegFile.scala 74:68:@42060.4]
  wire  _T_3286; // @[RegFile.scala 74:80:@42073.4]
  wire  _T_3287; // @[RegFile.scala 74:68:@42074.4]
  wire  _T_3293; // @[RegFile.scala 74:80:@42087.4]
  wire  _T_3294; // @[RegFile.scala 74:68:@42088.4]
  wire  _T_3300; // @[RegFile.scala 74:80:@42101.4]
  wire  _T_3301; // @[RegFile.scala 74:68:@42102.4]
  wire  _T_3307; // @[RegFile.scala 74:80:@42115.4]
  wire  _T_3308; // @[RegFile.scala 74:68:@42116.4]
  wire  _T_3314; // @[RegFile.scala 74:80:@42129.4]
  wire  _T_3315; // @[RegFile.scala 74:68:@42130.4]
  wire  _T_3321; // @[RegFile.scala 74:80:@42143.4]
  wire  _T_3322; // @[RegFile.scala 74:68:@42144.4]
  wire  _T_3328; // @[RegFile.scala 74:80:@42157.4]
  wire  _T_3329; // @[RegFile.scala 74:68:@42158.4]
  wire  _T_3335; // @[RegFile.scala 74:80:@42171.4]
  wire  _T_3336; // @[RegFile.scala 74:68:@42172.4]
  wire  _T_3342; // @[RegFile.scala 74:80:@42185.4]
  wire  _T_3343; // @[RegFile.scala 74:68:@42186.4]
  wire  _T_3349; // @[RegFile.scala 74:80:@42199.4]
  wire  _T_3350; // @[RegFile.scala 74:68:@42200.4]
  FringeFF regs_0 ( // @[RegFile.scala 66:20:@41887.4]
    .clock(regs_0_clock),
    .reset(regs_0_reset),
    .io_in(regs_0_io_in),
    .io_reset(regs_0_io_reset),
    .io_out(regs_0_io_out),
    .io_enable(regs_0_io_enable)
  );
  FringeFF regs_1 ( // @[RegFile.scala 66:20:@41899.4]
    .clock(regs_1_clock),
    .reset(regs_1_reset),
    .io_in(regs_1_io_in),
    .io_reset(regs_1_io_reset),
    .io_out(regs_1_io_out),
    .io_enable(regs_1_io_enable)
  );
  FringeFF regs_2 ( // @[RegFile.scala 66:20:@41918.4]
    .clock(regs_2_clock),
    .reset(regs_2_reset),
    .io_in(regs_2_io_in),
    .io_reset(regs_2_io_reset),
    .io_out(regs_2_io_out),
    .io_enable(regs_2_io_enable)
  );
  FringeFF regs_3 ( // @[RegFile.scala 66:20:@41930.4]
    .clock(regs_3_clock),
    .reset(regs_3_reset),
    .io_in(regs_3_io_in),
    .io_reset(regs_3_io_reset),
    .io_out(regs_3_io_out),
    .io_enable(regs_3_io_enable)
  );
  FringeFF regs_4 ( // @[RegFile.scala 66:20:@41944.4]
    .clock(regs_4_clock),
    .reset(regs_4_reset),
    .io_in(regs_4_io_in),
    .io_reset(regs_4_io_reset),
    .io_out(regs_4_io_out),
    .io_enable(regs_4_io_enable)
  );
  FringeFF regs_5 ( // @[RegFile.scala 66:20:@41958.4]
    .clock(regs_5_clock),
    .reset(regs_5_reset),
    .io_in(regs_5_io_in),
    .io_reset(regs_5_io_reset),
    .io_out(regs_5_io_out),
    .io_enable(regs_5_io_enable)
  );
  FringeFF regs_6 ( // @[RegFile.scala 66:20:@41972.4]
    .clock(regs_6_clock),
    .reset(regs_6_reset),
    .io_in(regs_6_io_in),
    .io_reset(regs_6_io_reset),
    .io_out(regs_6_io_out),
    .io_enable(regs_6_io_enable)
  );
  FringeFF regs_7 ( // @[RegFile.scala 66:20:@41986.4]
    .clock(regs_7_clock),
    .reset(regs_7_reset),
    .io_in(regs_7_io_in),
    .io_reset(regs_7_io_reset),
    .io_out(regs_7_io_out),
    .io_enable(regs_7_io_enable)
  );
  FringeFF regs_8 ( // @[RegFile.scala 66:20:@42000.4]
    .clock(regs_8_clock),
    .reset(regs_8_reset),
    .io_in(regs_8_io_in),
    .io_reset(regs_8_io_reset),
    .io_out(regs_8_io_out),
    .io_enable(regs_8_io_enable)
  );
  FringeFF regs_9 ( // @[RegFile.scala 66:20:@42014.4]
    .clock(regs_9_clock),
    .reset(regs_9_reset),
    .io_in(regs_9_io_in),
    .io_reset(regs_9_io_reset),
    .io_out(regs_9_io_out),
    .io_enable(regs_9_io_enable)
  );
  FringeFF regs_10 ( // @[RegFile.scala 66:20:@42028.4]
    .clock(regs_10_clock),
    .reset(regs_10_reset),
    .io_in(regs_10_io_in),
    .io_reset(regs_10_io_reset),
    .io_out(regs_10_io_out),
    .io_enable(regs_10_io_enable)
  );
  FringeFF regs_11 ( // @[RegFile.scala 66:20:@42042.4]
    .clock(regs_11_clock),
    .reset(regs_11_reset),
    .io_in(regs_11_io_in),
    .io_reset(regs_11_io_reset),
    .io_out(regs_11_io_out),
    .io_enable(regs_11_io_enable)
  );
  FringeFF regs_12 ( // @[RegFile.scala 66:20:@42056.4]
    .clock(regs_12_clock),
    .reset(regs_12_reset),
    .io_in(regs_12_io_in),
    .io_reset(regs_12_io_reset),
    .io_out(regs_12_io_out),
    .io_enable(regs_12_io_enable)
  );
  FringeFF regs_13 ( // @[RegFile.scala 66:20:@42070.4]
    .clock(regs_13_clock),
    .reset(regs_13_reset),
    .io_in(regs_13_io_in),
    .io_reset(regs_13_io_reset),
    .io_out(regs_13_io_out),
    .io_enable(regs_13_io_enable)
  );
  FringeFF regs_14 ( // @[RegFile.scala 66:20:@42084.4]
    .clock(regs_14_clock),
    .reset(regs_14_reset),
    .io_in(regs_14_io_in),
    .io_reset(regs_14_io_reset),
    .io_out(regs_14_io_out),
    .io_enable(regs_14_io_enable)
  );
  FringeFF regs_15 ( // @[RegFile.scala 66:20:@42098.4]
    .clock(regs_15_clock),
    .reset(regs_15_reset),
    .io_in(regs_15_io_in),
    .io_reset(regs_15_io_reset),
    .io_out(regs_15_io_out),
    .io_enable(regs_15_io_enable)
  );
  FringeFF regs_16 ( // @[RegFile.scala 66:20:@42112.4]
    .clock(regs_16_clock),
    .reset(regs_16_reset),
    .io_in(regs_16_io_in),
    .io_reset(regs_16_io_reset),
    .io_out(regs_16_io_out),
    .io_enable(regs_16_io_enable)
  );
  FringeFF regs_17 ( // @[RegFile.scala 66:20:@42126.4]
    .clock(regs_17_clock),
    .reset(regs_17_reset),
    .io_in(regs_17_io_in),
    .io_reset(regs_17_io_reset),
    .io_out(regs_17_io_out),
    .io_enable(regs_17_io_enable)
  );
  FringeFF regs_18 ( // @[RegFile.scala 66:20:@42140.4]
    .clock(regs_18_clock),
    .reset(regs_18_reset),
    .io_in(regs_18_io_in),
    .io_reset(regs_18_io_reset),
    .io_out(regs_18_io_out),
    .io_enable(regs_18_io_enable)
  );
  FringeFF regs_19 ( // @[RegFile.scala 66:20:@42154.4]
    .clock(regs_19_clock),
    .reset(regs_19_reset),
    .io_in(regs_19_io_in),
    .io_reset(regs_19_io_reset),
    .io_out(regs_19_io_out),
    .io_enable(regs_19_io_enable)
  );
  FringeFF regs_20 ( // @[RegFile.scala 66:20:@42168.4]
    .clock(regs_20_clock),
    .reset(regs_20_reset),
    .io_in(regs_20_io_in),
    .io_reset(regs_20_io_reset),
    .io_out(regs_20_io_out),
    .io_enable(regs_20_io_enable)
  );
  FringeFF regs_21 ( // @[RegFile.scala 66:20:@42182.4]
    .clock(regs_21_clock),
    .reset(regs_21_reset),
    .io_in(regs_21_io_in),
    .io_reset(regs_21_io_reset),
    .io_out(regs_21_io_out),
    .io_enable(regs_21_io_enable)
  );
  FringeFF regs_22 ( // @[RegFile.scala 66:20:@42196.4]
    .clock(regs_22_clock),
    .reset(regs_22_reset),
    .io_in(regs_22_io_in),
    .io_reset(regs_22_io_reset),
    .io_out(regs_22_io_out),
    .io_enable(regs_22_io_enable)
  );
  FringeFF regs_23 ( // @[RegFile.scala 66:20:@42210.4]
    .clock(regs_23_clock),
    .reset(regs_23_reset),
    .io_in(regs_23_io_in),
    .io_reset(regs_23_io_reset),
    .io_out(regs_23_io_out),
    .io_enable(regs_23_io_enable)
  );
  FringeFF regs_24 ( // @[RegFile.scala 66:20:@42224.4]
    .clock(regs_24_clock),
    .reset(regs_24_reset),
    .io_in(regs_24_io_in),
    .io_reset(regs_24_io_reset),
    .io_out(regs_24_io_out),
    .io_enable(regs_24_io_enable)
  );
  FringeFF regs_25 ( // @[RegFile.scala 66:20:@42238.4]
    .clock(regs_25_clock),
    .reset(regs_25_reset),
    .io_in(regs_25_io_in),
    .io_reset(regs_25_io_reset),
    .io_out(regs_25_io_out),
    .io_enable(regs_25_io_enable)
  );
  FringeFF regs_26 ( // @[RegFile.scala 66:20:@42252.4]
    .clock(regs_26_clock),
    .reset(regs_26_reset),
    .io_in(regs_26_io_in),
    .io_reset(regs_26_io_reset),
    .io_out(regs_26_io_out),
    .io_enable(regs_26_io_enable)
  );
  FringeFF regs_27 ( // @[RegFile.scala 66:20:@42266.4]
    .clock(regs_27_clock),
    .reset(regs_27_reset),
    .io_in(regs_27_io_in),
    .io_reset(regs_27_io_reset),
    .io_out(regs_27_io_out),
    .io_enable(regs_27_io_enable)
  );
  FringeFF regs_28 ( // @[RegFile.scala 66:20:@42280.4]
    .clock(regs_28_clock),
    .reset(regs_28_reset),
    .io_in(regs_28_io_in),
    .io_reset(regs_28_io_reset),
    .io_out(regs_28_io_out),
    .io_enable(regs_28_io_enable)
  );
  FringeFF regs_29 ( // @[RegFile.scala 66:20:@42294.4]
    .clock(regs_29_clock),
    .reset(regs_29_reset),
    .io_in(regs_29_io_in),
    .io_reset(regs_29_io_reset),
    .io_out(regs_29_io_out),
    .io_enable(regs_29_io_enable)
  );
  FringeFF regs_30 ( // @[RegFile.scala 66:20:@42308.4]
    .clock(regs_30_clock),
    .reset(regs_30_reset),
    .io_in(regs_30_io_in),
    .io_reset(regs_30_io_reset),
    .io_out(regs_30_io_out),
    .io_enable(regs_30_io_enable)
  );
  FringeFF regs_31 ( // @[RegFile.scala 66:20:@42322.4]
    .clock(regs_31_clock),
    .reset(regs_31_reset),
    .io_in(regs_31_io_in),
    .io_reset(regs_31_io_reset),
    .io_out(regs_31_io_out),
    .io_enable(regs_31_io_enable)
  );
  FringeFF regs_32 ( // @[RegFile.scala 66:20:@42336.4]
    .clock(regs_32_clock),
    .reset(regs_32_reset),
    .io_in(regs_32_io_in),
    .io_reset(regs_32_io_reset),
    .io_out(regs_32_io_out),
    .io_enable(regs_32_io_enable)
  );
  FringeFF regs_33 ( // @[RegFile.scala 66:20:@42350.4]
    .clock(regs_33_clock),
    .reset(regs_33_reset),
    .io_in(regs_33_io_in),
    .io_reset(regs_33_io_reset),
    .io_out(regs_33_io_out),
    .io_enable(regs_33_io_enable)
  );
  FringeFF regs_34 ( // @[RegFile.scala 66:20:@42364.4]
    .clock(regs_34_clock),
    .reset(regs_34_reset),
    .io_in(regs_34_io_in),
    .io_reset(regs_34_io_reset),
    .io_out(regs_34_io_out),
    .io_enable(regs_34_io_enable)
  );
  FringeFF regs_35 ( // @[RegFile.scala 66:20:@42378.4]
    .clock(regs_35_clock),
    .reset(regs_35_reset),
    .io_in(regs_35_io_in),
    .io_reset(regs_35_io_reset),
    .io_out(regs_35_io_out),
    .io_enable(regs_35_io_enable)
  );
  FringeFF regs_36 ( // @[RegFile.scala 66:20:@42392.4]
    .clock(regs_36_clock),
    .reset(regs_36_reset),
    .io_in(regs_36_io_in),
    .io_reset(regs_36_io_reset),
    .io_out(regs_36_io_out),
    .io_enable(regs_36_io_enable)
  );
  FringeFF regs_37 ( // @[RegFile.scala 66:20:@42406.4]
    .clock(regs_37_clock),
    .reset(regs_37_reset),
    .io_in(regs_37_io_in),
    .io_reset(regs_37_io_reset),
    .io_out(regs_37_io_out),
    .io_enable(regs_37_io_enable)
  );
  FringeFF regs_38 ( // @[RegFile.scala 66:20:@42420.4]
    .clock(regs_38_clock),
    .reset(regs_38_reset),
    .io_in(regs_38_io_in),
    .io_reset(regs_38_io_reset),
    .io_out(regs_38_io_out),
    .io_enable(regs_38_io_enable)
  );
  FringeFF regs_39 ( // @[RegFile.scala 66:20:@42434.4]
    .clock(regs_39_clock),
    .reset(regs_39_reset),
    .io_in(regs_39_io_in),
    .io_reset(regs_39_io_reset),
    .io_out(regs_39_io_out),
    .io_enable(regs_39_io_enable)
  );
  FringeFF regs_40 ( // @[RegFile.scala 66:20:@42448.4]
    .clock(regs_40_clock),
    .reset(regs_40_reset),
    .io_in(regs_40_io_in),
    .io_reset(regs_40_io_reset),
    .io_out(regs_40_io_out),
    .io_enable(regs_40_io_enable)
  );
  FringeFF regs_41 ( // @[RegFile.scala 66:20:@42462.4]
    .clock(regs_41_clock),
    .reset(regs_41_reset),
    .io_in(regs_41_io_in),
    .io_reset(regs_41_io_reset),
    .io_out(regs_41_io_out),
    .io_enable(regs_41_io_enable)
  );
  FringeFF regs_42 ( // @[RegFile.scala 66:20:@42476.4]
    .clock(regs_42_clock),
    .reset(regs_42_reset),
    .io_in(regs_42_io_in),
    .io_reset(regs_42_io_reset),
    .io_out(regs_42_io_out),
    .io_enable(regs_42_io_enable)
  );
  FringeFF regs_43 ( // @[RegFile.scala 66:20:@42490.4]
    .clock(regs_43_clock),
    .reset(regs_43_reset),
    .io_in(regs_43_io_in),
    .io_reset(regs_43_io_reset),
    .io_out(regs_43_io_out),
    .io_enable(regs_43_io_enable)
  );
  FringeFF regs_44 ( // @[RegFile.scala 66:20:@42504.4]
    .clock(regs_44_clock),
    .reset(regs_44_reset),
    .io_in(regs_44_io_in),
    .io_reset(regs_44_io_reset),
    .io_out(regs_44_io_out),
    .io_enable(regs_44_io_enable)
  );
  FringeFF regs_45 ( // @[RegFile.scala 66:20:@42518.4]
    .clock(regs_45_clock),
    .reset(regs_45_reset),
    .io_in(regs_45_io_in),
    .io_reset(regs_45_io_reset),
    .io_out(regs_45_io_out),
    .io_enable(regs_45_io_enable)
  );
  FringeFF regs_46 ( // @[RegFile.scala 66:20:@42532.4]
    .clock(regs_46_clock),
    .reset(regs_46_reset),
    .io_in(regs_46_io_in),
    .io_reset(regs_46_io_reset),
    .io_out(regs_46_io_out),
    .io_enable(regs_46_io_enable)
  );
  FringeFF regs_47 ( // @[RegFile.scala 66:20:@42546.4]
    .clock(regs_47_clock),
    .reset(regs_47_reset),
    .io_in(regs_47_io_in),
    .io_reset(regs_47_io_reset),
    .io_out(regs_47_io_out),
    .io_enable(regs_47_io_enable)
  );
  FringeFF regs_48 ( // @[RegFile.scala 66:20:@42560.4]
    .clock(regs_48_clock),
    .reset(regs_48_reset),
    .io_in(regs_48_io_in),
    .io_reset(regs_48_io_reset),
    .io_out(regs_48_io_out),
    .io_enable(regs_48_io_enable)
  );
  FringeFF regs_49 ( // @[RegFile.scala 66:20:@42574.4]
    .clock(regs_49_clock),
    .reset(regs_49_reset),
    .io_in(regs_49_io_in),
    .io_reset(regs_49_io_reset),
    .io_out(regs_49_io_out),
    .io_enable(regs_49_io_enable)
  );
  FringeFF regs_50 ( // @[RegFile.scala 66:20:@42588.4]
    .clock(regs_50_clock),
    .reset(regs_50_reset),
    .io_in(regs_50_io_in),
    .io_reset(regs_50_io_reset),
    .io_out(regs_50_io_out),
    .io_enable(regs_50_io_enable)
  );
  FringeFF regs_51 ( // @[RegFile.scala 66:20:@42602.4]
    .clock(regs_51_clock),
    .reset(regs_51_reset),
    .io_in(regs_51_io_in),
    .io_reset(regs_51_io_reset),
    .io_out(regs_51_io_out),
    .io_enable(regs_51_io_enable)
  );
  FringeFF regs_52 ( // @[RegFile.scala 66:20:@42616.4]
    .clock(regs_52_clock),
    .reset(regs_52_reset),
    .io_in(regs_52_io_in),
    .io_reset(regs_52_io_reset),
    .io_out(regs_52_io_out),
    .io_enable(regs_52_io_enable)
  );
  FringeFF regs_53 ( // @[RegFile.scala 66:20:@42630.4]
    .clock(regs_53_clock),
    .reset(regs_53_reset),
    .io_in(regs_53_io_in),
    .io_reset(regs_53_io_reset),
    .io_out(regs_53_io_out),
    .io_enable(regs_53_io_enable)
  );
  FringeFF regs_54 ( // @[RegFile.scala 66:20:@42644.4]
    .clock(regs_54_clock),
    .reset(regs_54_reset),
    .io_in(regs_54_io_in),
    .io_reset(regs_54_io_reset),
    .io_out(regs_54_io_out),
    .io_enable(regs_54_io_enable)
  );
  FringeFF regs_55 ( // @[RegFile.scala 66:20:@42658.4]
    .clock(regs_55_clock),
    .reset(regs_55_reset),
    .io_in(regs_55_io_in),
    .io_reset(regs_55_io_reset),
    .io_out(regs_55_io_out),
    .io_enable(regs_55_io_enable)
  );
  FringeFF regs_56 ( // @[RegFile.scala 66:20:@42672.4]
    .clock(regs_56_clock),
    .reset(regs_56_reset),
    .io_in(regs_56_io_in),
    .io_reset(regs_56_io_reset),
    .io_out(regs_56_io_out),
    .io_enable(regs_56_io_enable)
  );
  FringeFF regs_57 ( // @[RegFile.scala 66:20:@42686.4]
    .clock(regs_57_clock),
    .reset(regs_57_reset),
    .io_in(regs_57_io_in),
    .io_reset(regs_57_io_reset),
    .io_out(regs_57_io_out),
    .io_enable(regs_57_io_enable)
  );
  FringeFF regs_58 ( // @[RegFile.scala 66:20:@42700.4]
    .clock(regs_58_clock),
    .reset(regs_58_reset),
    .io_in(regs_58_io_in),
    .io_reset(regs_58_io_reset),
    .io_out(regs_58_io_out),
    .io_enable(regs_58_io_enable)
  );
  FringeFF regs_59 ( // @[RegFile.scala 66:20:@42714.4]
    .clock(regs_59_clock),
    .reset(regs_59_reset),
    .io_in(regs_59_io_in),
    .io_reset(regs_59_io_reset),
    .io_out(regs_59_io_out),
    .io_enable(regs_59_io_enable)
  );
  FringeFF regs_60 ( // @[RegFile.scala 66:20:@42728.4]
    .clock(regs_60_clock),
    .reset(regs_60_reset),
    .io_in(regs_60_io_in),
    .io_reset(regs_60_io_reset),
    .io_out(regs_60_io_out),
    .io_enable(regs_60_io_enable)
  );
  FringeFF regs_61 ( // @[RegFile.scala 66:20:@42742.4]
    .clock(regs_61_clock),
    .reset(regs_61_reset),
    .io_in(regs_61_io_in),
    .io_reset(regs_61_io_reset),
    .io_out(regs_61_io_out),
    .io_enable(regs_61_io_enable)
  );
  FringeFF regs_62 ( // @[RegFile.scala 66:20:@42756.4]
    .clock(regs_62_clock),
    .reset(regs_62_reset),
    .io_in(regs_62_io_in),
    .io_reset(regs_62_io_reset),
    .io_out(regs_62_io_out),
    .io_enable(regs_62_io_enable)
  );
  FringeFF regs_63 ( // @[RegFile.scala 66:20:@42770.4]
    .clock(regs_63_clock),
    .reset(regs_63_reset),
    .io_in(regs_63_io_in),
    .io_reset(regs_63_io_reset),
    .io_out(regs_63_io_out),
    .io_enable(regs_63_io_enable)
  );
  FringeFF regs_64 ( // @[RegFile.scala 66:20:@42784.4]
    .clock(regs_64_clock),
    .reset(regs_64_reset),
    .io_in(regs_64_io_in),
    .io_reset(regs_64_io_reset),
    .io_out(regs_64_io_out),
    .io_enable(regs_64_io_enable)
  );
  FringeFF regs_65 ( // @[RegFile.scala 66:20:@42798.4]
    .clock(regs_65_clock),
    .reset(regs_65_reset),
    .io_in(regs_65_io_in),
    .io_reset(regs_65_io_reset),
    .io_out(regs_65_io_out),
    .io_enable(regs_65_io_enable)
  );
  FringeFF regs_66 ( // @[RegFile.scala 66:20:@42812.4]
    .clock(regs_66_clock),
    .reset(regs_66_reset),
    .io_in(regs_66_io_in),
    .io_reset(regs_66_io_reset),
    .io_out(regs_66_io_out),
    .io_enable(regs_66_io_enable)
  );
  FringeFF regs_67 ( // @[RegFile.scala 66:20:@42826.4]
    .clock(regs_67_clock),
    .reset(regs_67_reset),
    .io_in(regs_67_io_in),
    .io_reset(regs_67_io_reset),
    .io_out(regs_67_io_out),
    .io_enable(regs_67_io_enable)
  );
  FringeFF regs_68 ( // @[RegFile.scala 66:20:@42840.4]
    .clock(regs_68_clock),
    .reset(regs_68_reset),
    .io_in(regs_68_io_in),
    .io_reset(regs_68_io_reset),
    .io_out(regs_68_io_out),
    .io_enable(regs_68_io_enable)
  );
  FringeFF regs_69 ( // @[RegFile.scala 66:20:@42854.4]
    .clock(regs_69_clock),
    .reset(regs_69_reset),
    .io_in(regs_69_io_in),
    .io_reset(regs_69_io_reset),
    .io_out(regs_69_io_out),
    .io_enable(regs_69_io_enable)
  );
  FringeFF regs_70 ( // @[RegFile.scala 66:20:@42868.4]
    .clock(regs_70_clock),
    .reset(regs_70_reset),
    .io_in(regs_70_io_in),
    .io_reset(regs_70_io_reset),
    .io_out(regs_70_io_out),
    .io_enable(regs_70_io_enable)
  );
  FringeFF regs_71 ( // @[RegFile.scala 66:20:@42882.4]
    .clock(regs_71_clock),
    .reset(regs_71_reset),
    .io_in(regs_71_io_in),
    .io_reset(regs_71_io_reset),
    .io_out(regs_71_io_out),
    .io_enable(regs_71_io_enable)
  );
  FringeFF regs_72 ( // @[RegFile.scala 66:20:@42896.4]
    .clock(regs_72_clock),
    .reset(regs_72_reset),
    .io_in(regs_72_io_in),
    .io_reset(regs_72_io_reset),
    .io_out(regs_72_io_out),
    .io_enable(regs_72_io_enable)
  );
  FringeFF regs_73 ( // @[RegFile.scala 66:20:@42910.4]
    .clock(regs_73_clock),
    .reset(regs_73_reset),
    .io_in(regs_73_io_in),
    .io_reset(regs_73_io_reset),
    .io_out(regs_73_io_out),
    .io_enable(regs_73_io_enable)
  );
  FringeFF regs_74 ( // @[RegFile.scala 66:20:@42924.4]
    .clock(regs_74_clock),
    .reset(regs_74_reset),
    .io_in(regs_74_io_in),
    .io_reset(regs_74_io_reset),
    .io_out(regs_74_io_out),
    .io_enable(regs_74_io_enable)
  );
  FringeFF regs_75 ( // @[RegFile.scala 66:20:@42938.4]
    .clock(regs_75_clock),
    .reset(regs_75_reset),
    .io_in(regs_75_io_in),
    .io_reset(regs_75_io_reset),
    .io_out(regs_75_io_out),
    .io_enable(regs_75_io_enable)
  );
  FringeFF regs_76 ( // @[RegFile.scala 66:20:@42952.4]
    .clock(regs_76_clock),
    .reset(regs_76_reset),
    .io_in(regs_76_io_in),
    .io_reset(regs_76_io_reset),
    .io_out(regs_76_io_out),
    .io_enable(regs_76_io_enable)
  );
  FringeFF regs_77 ( // @[RegFile.scala 66:20:@42966.4]
    .clock(regs_77_clock),
    .reset(regs_77_reset),
    .io_in(regs_77_io_in),
    .io_reset(regs_77_io_reset),
    .io_out(regs_77_io_out),
    .io_enable(regs_77_io_enable)
  );
  FringeFF regs_78 ( // @[RegFile.scala 66:20:@42980.4]
    .clock(regs_78_clock),
    .reset(regs_78_reset),
    .io_in(regs_78_io_in),
    .io_reset(regs_78_io_reset),
    .io_out(regs_78_io_out),
    .io_enable(regs_78_io_enable)
  );
  FringeFF regs_79 ( // @[RegFile.scala 66:20:@42994.4]
    .clock(regs_79_clock),
    .reset(regs_79_reset),
    .io_in(regs_79_io_in),
    .io_reset(regs_79_io_reset),
    .io_out(regs_79_io_out),
    .io_enable(regs_79_io_enable)
  );
  FringeFF regs_80 ( // @[RegFile.scala 66:20:@43008.4]
    .clock(regs_80_clock),
    .reset(regs_80_reset),
    .io_in(regs_80_io_in),
    .io_reset(regs_80_io_reset),
    .io_out(regs_80_io_out),
    .io_enable(regs_80_io_enable)
  );
  FringeFF regs_81 ( // @[RegFile.scala 66:20:@43022.4]
    .clock(regs_81_clock),
    .reset(regs_81_reset),
    .io_in(regs_81_io_in),
    .io_reset(regs_81_io_reset),
    .io_out(regs_81_io_out),
    .io_enable(regs_81_io_enable)
  );
  FringeFF regs_82 ( // @[RegFile.scala 66:20:@43036.4]
    .clock(regs_82_clock),
    .reset(regs_82_reset),
    .io_in(regs_82_io_in),
    .io_reset(regs_82_io_reset),
    .io_out(regs_82_io_out),
    .io_enable(regs_82_io_enable)
  );
  FringeFF regs_83 ( // @[RegFile.scala 66:20:@43050.4]
    .clock(regs_83_clock),
    .reset(regs_83_reset),
    .io_in(regs_83_io_in),
    .io_reset(regs_83_io_reset),
    .io_out(regs_83_io_out),
    .io_enable(regs_83_io_enable)
  );
  FringeFF regs_84 ( // @[RegFile.scala 66:20:@43064.4]
    .clock(regs_84_clock),
    .reset(regs_84_reset),
    .io_in(regs_84_io_in),
    .io_reset(regs_84_io_reset),
    .io_out(regs_84_io_out),
    .io_enable(regs_84_io_enable)
  );
  FringeFF regs_85 ( // @[RegFile.scala 66:20:@43078.4]
    .clock(regs_85_clock),
    .reset(regs_85_reset),
    .io_in(regs_85_io_in),
    .io_reset(regs_85_io_reset),
    .io_out(regs_85_io_out),
    .io_enable(regs_85_io_enable)
  );
  FringeFF regs_86 ( // @[RegFile.scala 66:20:@43092.4]
    .clock(regs_86_clock),
    .reset(regs_86_reset),
    .io_in(regs_86_io_in),
    .io_reset(regs_86_io_reset),
    .io_out(regs_86_io_out),
    .io_enable(regs_86_io_enable)
  );
  FringeFF regs_87 ( // @[RegFile.scala 66:20:@43106.4]
    .clock(regs_87_clock),
    .reset(regs_87_reset),
    .io_in(regs_87_io_in),
    .io_reset(regs_87_io_reset),
    .io_out(regs_87_io_out),
    .io_enable(regs_87_io_enable)
  );
  FringeFF regs_88 ( // @[RegFile.scala 66:20:@43120.4]
    .clock(regs_88_clock),
    .reset(regs_88_reset),
    .io_in(regs_88_io_in),
    .io_reset(regs_88_io_reset),
    .io_out(regs_88_io_out),
    .io_enable(regs_88_io_enable)
  );
  FringeFF regs_89 ( // @[RegFile.scala 66:20:@43134.4]
    .clock(regs_89_clock),
    .reset(regs_89_reset),
    .io_in(regs_89_io_in),
    .io_reset(regs_89_io_reset),
    .io_out(regs_89_io_out),
    .io_enable(regs_89_io_enable)
  );
  FringeFF regs_90 ( // @[RegFile.scala 66:20:@43148.4]
    .clock(regs_90_clock),
    .reset(regs_90_reset),
    .io_in(regs_90_io_in),
    .io_reset(regs_90_io_reset),
    .io_out(regs_90_io_out),
    .io_enable(regs_90_io_enable)
  );
  FringeFF regs_91 ( // @[RegFile.scala 66:20:@43162.4]
    .clock(regs_91_clock),
    .reset(regs_91_reset),
    .io_in(regs_91_io_in),
    .io_reset(regs_91_io_reset),
    .io_out(regs_91_io_out),
    .io_enable(regs_91_io_enable)
  );
  FringeFF regs_92 ( // @[RegFile.scala 66:20:@43176.4]
    .clock(regs_92_clock),
    .reset(regs_92_reset),
    .io_in(regs_92_io_in),
    .io_reset(regs_92_io_reset),
    .io_out(regs_92_io_out),
    .io_enable(regs_92_io_enable)
  );
  FringeFF regs_93 ( // @[RegFile.scala 66:20:@43190.4]
    .clock(regs_93_clock),
    .reset(regs_93_reset),
    .io_in(regs_93_io_in),
    .io_reset(regs_93_io_reset),
    .io_out(regs_93_io_out),
    .io_enable(regs_93_io_enable)
  );
  FringeFF regs_94 ( // @[RegFile.scala 66:20:@43204.4]
    .clock(regs_94_clock),
    .reset(regs_94_reset),
    .io_in(regs_94_io_in),
    .io_reset(regs_94_io_reset),
    .io_out(regs_94_io_out),
    .io_enable(regs_94_io_enable)
  );
  FringeFF regs_95 ( // @[RegFile.scala 66:20:@43218.4]
    .clock(regs_95_clock),
    .reset(regs_95_reset),
    .io_in(regs_95_io_in),
    .io_reset(regs_95_io_reset),
    .io_out(regs_95_io_out),
    .io_enable(regs_95_io_enable)
  );
  FringeFF regs_96 ( // @[RegFile.scala 66:20:@43232.4]
    .clock(regs_96_clock),
    .reset(regs_96_reset),
    .io_in(regs_96_io_in),
    .io_reset(regs_96_io_reset),
    .io_out(regs_96_io_out),
    .io_enable(regs_96_io_enable)
  );
  FringeFF regs_97 ( // @[RegFile.scala 66:20:@43246.4]
    .clock(regs_97_clock),
    .reset(regs_97_reset),
    .io_in(regs_97_io_in),
    .io_reset(regs_97_io_reset),
    .io_out(regs_97_io_out),
    .io_enable(regs_97_io_enable)
  );
  FringeFF regs_98 ( // @[RegFile.scala 66:20:@43260.4]
    .clock(regs_98_clock),
    .reset(regs_98_reset),
    .io_in(regs_98_io_in),
    .io_reset(regs_98_io_reset),
    .io_out(regs_98_io_out),
    .io_enable(regs_98_io_enable)
  );
  FringeFF regs_99 ( // @[RegFile.scala 66:20:@43274.4]
    .clock(regs_99_clock),
    .reset(regs_99_reset),
    .io_in(regs_99_io_in),
    .io_reset(regs_99_io_reset),
    .io_out(regs_99_io_out),
    .io_enable(regs_99_io_enable)
  );
  FringeFF regs_100 ( // @[RegFile.scala 66:20:@43288.4]
    .clock(regs_100_clock),
    .reset(regs_100_reset),
    .io_in(regs_100_io_in),
    .io_reset(regs_100_io_reset),
    .io_out(regs_100_io_out),
    .io_enable(regs_100_io_enable)
  );
  FringeFF regs_101 ( // @[RegFile.scala 66:20:@43302.4]
    .clock(regs_101_clock),
    .reset(regs_101_reset),
    .io_in(regs_101_io_in),
    .io_reset(regs_101_io_reset),
    .io_out(regs_101_io_out),
    .io_enable(regs_101_io_enable)
  );
  FringeFF regs_102 ( // @[RegFile.scala 66:20:@43316.4]
    .clock(regs_102_clock),
    .reset(regs_102_reset),
    .io_in(regs_102_io_in),
    .io_reset(regs_102_io_reset),
    .io_out(regs_102_io_out),
    .io_enable(regs_102_io_enable)
  );
  FringeFF regs_103 ( // @[RegFile.scala 66:20:@43330.4]
    .clock(regs_103_clock),
    .reset(regs_103_reset),
    .io_in(regs_103_io_in),
    .io_reset(regs_103_io_reset),
    .io_out(regs_103_io_out),
    .io_enable(regs_103_io_enable)
  );
  FringeFF regs_104 ( // @[RegFile.scala 66:20:@43344.4]
    .clock(regs_104_clock),
    .reset(regs_104_reset),
    .io_in(regs_104_io_in),
    .io_reset(regs_104_io_reset),
    .io_out(regs_104_io_out),
    .io_enable(regs_104_io_enable)
  );
  FringeFF regs_105 ( // @[RegFile.scala 66:20:@43358.4]
    .clock(regs_105_clock),
    .reset(regs_105_reset),
    .io_in(regs_105_io_in),
    .io_reset(regs_105_io_reset),
    .io_out(regs_105_io_out),
    .io_enable(regs_105_io_enable)
  );
  FringeFF regs_106 ( // @[RegFile.scala 66:20:@43372.4]
    .clock(regs_106_clock),
    .reset(regs_106_reset),
    .io_in(regs_106_io_in),
    .io_reset(regs_106_io_reset),
    .io_out(regs_106_io_out),
    .io_enable(regs_106_io_enable)
  );
  FringeFF regs_107 ( // @[RegFile.scala 66:20:@43386.4]
    .clock(regs_107_clock),
    .reset(regs_107_reset),
    .io_in(regs_107_io_in),
    .io_reset(regs_107_io_reset),
    .io_out(regs_107_io_out),
    .io_enable(regs_107_io_enable)
  );
  FringeFF regs_108 ( // @[RegFile.scala 66:20:@43400.4]
    .clock(regs_108_clock),
    .reset(regs_108_reset),
    .io_in(regs_108_io_in),
    .io_reset(regs_108_io_reset),
    .io_out(regs_108_io_out),
    .io_enable(regs_108_io_enable)
  );
  FringeFF regs_109 ( // @[RegFile.scala 66:20:@43414.4]
    .clock(regs_109_clock),
    .reset(regs_109_reset),
    .io_in(regs_109_io_in),
    .io_reset(regs_109_io_reset),
    .io_out(regs_109_io_out),
    .io_enable(regs_109_io_enable)
  );
  FringeFF regs_110 ( // @[RegFile.scala 66:20:@43428.4]
    .clock(regs_110_clock),
    .reset(regs_110_reset),
    .io_in(regs_110_io_in),
    .io_reset(regs_110_io_reset),
    .io_out(regs_110_io_out),
    .io_enable(regs_110_io_enable)
  );
  FringeFF regs_111 ( // @[RegFile.scala 66:20:@43442.4]
    .clock(regs_111_clock),
    .reset(regs_111_reset),
    .io_in(regs_111_io_in),
    .io_reset(regs_111_io_reset),
    .io_out(regs_111_io_out),
    .io_enable(regs_111_io_enable)
  );
  FringeFF regs_112 ( // @[RegFile.scala 66:20:@43456.4]
    .clock(regs_112_clock),
    .reset(regs_112_reset),
    .io_in(regs_112_io_in),
    .io_reset(regs_112_io_reset),
    .io_out(regs_112_io_out),
    .io_enable(regs_112_io_enable)
  );
  FringeFF regs_113 ( // @[RegFile.scala 66:20:@43470.4]
    .clock(regs_113_clock),
    .reset(regs_113_reset),
    .io_in(regs_113_io_in),
    .io_reset(regs_113_io_reset),
    .io_out(regs_113_io_out),
    .io_enable(regs_113_io_enable)
  );
  FringeFF regs_114 ( // @[RegFile.scala 66:20:@43484.4]
    .clock(regs_114_clock),
    .reset(regs_114_reset),
    .io_in(regs_114_io_in),
    .io_reset(regs_114_io_reset),
    .io_out(regs_114_io_out),
    .io_enable(regs_114_io_enable)
  );
  FringeFF regs_115 ( // @[RegFile.scala 66:20:@43498.4]
    .clock(regs_115_clock),
    .reset(regs_115_reset),
    .io_in(regs_115_io_in),
    .io_reset(regs_115_io_reset),
    .io_out(regs_115_io_out),
    .io_enable(regs_115_io_enable)
  );
  FringeFF regs_116 ( // @[RegFile.scala 66:20:@43512.4]
    .clock(regs_116_clock),
    .reset(regs_116_reset),
    .io_in(regs_116_io_in),
    .io_reset(regs_116_io_reset),
    .io_out(regs_116_io_out),
    .io_enable(regs_116_io_enable)
  );
  FringeFF regs_117 ( // @[RegFile.scala 66:20:@43526.4]
    .clock(regs_117_clock),
    .reset(regs_117_reset),
    .io_in(regs_117_io_in),
    .io_reset(regs_117_io_reset),
    .io_out(regs_117_io_out),
    .io_enable(regs_117_io_enable)
  );
  FringeFF regs_118 ( // @[RegFile.scala 66:20:@43540.4]
    .clock(regs_118_clock),
    .reset(regs_118_reset),
    .io_in(regs_118_io_in),
    .io_reset(regs_118_io_reset),
    .io_out(regs_118_io_out),
    .io_enable(regs_118_io_enable)
  );
  FringeFF regs_119 ( // @[RegFile.scala 66:20:@43554.4]
    .clock(regs_119_clock),
    .reset(regs_119_reset),
    .io_in(regs_119_io_in),
    .io_reset(regs_119_io_reset),
    .io_out(regs_119_io_out),
    .io_enable(regs_119_io_enable)
  );
  FringeFF regs_120 ( // @[RegFile.scala 66:20:@43568.4]
    .clock(regs_120_clock),
    .reset(regs_120_reset),
    .io_in(regs_120_io_in),
    .io_reset(regs_120_io_reset),
    .io_out(regs_120_io_out),
    .io_enable(regs_120_io_enable)
  );
  FringeFF regs_121 ( // @[RegFile.scala 66:20:@43582.4]
    .clock(regs_121_clock),
    .reset(regs_121_reset),
    .io_in(regs_121_io_in),
    .io_reset(regs_121_io_reset),
    .io_out(regs_121_io_out),
    .io_enable(regs_121_io_enable)
  );
  FringeFF regs_122 ( // @[RegFile.scala 66:20:@43596.4]
    .clock(regs_122_clock),
    .reset(regs_122_reset),
    .io_in(regs_122_io_in),
    .io_reset(regs_122_io_reset),
    .io_out(regs_122_io_out),
    .io_enable(regs_122_io_enable)
  );
  FringeFF regs_123 ( // @[RegFile.scala 66:20:@43610.4]
    .clock(regs_123_clock),
    .reset(regs_123_reset),
    .io_in(regs_123_io_in),
    .io_reset(regs_123_io_reset),
    .io_out(regs_123_io_out),
    .io_enable(regs_123_io_enable)
  );
  FringeFF regs_124 ( // @[RegFile.scala 66:20:@43624.4]
    .clock(regs_124_clock),
    .reset(regs_124_reset),
    .io_in(regs_124_io_in),
    .io_reset(regs_124_io_reset),
    .io_out(regs_124_io_out),
    .io_enable(regs_124_io_enable)
  );
  FringeFF regs_125 ( // @[RegFile.scala 66:20:@43638.4]
    .clock(regs_125_clock),
    .reset(regs_125_reset),
    .io_in(regs_125_io_in),
    .io_reset(regs_125_io_reset),
    .io_out(regs_125_io_out),
    .io_enable(regs_125_io_enable)
  );
  FringeFF regs_126 ( // @[RegFile.scala 66:20:@43652.4]
    .clock(regs_126_clock),
    .reset(regs_126_reset),
    .io_in(regs_126_io_in),
    .io_reset(regs_126_io_reset),
    .io_out(regs_126_io_out),
    .io_enable(regs_126_io_enable)
  );
  FringeFF regs_127 ( // @[RegFile.scala 66:20:@43666.4]
    .clock(regs_127_clock),
    .reset(regs_127_reset),
    .io_in(regs_127_io_in),
    .io_reset(regs_127_io_reset),
    .io_out(regs_127_io_out),
    .io_enable(regs_127_io_enable)
  );
  FringeFF regs_128 ( // @[RegFile.scala 66:20:@43680.4]
    .clock(regs_128_clock),
    .reset(regs_128_reset),
    .io_in(regs_128_io_in),
    .io_reset(regs_128_io_reset),
    .io_out(regs_128_io_out),
    .io_enable(regs_128_io_enable)
  );
  FringeFF regs_129 ( // @[RegFile.scala 66:20:@43694.4]
    .clock(regs_129_clock),
    .reset(regs_129_reset),
    .io_in(regs_129_io_in),
    .io_reset(regs_129_io_reset),
    .io_out(regs_129_io_out),
    .io_enable(regs_129_io_enable)
  );
  FringeFF regs_130 ( // @[RegFile.scala 66:20:@43708.4]
    .clock(regs_130_clock),
    .reset(regs_130_reset),
    .io_in(regs_130_io_in),
    .io_reset(regs_130_io_reset),
    .io_out(regs_130_io_out),
    .io_enable(regs_130_io_enable)
  );
  FringeFF regs_131 ( // @[RegFile.scala 66:20:@43722.4]
    .clock(regs_131_clock),
    .reset(regs_131_reset),
    .io_in(regs_131_io_in),
    .io_reset(regs_131_io_reset),
    .io_out(regs_131_io_out),
    .io_enable(regs_131_io_enable)
  );
  FringeFF regs_132 ( // @[RegFile.scala 66:20:@43736.4]
    .clock(regs_132_clock),
    .reset(regs_132_reset),
    .io_in(regs_132_io_in),
    .io_reset(regs_132_io_reset),
    .io_out(regs_132_io_out),
    .io_enable(regs_132_io_enable)
  );
  FringeFF regs_133 ( // @[RegFile.scala 66:20:@43750.4]
    .clock(regs_133_clock),
    .reset(regs_133_reset),
    .io_in(regs_133_io_in),
    .io_reset(regs_133_io_reset),
    .io_out(regs_133_io_out),
    .io_enable(regs_133_io_enable)
  );
  FringeFF regs_134 ( // @[RegFile.scala 66:20:@43764.4]
    .clock(regs_134_clock),
    .reset(regs_134_reset),
    .io_in(regs_134_io_in),
    .io_reset(regs_134_io_reset),
    .io_out(regs_134_io_out),
    .io_enable(regs_134_io_enable)
  );
  FringeFF regs_135 ( // @[RegFile.scala 66:20:@43778.4]
    .clock(regs_135_clock),
    .reset(regs_135_reset),
    .io_in(regs_135_io_in),
    .io_reset(regs_135_io_reset),
    .io_out(regs_135_io_out),
    .io_enable(regs_135_io_enable)
  );
  FringeFF regs_136 ( // @[RegFile.scala 66:20:@43792.4]
    .clock(regs_136_clock),
    .reset(regs_136_reset),
    .io_in(regs_136_io_in),
    .io_reset(regs_136_io_reset),
    .io_out(regs_136_io_out),
    .io_enable(regs_136_io_enable)
  );
  FringeFF regs_137 ( // @[RegFile.scala 66:20:@43806.4]
    .clock(regs_137_clock),
    .reset(regs_137_reset),
    .io_in(regs_137_io_in),
    .io_reset(regs_137_io_reset),
    .io_out(regs_137_io_out),
    .io_enable(regs_137_io_enable)
  );
  FringeFF regs_138 ( // @[RegFile.scala 66:20:@43820.4]
    .clock(regs_138_clock),
    .reset(regs_138_reset),
    .io_in(regs_138_io_in),
    .io_reset(regs_138_io_reset),
    .io_out(regs_138_io_out),
    .io_enable(regs_138_io_enable)
  );
  FringeFF regs_139 ( // @[RegFile.scala 66:20:@43834.4]
    .clock(regs_139_clock),
    .reset(regs_139_reset),
    .io_in(regs_139_io_in),
    .io_reset(regs_139_io_reset),
    .io_out(regs_139_io_out),
    .io_enable(regs_139_io_enable)
  );
  FringeFF regs_140 ( // @[RegFile.scala 66:20:@43848.4]
    .clock(regs_140_clock),
    .reset(regs_140_reset),
    .io_in(regs_140_io_in),
    .io_reset(regs_140_io_reset),
    .io_out(regs_140_io_out),
    .io_enable(regs_140_io_enable)
  );
  FringeFF regs_141 ( // @[RegFile.scala 66:20:@43862.4]
    .clock(regs_141_clock),
    .reset(regs_141_reset),
    .io_in(regs_141_io_in),
    .io_reset(regs_141_io_reset),
    .io_out(regs_141_io_out),
    .io_enable(regs_141_io_enable)
  );
  FringeFF regs_142 ( // @[RegFile.scala 66:20:@43876.4]
    .clock(regs_142_clock),
    .reset(regs_142_reset),
    .io_in(regs_142_io_in),
    .io_reset(regs_142_io_reset),
    .io_out(regs_142_io_out),
    .io_enable(regs_142_io_enable)
  );
  FringeFF regs_143 ( // @[RegFile.scala 66:20:@43890.4]
    .clock(regs_143_clock),
    .reset(regs_143_reset),
    .io_in(regs_143_io_in),
    .io_reset(regs_143_io_reset),
    .io_out(regs_143_io_out),
    .io_enable(regs_143_io_enable)
  );
  FringeFF regs_144 ( // @[RegFile.scala 66:20:@43904.4]
    .clock(regs_144_clock),
    .reset(regs_144_reset),
    .io_in(regs_144_io_in),
    .io_reset(regs_144_io_reset),
    .io_out(regs_144_io_out),
    .io_enable(regs_144_io_enable)
  );
  FringeFF regs_145 ( // @[RegFile.scala 66:20:@43918.4]
    .clock(regs_145_clock),
    .reset(regs_145_reset),
    .io_in(regs_145_io_in),
    .io_reset(regs_145_io_reset),
    .io_out(regs_145_io_out),
    .io_enable(regs_145_io_enable)
  );
  FringeFF regs_146 ( // @[RegFile.scala 66:20:@43932.4]
    .clock(regs_146_clock),
    .reset(regs_146_reset),
    .io_in(regs_146_io_in),
    .io_reset(regs_146_io_reset),
    .io_out(regs_146_io_out),
    .io_enable(regs_146_io_enable)
  );
  FringeFF regs_147 ( // @[RegFile.scala 66:20:@43946.4]
    .clock(regs_147_clock),
    .reset(regs_147_reset),
    .io_in(regs_147_io_in),
    .io_reset(regs_147_io_reset),
    .io_out(regs_147_io_out),
    .io_enable(regs_147_io_enable)
  );
  FringeFF regs_148 ( // @[RegFile.scala 66:20:@43960.4]
    .clock(regs_148_clock),
    .reset(regs_148_reset),
    .io_in(regs_148_io_in),
    .io_reset(regs_148_io_reset),
    .io_out(regs_148_io_out),
    .io_enable(regs_148_io_enable)
  );
  FringeFF regs_149 ( // @[RegFile.scala 66:20:@43974.4]
    .clock(regs_149_clock),
    .reset(regs_149_reset),
    .io_in(regs_149_io_in),
    .io_reset(regs_149_io_reset),
    .io_out(regs_149_io_out),
    .io_enable(regs_149_io_enable)
  );
  FringeFF regs_150 ( // @[RegFile.scala 66:20:@43988.4]
    .clock(regs_150_clock),
    .reset(regs_150_reset),
    .io_in(regs_150_io_in),
    .io_reset(regs_150_io_reset),
    .io_out(regs_150_io_out),
    .io_enable(regs_150_io_enable)
  );
  FringeFF regs_151 ( // @[RegFile.scala 66:20:@44002.4]
    .clock(regs_151_clock),
    .reset(regs_151_reset),
    .io_in(regs_151_io_in),
    .io_reset(regs_151_io_reset),
    .io_out(regs_151_io_out),
    .io_enable(regs_151_io_enable)
  );
  FringeFF regs_152 ( // @[RegFile.scala 66:20:@44016.4]
    .clock(regs_152_clock),
    .reset(regs_152_reset),
    .io_in(regs_152_io_in),
    .io_reset(regs_152_io_reset),
    .io_out(regs_152_io_out),
    .io_enable(regs_152_io_enable)
  );
  FringeFF regs_153 ( // @[RegFile.scala 66:20:@44030.4]
    .clock(regs_153_clock),
    .reset(regs_153_reset),
    .io_in(regs_153_io_in),
    .io_reset(regs_153_io_reset),
    .io_out(regs_153_io_out),
    .io_enable(regs_153_io_enable)
  );
  FringeFF regs_154 ( // @[RegFile.scala 66:20:@44044.4]
    .clock(regs_154_clock),
    .reset(regs_154_reset),
    .io_in(regs_154_io_in),
    .io_reset(regs_154_io_reset),
    .io_out(regs_154_io_out),
    .io_enable(regs_154_io_enable)
  );
  FringeFF regs_155 ( // @[RegFile.scala 66:20:@44058.4]
    .clock(regs_155_clock),
    .reset(regs_155_reset),
    .io_in(regs_155_io_in),
    .io_reset(regs_155_io_reset),
    .io_out(regs_155_io_out),
    .io_enable(regs_155_io_enable)
  );
  FringeFF regs_156 ( // @[RegFile.scala 66:20:@44072.4]
    .clock(regs_156_clock),
    .reset(regs_156_reset),
    .io_in(regs_156_io_in),
    .io_reset(regs_156_io_reset),
    .io_out(regs_156_io_out),
    .io_enable(regs_156_io_enable)
  );
  FringeFF regs_157 ( // @[RegFile.scala 66:20:@44086.4]
    .clock(regs_157_clock),
    .reset(regs_157_reset),
    .io_in(regs_157_io_in),
    .io_reset(regs_157_io_reset),
    .io_out(regs_157_io_out),
    .io_enable(regs_157_io_enable)
  );
  FringeFF regs_158 ( // @[RegFile.scala 66:20:@44100.4]
    .clock(regs_158_clock),
    .reset(regs_158_reset),
    .io_in(regs_158_io_in),
    .io_reset(regs_158_io_reset),
    .io_out(regs_158_io_out),
    .io_enable(regs_158_io_enable)
  );
  FringeFF regs_159 ( // @[RegFile.scala 66:20:@44114.4]
    .clock(regs_159_clock),
    .reset(regs_159_reset),
    .io_in(regs_159_io_in),
    .io_reset(regs_159_io_reset),
    .io_out(regs_159_io_out),
    .io_enable(regs_159_io_enable)
  );
  FringeFF regs_160 ( // @[RegFile.scala 66:20:@44128.4]
    .clock(regs_160_clock),
    .reset(regs_160_reset),
    .io_in(regs_160_io_in),
    .io_reset(regs_160_io_reset),
    .io_out(regs_160_io_out),
    .io_enable(regs_160_io_enable)
  );
  FringeFF regs_161 ( // @[RegFile.scala 66:20:@44142.4]
    .clock(regs_161_clock),
    .reset(regs_161_reset),
    .io_in(regs_161_io_in),
    .io_reset(regs_161_io_reset),
    .io_out(regs_161_io_out),
    .io_enable(regs_161_io_enable)
  );
  FringeFF regs_162 ( // @[RegFile.scala 66:20:@44156.4]
    .clock(regs_162_clock),
    .reset(regs_162_reset),
    .io_in(regs_162_io_in),
    .io_reset(regs_162_io_reset),
    .io_out(regs_162_io_out),
    .io_enable(regs_162_io_enable)
  );
  FringeFF regs_163 ( // @[RegFile.scala 66:20:@44170.4]
    .clock(regs_163_clock),
    .reset(regs_163_reset),
    .io_in(regs_163_io_in),
    .io_reset(regs_163_io_reset),
    .io_out(regs_163_io_out),
    .io_enable(regs_163_io_enable)
  );
  FringeFF regs_164 ( // @[RegFile.scala 66:20:@44184.4]
    .clock(regs_164_clock),
    .reset(regs_164_reset),
    .io_in(regs_164_io_in),
    .io_reset(regs_164_io_reset),
    .io_out(regs_164_io_out),
    .io_enable(regs_164_io_enable)
  );
  FringeFF regs_165 ( // @[RegFile.scala 66:20:@44198.4]
    .clock(regs_165_clock),
    .reset(regs_165_reset),
    .io_in(regs_165_io_in),
    .io_reset(regs_165_io_reset),
    .io_out(regs_165_io_out),
    .io_enable(regs_165_io_enable)
  );
  FringeFF regs_166 ( // @[RegFile.scala 66:20:@44212.4]
    .clock(regs_166_clock),
    .reset(regs_166_reset),
    .io_in(regs_166_io_in),
    .io_reset(regs_166_io_reset),
    .io_out(regs_166_io_out),
    .io_enable(regs_166_io_enable)
  );
  FringeFF regs_167 ( // @[RegFile.scala 66:20:@44226.4]
    .clock(regs_167_clock),
    .reset(regs_167_reset),
    .io_in(regs_167_io_in),
    .io_reset(regs_167_io_reset),
    .io_out(regs_167_io_out),
    .io_enable(regs_167_io_enable)
  );
  FringeFF regs_168 ( // @[RegFile.scala 66:20:@44240.4]
    .clock(regs_168_clock),
    .reset(regs_168_reset),
    .io_in(regs_168_io_in),
    .io_reset(regs_168_io_reset),
    .io_out(regs_168_io_out),
    .io_enable(regs_168_io_enable)
  );
  FringeFF regs_169 ( // @[RegFile.scala 66:20:@44254.4]
    .clock(regs_169_clock),
    .reset(regs_169_reset),
    .io_in(regs_169_io_in),
    .io_reset(regs_169_io_reset),
    .io_out(regs_169_io_out),
    .io_enable(regs_169_io_enable)
  );
  FringeFF regs_170 ( // @[RegFile.scala 66:20:@44268.4]
    .clock(regs_170_clock),
    .reset(regs_170_reset),
    .io_in(regs_170_io_in),
    .io_reset(regs_170_io_reset),
    .io_out(regs_170_io_out),
    .io_enable(regs_170_io_enable)
  );
  FringeFF regs_171 ( // @[RegFile.scala 66:20:@44282.4]
    .clock(regs_171_clock),
    .reset(regs_171_reset),
    .io_in(regs_171_io_in),
    .io_reset(regs_171_io_reset),
    .io_out(regs_171_io_out),
    .io_enable(regs_171_io_enable)
  );
  FringeFF regs_172 ( // @[RegFile.scala 66:20:@44296.4]
    .clock(regs_172_clock),
    .reset(regs_172_reset),
    .io_in(regs_172_io_in),
    .io_reset(regs_172_io_reset),
    .io_out(regs_172_io_out),
    .io_enable(regs_172_io_enable)
  );
  FringeFF regs_173 ( // @[RegFile.scala 66:20:@44310.4]
    .clock(regs_173_clock),
    .reset(regs_173_reset),
    .io_in(regs_173_io_in),
    .io_reset(regs_173_io_reset),
    .io_out(regs_173_io_out),
    .io_enable(regs_173_io_enable)
  );
  FringeFF regs_174 ( // @[RegFile.scala 66:20:@44324.4]
    .clock(regs_174_clock),
    .reset(regs_174_reset),
    .io_in(regs_174_io_in),
    .io_reset(regs_174_io_reset),
    .io_out(regs_174_io_out),
    .io_enable(regs_174_io_enable)
  );
  FringeFF regs_175 ( // @[RegFile.scala 66:20:@44338.4]
    .clock(regs_175_clock),
    .reset(regs_175_reset),
    .io_in(regs_175_io_in),
    .io_reset(regs_175_io_reset),
    .io_out(regs_175_io_out),
    .io_enable(regs_175_io_enable)
  );
  FringeFF regs_176 ( // @[RegFile.scala 66:20:@44352.4]
    .clock(regs_176_clock),
    .reset(regs_176_reset),
    .io_in(regs_176_io_in),
    .io_reset(regs_176_io_reset),
    .io_out(regs_176_io_out),
    .io_enable(regs_176_io_enable)
  );
  FringeFF regs_177 ( // @[RegFile.scala 66:20:@44366.4]
    .clock(regs_177_clock),
    .reset(regs_177_reset),
    .io_in(regs_177_io_in),
    .io_reset(regs_177_io_reset),
    .io_out(regs_177_io_out),
    .io_enable(regs_177_io_enable)
  );
  FringeFF regs_178 ( // @[RegFile.scala 66:20:@44380.4]
    .clock(regs_178_clock),
    .reset(regs_178_reset),
    .io_in(regs_178_io_in),
    .io_reset(regs_178_io_reset),
    .io_out(regs_178_io_out),
    .io_enable(regs_178_io_enable)
  );
  FringeFF regs_179 ( // @[RegFile.scala 66:20:@44394.4]
    .clock(regs_179_clock),
    .reset(regs_179_reset),
    .io_in(regs_179_io_in),
    .io_reset(regs_179_io_reset),
    .io_out(regs_179_io_out),
    .io_enable(regs_179_io_enable)
  );
  FringeFF regs_180 ( // @[RegFile.scala 66:20:@44408.4]
    .clock(regs_180_clock),
    .reset(regs_180_reset),
    .io_in(regs_180_io_in),
    .io_reset(regs_180_io_reset),
    .io_out(regs_180_io_out),
    .io_enable(regs_180_io_enable)
  );
  FringeFF regs_181 ( // @[RegFile.scala 66:20:@44422.4]
    .clock(regs_181_clock),
    .reset(regs_181_reset),
    .io_in(regs_181_io_in),
    .io_reset(regs_181_io_reset),
    .io_out(regs_181_io_out),
    .io_enable(regs_181_io_enable)
  );
  FringeFF regs_182 ( // @[RegFile.scala 66:20:@44436.4]
    .clock(regs_182_clock),
    .reset(regs_182_reset),
    .io_in(regs_182_io_in),
    .io_reset(regs_182_io_reset),
    .io_out(regs_182_io_out),
    .io_enable(regs_182_io_enable)
  );
  FringeFF regs_183 ( // @[RegFile.scala 66:20:@44450.4]
    .clock(regs_183_clock),
    .reset(regs_183_reset),
    .io_in(regs_183_io_in),
    .io_reset(regs_183_io_reset),
    .io_out(regs_183_io_out),
    .io_enable(regs_183_io_enable)
  );
  FringeFF regs_184 ( // @[RegFile.scala 66:20:@44464.4]
    .clock(regs_184_clock),
    .reset(regs_184_reset),
    .io_in(regs_184_io_in),
    .io_reset(regs_184_io_reset),
    .io_out(regs_184_io_out),
    .io_enable(regs_184_io_enable)
  );
  FringeFF regs_185 ( // @[RegFile.scala 66:20:@44478.4]
    .clock(regs_185_clock),
    .reset(regs_185_reset),
    .io_in(regs_185_io_in),
    .io_reset(regs_185_io_reset),
    .io_out(regs_185_io_out),
    .io_enable(regs_185_io_enable)
  );
  FringeFF regs_186 ( // @[RegFile.scala 66:20:@44492.4]
    .clock(regs_186_clock),
    .reset(regs_186_reset),
    .io_in(regs_186_io_in),
    .io_reset(regs_186_io_reset),
    .io_out(regs_186_io_out),
    .io_enable(regs_186_io_enable)
  );
  FringeFF regs_187 ( // @[RegFile.scala 66:20:@44506.4]
    .clock(regs_187_clock),
    .reset(regs_187_reset),
    .io_in(regs_187_io_in),
    .io_reset(regs_187_io_reset),
    .io_out(regs_187_io_out),
    .io_enable(regs_187_io_enable)
  );
  FringeFF regs_188 ( // @[RegFile.scala 66:20:@44520.4]
    .clock(regs_188_clock),
    .reset(regs_188_reset),
    .io_in(regs_188_io_in),
    .io_reset(regs_188_io_reset),
    .io_out(regs_188_io_out),
    .io_enable(regs_188_io_enable)
  );
  FringeFF regs_189 ( // @[RegFile.scala 66:20:@44534.4]
    .clock(regs_189_clock),
    .reset(regs_189_reset),
    .io_in(regs_189_io_in),
    .io_reset(regs_189_io_reset),
    .io_out(regs_189_io_out),
    .io_enable(regs_189_io_enable)
  );
  FringeFF regs_190 ( // @[RegFile.scala 66:20:@44548.4]
    .clock(regs_190_clock),
    .reset(regs_190_reset),
    .io_in(regs_190_io_in),
    .io_reset(regs_190_io_reset),
    .io_out(regs_190_io_out),
    .io_enable(regs_190_io_enable)
  );
  FringeFF regs_191 ( // @[RegFile.scala 66:20:@44562.4]
    .clock(regs_191_clock),
    .reset(regs_191_reset),
    .io_in(regs_191_io_in),
    .io_reset(regs_191_io_reset),
    .io_out(regs_191_io_out),
    .io_enable(regs_191_io_enable)
  );
  FringeFF regs_192 ( // @[RegFile.scala 66:20:@44576.4]
    .clock(regs_192_clock),
    .reset(regs_192_reset),
    .io_in(regs_192_io_in),
    .io_reset(regs_192_io_reset),
    .io_out(regs_192_io_out),
    .io_enable(regs_192_io_enable)
  );
  FringeFF regs_193 ( // @[RegFile.scala 66:20:@44590.4]
    .clock(regs_193_clock),
    .reset(regs_193_reset),
    .io_in(regs_193_io_in),
    .io_reset(regs_193_io_reset),
    .io_out(regs_193_io_out),
    .io_enable(regs_193_io_enable)
  );
  FringeFF regs_194 ( // @[RegFile.scala 66:20:@44604.4]
    .clock(regs_194_clock),
    .reset(regs_194_reset),
    .io_in(regs_194_io_in),
    .io_reset(regs_194_io_reset),
    .io_out(regs_194_io_out),
    .io_enable(regs_194_io_enable)
  );
  FringeFF regs_195 ( // @[RegFile.scala 66:20:@44618.4]
    .clock(regs_195_clock),
    .reset(regs_195_reset),
    .io_in(regs_195_io_in),
    .io_reset(regs_195_io_reset),
    .io_out(regs_195_io_out),
    .io_enable(regs_195_io_enable)
  );
  FringeFF regs_196 ( // @[RegFile.scala 66:20:@44632.4]
    .clock(regs_196_clock),
    .reset(regs_196_reset),
    .io_in(regs_196_io_in),
    .io_reset(regs_196_io_reset),
    .io_out(regs_196_io_out),
    .io_enable(regs_196_io_enable)
  );
  FringeFF regs_197 ( // @[RegFile.scala 66:20:@44646.4]
    .clock(regs_197_clock),
    .reset(regs_197_reset),
    .io_in(regs_197_io_in),
    .io_reset(regs_197_io_reset),
    .io_out(regs_197_io_out),
    .io_enable(regs_197_io_enable)
  );
  FringeFF regs_198 ( // @[RegFile.scala 66:20:@44660.4]
    .clock(regs_198_clock),
    .reset(regs_198_reset),
    .io_in(regs_198_io_in),
    .io_reset(regs_198_io_reset),
    .io_out(regs_198_io_out),
    .io_enable(regs_198_io_enable)
  );
  FringeFF regs_199 ( // @[RegFile.scala 66:20:@44674.4]
    .clock(regs_199_clock),
    .reset(regs_199_reset),
    .io_in(regs_199_io_in),
    .io_reset(regs_199_io_reset),
    .io_out(regs_199_io_out),
    .io_enable(regs_199_io_enable)
  );
  FringeFF regs_200 ( // @[RegFile.scala 66:20:@44688.4]
    .clock(regs_200_clock),
    .reset(regs_200_reset),
    .io_in(regs_200_io_in),
    .io_reset(regs_200_io_reset),
    .io_out(regs_200_io_out),
    .io_enable(regs_200_io_enable)
  );
  FringeFF regs_201 ( // @[RegFile.scala 66:20:@44702.4]
    .clock(regs_201_clock),
    .reset(regs_201_reset),
    .io_in(regs_201_io_in),
    .io_reset(regs_201_io_reset),
    .io_out(regs_201_io_out),
    .io_enable(regs_201_io_enable)
  );
  FringeFF regs_202 ( // @[RegFile.scala 66:20:@44716.4]
    .clock(regs_202_clock),
    .reset(regs_202_reset),
    .io_in(regs_202_io_in),
    .io_reset(regs_202_io_reset),
    .io_out(regs_202_io_out),
    .io_enable(regs_202_io_enable)
  );
  FringeFF regs_203 ( // @[RegFile.scala 66:20:@44730.4]
    .clock(regs_203_clock),
    .reset(regs_203_reset),
    .io_in(regs_203_io_in),
    .io_reset(regs_203_io_reset),
    .io_out(regs_203_io_out),
    .io_enable(regs_203_io_enable)
  );
  FringeFF regs_204 ( // @[RegFile.scala 66:20:@44744.4]
    .clock(regs_204_clock),
    .reset(regs_204_reset),
    .io_in(regs_204_io_in),
    .io_reset(regs_204_io_reset),
    .io_out(regs_204_io_out),
    .io_enable(regs_204_io_enable)
  );
  FringeFF regs_205 ( // @[RegFile.scala 66:20:@44758.4]
    .clock(regs_205_clock),
    .reset(regs_205_reset),
    .io_in(regs_205_io_in),
    .io_reset(regs_205_io_reset),
    .io_out(regs_205_io_out),
    .io_enable(regs_205_io_enable)
  );
  FringeFF regs_206 ( // @[RegFile.scala 66:20:@44772.4]
    .clock(regs_206_clock),
    .reset(regs_206_reset),
    .io_in(regs_206_io_in),
    .io_reset(regs_206_io_reset),
    .io_out(regs_206_io_out),
    .io_enable(regs_206_io_enable)
  );
  FringeFF regs_207 ( // @[RegFile.scala 66:20:@44786.4]
    .clock(regs_207_clock),
    .reset(regs_207_reset),
    .io_in(regs_207_io_in),
    .io_reset(regs_207_io_reset),
    .io_out(regs_207_io_out),
    .io_enable(regs_207_io_enable)
  );
  FringeFF regs_208 ( // @[RegFile.scala 66:20:@44800.4]
    .clock(regs_208_clock),
    .reset(regs_208_reset),
    .io_in(regs_208_io_in),
    .io_reset(regs_208_io_reset),
    .io_out(regs_208_io_out),
    .io_enable(regs_208_io_enable)
  );
  FringeFF regs_209 ( // @[RegFile.scala 66:20:@44814.4]
    .clock(regs_209_clock),
    .reset(regs_209_reset),
    .io_in(regs_209_io_in),
    .io_reset(regs_209_io_reset),
    .io_out(regs_209_io_out),
    .io_enable(regs_209_io_enable)
  );
  FringeFF regs_210 ( // @[RegFile.scala 66:20:@44828.4]
    .clock(regs_210_clock),
    .reset(regs_210_reset),
    .io_in(regs_210_io_in),
    .io_reset(regs_210_io_reset),
    .io_out(regs_210_io_out),
    .io_enable(regs_210_io_enable)
  );
  FringeFF regs_211 ( // @[RegFile.scala 66:20:@44842.4]
    .clock(regs_211_clock),
    .reset(regs_211_reset),
    .io_in(regs_211_io_in),
    .io_reset(regs_211_io_reset),
    .io_out(regs_211_io_out),
    .io_enable(regs_211_io_enable)
  );
  FringeFF regs_212 ( // @[RegFile.scala 66:20:@44856.4]
    .clock(regs_212_clock),
    .reset(regs_212_reset),
    .io_in(regs_212_io_in),
    .io_reset(regs_212_io_reset),
    .io_out(regs_212_io_out),
    .io_enable(regs_212_io_enable)
  );
  FringeFF regs_213 ( // @[RegFile.scala 66:20:@44870.4]
    .clock(regs_213_clock),
    .reset(regs_213_reset),
    .io_in(regs_213_io_in),
    .io_reset(regs_213_io_reset),
    .io_out(regs_213_io_out),
    .io_enable(regs_213_io_enable)
  );
  FringeFF regs_214 ( // @[RegFile.scala 66:20:@44884.4]
    .clock(regs_214_clock),
    .reset(regs_214_reset),
    .io_in(regs_214_io_in),
    .io_reset(regs_214_io_reset),
    .io_out(regs_214_io_out),
    .io_enable(regs_214_io_enable)
  );
  FringeFF regs_215 ( // @[RegFile.scala 66:20:@44898.4]
    .clock(regs_215_clock),
    .reset(regs_215_reset),
    .io_in(regs_215_io_in),
    .io_reset(regs_215_io_reset),
    .io_out(regs_215_io_out),
    .io_enable(regs_215_io_enable)
  );
  FringeFF regs_216 ( // @[RegFile.scala 66:20:@44912.4]
    .clock(regs_216_clock),
    .reset(regs_216_reset),
    .io_in(regs_216_io_in),
    .io_reset(regs_216_io_reset),
    .io_out(regs_216_io_out),
    .io_enable(regs_216_io_enable)
  );
  FringeFF regs_217 ( // @[RegFile.scala 66:20:@44926.4]
    .clock(regs_217_clock),
    .reset(regs_217_reset),
    .io_in(regs_217_io_in),
    .io_reset(regs_217_io_reset),
    .io_out(regs_217_io_out),
    .io_enable(regs_217_io_enable)
  );
  FringeFF regs_218 ( // @[RegFile.scala 66:20:@44940.4]
    .clock(regs_218_clock),
    .reset(regs_218_reset),
    .io_in(regs_218_io_in),
    .io_reset(regs_218_io_reset),
    .io_out(regs_218_io_out),
    .io_enable(regs_218_io_enable)
  );
  FringeFF regs_219 ( // @[RegFile.scala 66:20:@44954.4]
    .clock(regs_219_clock),
    .reset(regs_219_reset),
    .io_in(regs_219_io_in),
    .io_reset(regs_219_io_reset),
    .io_out(regs_219_io_out),
    .io_enable(regs_219_io_enable)
  );
  FringeFF regs_220 ( // @[RegFile.scala 66:20:@44968.4]
    .clock(regs_220_clock),
    .reset(regs_220_reset),
    .io_in(regs_220_io_in),
    .io_reset(regs_220_io_reset),
    .io_out(regs_220_io_out),
    .io_enable(regs_220_io_enable)
  );
  FringeFF regs_221 ( // @[RegFile.scala 66:20:@44982.4]
    .clock(regs_221_clock),
    .reset(regs_221_reset),
    .io_in(regs_221_io_in),
    .io_reset(regs_221_io_reset),
    .io_out(regs_221_io_out),
    .io_enable(regs_221_io_enable)
  );
  FringeFF regs_222 ( // @[RegFile.scala 66:20:@44996.4]
    .clock(regs_222_clock),
    .reset(regs_222_reset),
    .io_in(regs_222_io_in),
    .io_reset(regs_222_io_reset),
    .io_out(regs_222_io_out),
    .io_enable(regs_222_io_enable)
  );
  FringeFF regs_223 ( // @[RegFile.scala 66:20:@45010.4]
    .clock(regs_223_clock),
    .reset(regs_223_reset),
    .io_in(regs_223_io_in),
    .io_reset(regs_223_io_reset),
    .io_out(regs_223_io_out),
    .io_enable(regs_223_io_enable)
  );
  FringeFF regs_224 ( // @[RegFile.scala 66:20:@45024.4]
    .clock(regs_224_clock),
    .reset(regs_224_reset),
    .io_in(regs_224_io_in),
    .io_reset(regs_224_io_reset),
    .io_out(regs_224_io_out),
    .io_enable(regs_224_io_enable)
  );
  FringeFF regs_225 ( // @[RegFile.scala 66:20:@45038.4]
    .clock(regs_225_clock),
    .reset(regs_225_reset),
    .io_in(regs_225_io_in),
    .io_reset(regs_225_io_reset),
    .io_out(regs_225_io_out),
    .io_enable(regs_225_io_enable)
  );
  FringeFF regs_226 ( // @[RegFile.scala 66:20:@45052.4]
    .clock(regs_226_clock),
    .reset(regs_226_reset),
    .io_in(regs_226_io_in),
    .io_reset(regs_226_io_reset),
    .io_out(regs_226_io_out),
    .io_enable(regs_226_io_enable)
  );
  FringeFF regs_227 ( // @[RegFile.scala 66:20:@45066.4]
    .clock(regs_227_clock),
    .reset(regs_227_reset),
    .io_in(regs_227_io_in),
    .io_reset(regs_227_io_reset),
    .io_out(regs_227_io_out),
    .io_enable(regs_227_io_enable)
  );
  FringeFF regs_228 ( // @[RegFile.scala 66:20:@45080.4]
    .clock(regs_228_clock),
    .reset(regs_228_reset),
    .io_in(regs_228_io_in),
    .io_reset(regs_228_io_reset),
    .io_out(regs_228_io_out),
    .io_enable(regs_228_io_enable)
  );
  FringeFF regs_229 ( // @[RegFile.scala 66:20:@45094.4]
    .clock(regs_229_clock),
    .reset(regs_229_reset),
    .io_in(regs_229_io_in),
    .io_reset(regs_229_io_reset),
    .io_out(regs_229_io_out),
    .io_enable(regs_229_io_enable)
  );
  FringeFF regs_230 ( // @[RegFile.scala 66:20:@45108.4]
    .clock(regs_230_clock),
    .reset(regs_230_reset),
    .io_in(regs_230_io_in),
    .io_reset(regs_230_io_reset),
    .io_out(regs_230_io_out),
    .io_enable(regs_230_io_enable)
  );
  FringeFF regs_231 ( // @[RegFile.scala 66:20:@45122.4]
    .clock(regs_231_clock),
    .reset(regs_231_reset),
    .io_in(regs_231_io_in),
    .io_reset(regs_231_io_reset),
    .io_out(regs_231_io_out),
    .io_enable(regs_231_io_enable)
  );
  FringeFF regs_232 ( // @[RegFile.scala 66:20:@45136.4]
    .clock(regs_232_clock),
    .reset(regs_232_reset),
    .io_in(regs_232_io_in),
    .io_reset(regs_232_io_reset),
    .io_out(regs_232_io_out),
    .io_enable(regs_232_io_enable)
  );
  FringeFF regs_233 ( // @[RegFile.scala 66:20:@45150.4]
    .clock(regs_233_clock),
    .reset(regs_233_reset),
    .io_in(regs_233_io_in),
    .io_reset(regs_233_io_reset),
    .io_out(regs_233_io_out),
    .io_enable(regs_233_io_enable)
  );
  FringeFF regs_234 ( // @[RegFile.scala 66:20:@45164.4]
    .clock(regs_234_clock),
    .reset(regs_234_reset),
    .io_in(regs_234_io_in),
    .io_reset(regs_234_io_reset),
    .io_out(regs_234_io_out),
    .io_enable(regs_234_io_enable)
  );
  FringeFF regs_235 ( // @[RegFile.scala 66:20:@45178.4]
    .clock(regs_235_clock),
    .reset(regs_235_reset),
    .io_in(regs_235_io_in),
    .io_reset(regs_235_io_reset),
    .io_out(regs_235_io_out),
    .io_enable(regs_235_io_enable)
  );
  FringeFF regs_236 ( // @[RegFile.scala 66:20:@45192.4]
    .clock(regs_236_clock),
    .reset(regs_236_reset),
    .io_in(regs_236_io_in),
    .io_reset(regs_236_io_reset),
    .io_out(regs_236_io_out),
    .io_enable(regs_236_io_enable)
  );
  FringeFF regs_237 ( // @[RegFile.scala 66:20:@45206.4]
    .clock(regs_237_clock),
    .reset(regs_237_reset),
    .io_in(regs_237_io_in),
    .io_reset(regs_237_io_reset),
    .io_out(regs_237_io_out),
    .io_enable(regs_237_io_enable)
  );
  FringeFF regs_238 ( // @[RegFile.scala 66:20:@45220.4]
    .clock(regs_238_clock),
    .reset(regs_238_reset),
    .io_in(regs_238_io_in),
    .io_reset(regs_238_io_reset),
    .io_out(regs_238_io_out),
    .io_enable(regs_238_io_enable)
  );
  FringeFF regs_239 ( // @[RegFile.scala 66:20:@45234.4]
    .clock(regs_239_clock),
    .reset(regs_239_reset),
    .io_in(regs_239_io_in),
    .io_reset(regs_239_io_reset),
    .io_out(regs_239_io_out),
    .io_enable(regs_239_io_enable)
  );
  FringeFF regs_240 ( // @[RegFile.scala 66:20:@45248.4]
    .clock(regs_240_clock),
    .reset(regs_240_reset),
    .io_in(regs_240_io_in),
    .io_reset(regs_240_io_reset),
    .io_out(regs_240_io_out),
    .io_enable(regs_240_io_enable)
  );
  FringeFF regs_241 ( // @[RegFile.scala 66:20:@45262.4]
    .clock(regs_241_clock),
    .reset(regs_241_reset),
    .io_in(regs_241_io_in),
    .io_reset(regs_241_io_reset),
    .io_out(regs_241_io_out),
    .io_enable(regs_241_io_enable)
  );
  FringeFF regs_242 ( // @[RegFile.scala 66:20:@45276.4]
    .clock(regs_242_clock),
    .reset(regs_242_reset),
    .io_in(regs_242_io_in),
    .io_reset(regs_242_io_reset),
    .io_out(regs_242_io_out),
    .io_enable(regs_242_io_enable)
  );
  FringeFF regs_243 ( // @[RegFile.scala 66:20:@45290.4]
    .clock(regs_243_clock),
    .reset(regs_243_reset),
    .io_in(regs_243_io_in),
    .io_reset(regs_243_io_reset),
    .io_out(regs_243_io_out),
    .io_enable(regs_243_io_enable)
  );
  FringeFF regs_244 ( // @[RegFile.scala 66:20:@45304.4]
    .clock(regs_244_clock),
    .reset(regs_244_reset),
    .io_in(regs_244_io_in),
    .io_reset(regs_244_io_reset),
    .io_out(regs_244_io_out),
    .io_enable(regs_244_io_enable)
  );
  FringeFF regs_245 ( // @[RegFile.scala 66:20:@45318.4]
    .clock(regs_245_clock),
    .reset(regs_245_reset),
    .io_in(regs_245_io_in),
    .io_reset(regs_245_io_reset),
    .io_out(regs_245_io_out),
    .io_enable(regs_245_io_enable)
  );
  FringeFF regs_246 ( // @[RegFile.scala 66:20:@45332.4]
    .clock(regs_246_clock),
    .reset(regs_246_reset),
    .io_in(regs_246_io_in),
    .io_reset(regs_246_io_reset),
    .io_out(regs_246_io_out),
    .io_enable(regs_246_io_enable)
  );
  FringeFF regs_247 ( // @[RegFile.scala 66:20:@45346.4]
    .clock(regs_247_clock),
    .reset(regs_247_reset),
    .io_in(regs_247_io_in),
    .io_reset(regs_247_io_reset),
    .io_out(regs_247_io_out),
    .io_enable(regs_247_io_enable)
  );
  FringeFF regs_248 ( // @[RegFile.scala 66:20:@45360.4]
    .clock(regs_248_clock),
    .reset(regs_248_reset),
    .io_in(regs_248_io_in),
    .io_reset(regs_248_io_reset),
    .io_out(regs_248_io_out),
    .io_enable(regs_248_io_enable)
  );
  FringeFF regs_249 ( // @[RegFile.scala 66:20:@45374.4]
    .clock(regs_249_clock),
    .reset(regs_249_reset),
    .io_in(regs_249_io_in),
    .io_reset(regs_249_io_reset),
    .io_out(regs_249_io_out),
    .io_enable(regs_249_io_enable)
  );
  FringeFF regs_250 ( // @[RegFile.scala 66:20:@45388.4]
    .clock(regs_250_clock),
    .reset(regs_250_reset),
    .io_in(regs_250_io_in),
    .io_reset(regs_250_io_reset),
    .io_out(regs_250_io_out),
    .io_enable(regs_250_io_enable)
  );
  FringeFF regs_251 ( // @[RegFile.scala 66:20:@45402.4]
    .clock(regs_251_clock),
    .reset(regs_251_reset),
    .io_in(regs_251_io_in),
    .io_reset(regs_251_io_reset),
    .io_out(regs_251_io_out),
    .io_enable(regs_251_io_enable)
  );
  FringeFF regs_252 ( // @[RegFile.scala 66:20:@45416.4]
    .clock(regs_252_clock),
    .reset(regs_252_reset),
    .io_in(regs_252_io_in),
    .io_reset(regs_252_io_reset),
    .io_out(regs_252_io_out),
    .io_enable(regs_252_io_enable)
  );
  FringeFF regs_253 ( // @[RegFile.scala 66:20:@45430.4]
    .clock(regs_253_clock),
    .reset(regs_253_reset),
    .io_in(regs_253_io_in),
    .io_reset(regs_253_io_reset),
    .io_out(regs_253_io_out),
    .io_enable(regs_253_io_enable)
  );
  FringeFF regs_254 ( // @[RegFile.scala 66:20:@45444.4]
    .clock(regs_254_clock),
    .reset(regs_254_reset),
    .io_in(regs_254_io_in),
    .io_reset(regs_254_io_reset),
    .io_out(regs_254_io_out),
    .io_enable(regs_254_io_enable)
  );
  FringeFF regs_255 ( // @[RegFile.scala 66:20:@45458.4]
    .clock(regs_255_clock),
    .reset(regs_255_reset),
    .io_in(regs_255_io_in),
    .io_reset(regs_255_io_reset),
    .io_out(regs_255_io_out),
    .io_enable(regs_255_io_enable)
  );
  FringeFF regs_256 ( // @[RegFile.scala 66:20:@45472.4]
    .clock(regs_256_clock),
    .reset(regs_256_reset),
    .io_in(regs_256_io_in),
    .io_reset(regs_256_io_reset),
    .io_out(regs_256_io_out),
    .io_enable(regs_256_io_enable)
  );
  FringeFF regs_257 ( // @[RegFile.scala 66:20:@45486.4]
    .clock(regs_257_clock),
    .reset(regs_257_reset),
    .io_in(regs_257_io_in),
    .io_reset(regs_257_io_reset),
    .io_out(regs_257_io_out),
    .io_enable(regs_257_io_enable)
  );
  FringeFF regs_258 ( // @[RegFile.scala 66:20:@45500.4]
    .clock(regs_258_clock),
    .reset(regs_258_reset),
    .io_in(regs_258_io_in),
    .io_reset(regs_258_io_reset),
    .io_out(regs_258_io_out),
    .io_enable(regs_258_io_enable)
  );
  FringeFF regs_259 ( // @[RegFile.scala 66:20:@45514.4]
    .clock(regs_259_clock),
    .reset(regs_259_reset),
    .io_in(regs_259_io_in),
    .io_reset(regs_259_io_reset),
    .io_out(regs_259_io_out),
    .io_enable(regs_259_io_enable)
  );
  FringeFF regs_260 ( // @[RegFile.scala 66:20:@45528.4]
    .clock(regs_260_clock),
    .reset(regs_260_reset),
    .io_in(regs_260_io_in),
    .io_reset(regs_260_io_reset),
    .io_out(regs_260_io_out),
    .io_enable(regs_260_io_enable)
  );
  FringeFF regs_261 ( // @[RegFile.scala 66:20:@45542.4]
    .clock(regs_261_clock),
    .reset(regs_261_reset),
    .io_in(regs_261_io_in),
    .io_reset(regs_261_io_reset),
    .io_out(regs_261_io_out),
    .io_enable(regs_261_io_enable)
  );
  FringeFF regs_262 ( // @[RegFile.scala 66:20:@45556.4]
    .clock(regs_262_clock),
    .reset(regs_262_reset),
    .io_in(regs_262_io_in),
    .io_reset(regs_262_io_reset),
    .io_out(regs_262_io_out),
    .io_enable(regs_262_io_enable)
  );
  FringeFF regs_263 ( // @[RegFile.scala 66:20:@45570.4]
    .clock(regs_263_clock),
    .reset(regs_263_reset),
    .io_in(regs_263_io_in),
    .io_reset(regs_263_io_reset),
    .io_out(regs_263_io_out),
    .io_enable(regs_263_io_enable)
  );
  FringeFF regs_264 ( // @[RegFile.scala 66:20:@45584.4]
    .clock(regs_264_clock),
    .reset(regs_264_reset),
    .io_in(regs_264_io_in),
    .io_reset(regs_264_io_reset),
    .io_out(regs_264_io_out),
    .io_enable(regs_264_io_enable)
  );
  FringeFF regs_265 ( // @[RegFile.scala 66:20:@45598.4]
    .clock(regs_265_clock),
    .reset(regs_265_reset),
    .io_in(regs_265_io_in),
    .io_reset(regs_265_io_reset),
    .io_out(regs_265_io_out),
    .io_enable(regs_265_io_enable)
  );
  FringeFF regs_266 ( // @[RegFile.scala 66:20:@45612.4]
    .clock(regs_266_clock),
    .reset(regs_266_reset),
    .io_in(regs_266_io_in),
    .io_reset(regs_266_io_reset),
    .io_out(regs_266_io_out),
    .io_enable(regs_266_io_enable)
  );
  FringeFF regs_267 ( // @[RegFile.scala 66:20:@45626.4]
    .clock(regs_267_clock),
    .reset(regs_267_reset),
    .io_in(regs_267_io_in),
    .io_reset(regs_267_io_reset),
    .io_out(regs_267_io_out),
    .io_enable(regs_267_io_enable)
  );
  FringeFF regs_268 ( // @[RegFile.scala 66:20:@45640.4]
    .clock(regs_268_clock),
    .reset(regs_268_reset),
    .io_in(regs_268_io_in),
    .io_reset(regs_268_io_reset),
    .io_out(regs_268_io_out),
    .io_enable(regs_268_io_enable)
  );
  FringeFF regs_269 ( // @[RegFile.scala 66:20:@45654.4]
    .clock(regs_269_clock),
    .reset(regs_269_reset),
    .io_in(regs_269_io_in),
    .io_reset(regs_269_io_reset),
    .io_out(regs_269_io_out),
    .io_enable(regs_269_io_enable)
  );
  FringeFF regs_270 ( // @[RegFile.scala 66:20:@45668.4]
    .clock(regs_270_clock),
    .reset(regs_270_reset),
    .io_in(regs_270_io_in),
    .io_reset(regs_270_io_reset),
    .io_out(regs_270_io_out),
    .io_enable(regs_270_io_enable)
  );
  FringeFF regs_271 ( // @[RegFile.scala 66:20:@45682.4]
    .clock(regs_271_clock),
    .reset(regs_271_reset),
    .io_in(regs_271_io_in),
    .io_reset(regs_271_io_reset),
    .io_out(regs_271_io_out),
    .io_enable(regs_271_io_enable)
  );
  FringeFF regs_272 ( // @[RegFile.scala 66:20:@45696.4]
    .clock(regs_272_clock),
    .reset(regs_272_reset),
    .io_in(regs_272_io_in),
    .io_reset(regs_272_io_reset),
    .io_out(regs_272_io_out),
    .io_enable(regs_272_io_enable)
  );
  FringeFF regs_273 ( // @[RegFile.scala 66:20:@45710.4]
    .clock(regs_273_clock),
    .reset(regs_273_reset),
    .io_in(regs_273_io_in),
    .io_reset(regs_273_io_reset),
    .io_out(regs_273_io_out),
    .io_enable(regs_273_io_enable)
  );
  FringeFF regs_274 ( // @[RegFile.scala 66:20:@45724.4]
    .clock(regs_274_clock),
    .reset(regs_274_reset),
    .io_in(regs_274_io_in),
    .io_reset(regs_274_io_reset),
    .io_out(regs_274_io_out),
    .io_enable(regs_274_io_enable)
  );
  FringeFF regs_275 ( // @[RegFile.scala 66:20:@45738.4]
    .clock(regs_275_clock),
    .reset(regs_275_reset),
    .io_in(regs_275_io_in),
    .io_reset(regs_275_io_reset),
    .io_out(regs_275_io_out),
    .io_enable(regs_275_io_enable)
  );
  FringeFF regs_276 ( // @[RegFile.scala 66:20:@45752.4]
    .clock(regs_276_clock),
    .reset(regs_276_reset),
    .io_in(regs_276_io_in),
    .io_reset(regs_276_io_reset),
    .io_out(regs_276_io_out),
    .io_enable(regs_276_io_enable)
  );
  FringeFF regs_277 ( // @[RegFile.scala 66:20:@45766.4]
    .clock(regs_277_clock),
    .reset(regs_277_reset),
    .io_in(regs_277_io_in),
    .io_reset(regs_277_io_reset),
    .io_out(regs_277_io_out),
    .io_enable(regs_277_io_enable)
  );
  FringeFF regs_278 ( // @[RegFile.scala 66:20:@45780.4]
    .clock(regs_278_clock),
    .reset(regs_278_reset),
    .io_in(regs_278_io_in),
    .io_reset(regs_278_io_reset),
    .io_out(regs_278_io_out),
    .io_enable(regs_278_io_enable)
  );
  FringeFF regs_279 ( // @[RegFile.scala 66:20:@45794.4]
    .clock(regs_279_clock),
    .reset(regs_279_reset),
    .io_in(regs_279_io_in),
    .io_reset(regs_279_io_reset),
    .io_out(regs_279_io_out),
    .io_enable(regs_279_io_enable)
  );
  FringeFF regs_280 ( // @[RegFile.scala 66:20:@45808.4]
    .clock(regs_280_clock),
    .reset(regs_280_reset),
    .io_in(regs_280_io_in),
    .io_reset(regs_280_io_reset),
    .io_out(regs_280_io_out),
    .io_enable(regs_280_io_enable)
  );
  FringeFF regs_281 ( // @[RegFile.scala 66:20:@45822.4]
    .clock(regs_281_clock),
    .reset(regs_281_reset),
    .io_in(regs_281_io_in),
    .io_reset(regs_281_io_reset),
    .io_out(regs_281_io_out),
    .io_enable(regs_281_io_enable)
  );
  FringeFF regs_282 ( // @[RegFile.scala 66:20:@45836.4]
    .clock(regs_282_clock),
    .reset(regs_282_reset),
    .io_in(regs_282_io_in),
    .io_reset(regs_282_io_reset),
    .io_out(regs_282_io_out),
    .io_enable(regs_282_io_enable)
  );
  FringeFF regs_283 ( // @[RegFile.scala 66:20:@45850.4]
    .clock(regs_283_clock),
    .reset(regs_283_reset),
    .io_in(regs_283_io_in),
    .io_reset(regs_283_io_reset),
    .io_out(regs_283_io_out),
    .io_enable(regs_283_io_enable)
  );
  FringeFF regs_284 ( // @[RegFile.scala 66:20:@45864.4]
    .clock(regs_284_clock),
    .reset(regs_284_reset),
    .io_in(regs_284_io_in),
    .io_reset(regs_284_io_reset),
    .io_out(regs_284_io_out),
    .io_enable(regs_284_io_enable)
  );
  FringeFF regs_285 ( // @[RegFile.scala 66:20:@45878.4]
    .clock(regs_285_clock),
    .reset(regs_285_reset),
    .io_in(regs_285_io_in),
    .io_reset(regs_285_io_reset),
    .io_out(regs_285_io_out),
    .io_enable(regs_285_io_enable)
  );
  FringeFF regs_286 ( // @[RegFile.scala 66:20:@45892.4]
    .clock(regs_286_clock),
    .reset(regs_286_reset),
    .io_in(regs_286_io_in),
    .io_reset(regs_286_io_reset),
    .io_out(regs_286_io_out),
    .io_enable(regs_286_io_enable)
  );
  FringeFF regs_287 ( // @[RegFile.scala 66:20:@45906.4]
    .clock(regs_287_clock),
    .reset(regs_287_reset),
    .io_in(regs_287_io_in),
    .io_reset(regs_287_io_reset),
    .io_out(regs_287_io_out),
    .io_enable(regs_287_io_enable)
  );
  FringeFF regs_288 ( // @[RegFile.scala 66:20:@45920.4]
    .clock(regs_288_clock),
    .reset(regs_288_reset),
    .io_in(regs_288_io_in),
    .io_reset(regs_288_io_reset),
    .io_out(regs_288_io_out),
    .io_enable(regs_288_io_enable)
  );
  FringeFF regs_289 ( // @[RegFile.scala 66:20:@45934.4]
    .clock(regs_289_clock),
    .reset(regs_289_reset),
    .io_in(regs_289_io_in),
    .io_reset(regs_289_io_reset),
    .io_out(regs_289_io_out),
    .io_enable(regs_289_io_enable)
  );
  FringeFF regs_290 ( // @[RegFile.scala 66:20:@45948.4]
    .clock(regs_290_clock),
    .reset(regs_290_reset),
    .io_in(regs_290_io_in),
    .io_reset(regs_290_io_reset),
    .io_out(regs_290_io_out),
    .io_enable(regs_290_io_enable)
  );
  FringeFF regs_291 ( // @[RegFile.scala 66:20:@45962.4]
    .clock(regs_291_clock),
    .reset(regs_291_reset),
    .io_in(regs_291_io_in),
    .io_reset(regs_291_io_reset),
    .io_out(regs_291_io_out),
    .io_enable(regs_291_io_enable)
  );
  FringeFF regs_292 ( // @[RegFile.scala 66:20:@45976.4]
    .clock(regs_292_clock),
    .reset(regs_292_reset),
    .io_in(regs_292_io_in),
    .io_reset(regs_292_io_reset),
    .io_out(regs_292_io_out),
    .io_enable(regs_292_io_enable)
  );
  FringeFF regs_293 ( // @[RegFile.scala 66:20:@45990.4]
    .clock(regs_293_clock),
    .reset(regs_293_reset),
    .io_in(regs_293_io_in),
    .io_reset(regs_293_io_reset),
    .io_out(regs_293_io_out),
    .io_enable(regs_293_io_enable)
  );
  FringeFF regs_294 ( // @[RegFile.scala 66:20:@46004.4]
    .clock(regs_294_clock),
    .reset(regs_294_reset),
    .io_in(regs_294_io_in),
    .io_reset(regs_294_io_reset),
    .io_out(regs_294_io_out),
    .io_enable(regs_294_io_enable)
  );
  FringeFF regs_295 ( // @[RegFile.scala 66:20:@46018.4]
    .clock(regs_295_clock),
    .reset(regs_295_reset),
    .io_in(regs_295_io_in),
    .io_reset(regs_295_io_reset),
    .io_out(regs_295_io_out),
    .io_enable(regs_295_io_enable)
  );
  FringeFF regs_296 ( // @[RegFile.scala 66:20:@46032.4]
    .clock(regs_296_clock),
    .reset(regs_296_reset),
    .io_in(regs_296_io_in),
    .io_reset(regs_296_io_reset),
    .io_out(regs_296_io_out),
    .io_enable(regs_296_io_enable)
  );
  FringeFF regs_297 ( // @[RegFile.scala 66:20:@46046.4]
    .clock(regs_297_clock),
    .reset(regs_297_reset),
    .io_in(regs_297_io_in),
    .io_reset(regs_297_io_reset),
    .io_out(regs_297_io_out),
    .io_enable(regs_297_io_enable)
  );
  FringeFF regs_298 ( // @[RegFile.scala 66:20:@46060.4]
    .clock(regs_298_clock),
    .reset(regs_298_reset),
    .io_in(regs_298_io_in),
    .io_reset(regs_298_io_reset),
    .io_out(regs_298_io_out),
    .io_enable(regs_298_io_enable)
  );
  FringeFF regs_299 ( // @[RegFile.scala 66:20:@46074.4]
    .clock(regs_299_clock),
    .reset(regs_299_reset),
    .io_in(regs_299_io_in),
    .io_reset(regs_299_io_reset),
    .io_out(regs_299_io_out),
    .io_enable(regs_299_io_enable)
  );
  FringeFF regs_300 ( // @[RegFile.scala 66:20:@46088.4]
    .clock(regs_300_clock),
    .reset(regs_300_reset),
    .io_in(regs_300_io_in),
    .io_reset(regs_300_io_reset),
    .io_out(regs_300_io_out),
    .io_enable(regs_300_io_enable)
  );
  FringeFF regs_301 ( // @[RegFile.scala 66:20:@46102.4]
    .clock(regs_301_clock),
    .reset(regs_301_reset),
    .io_in(regs_301_io_in),
    .io_reset(regs_301_io_reset),
    .io_out(regs_301_io_out),
    .io_enable(regs_301_io_enable)
  );
  FringeFF regs_302 ( // @[RegFile.scala 66:20:@46116.4]
    .clock(regs_302_clock),
    .reset(regs_302_reset),
    .io_in(regs_302_io_in),
    .io_reset(regs_302_io_reset),
    .io_out(regs_302_io_out),
    .io_enable(regs_302_io_enable)
  );
  FringeFF regs_303 ( // @[RegFile.scala 66:20:@46130.4]
    .clock(regs_303_clock),
    .reset(regs_303_reset),
    .io_in(regs_303_io_in),
    .io_reset(regs_303_io_reset),
    .io_out(regs_303_io_out),
    .io_enable(regs_303_io_enable)
  );
  FringeFF regs_304 ( // @[RegFile.scala 66:20:@46144.4]
    .clock(regs_304_clock),
    .reset(regs_304_reset),
    .io_in(regs_304_io_in),
    .io_reset(regs_304_io_reset),
    .io_out(regs_304_io_out),
    .io_enable(regs_304_io_enable)
  );
  FringeFF regs_305 ( // @[RegFile.scala 66:20:@46158.4]
    .clock(regs_305_clock),
    .reset(regs_305_reset),
    .io_in(regs_305_io_in),
    .io_reset(regs_305_io_reset),
    .io_out(regs_305_io_out),
    .io_enable(regs_305_io_enable)
  );
  FringeFF regs_306 ( // @[RegFile.scala 66:20:@46172.4]
    .clock(regs_306_clock),
    .reset(regs_306_reset),
    .io_in(regs_306_io_in),
    .io_reset(regs_306_io_reset),
    .io_out(regs_306_io_out),
    .io_enable(regs_306_io_enable)
  );
  FringeFF regs_307 ( // @[RegFile.scala 66:20:@46186.4]
    .clock(regs_307_clock),
    .reset(regs_307_reset),
    .io_in(regs_307_io_in),
    .io_reset(regs_307_io_reset),
    .io_out(regs_307_io_out),
    .io_enable(regs_307_io_enable)
  );
  FringeFF regs_308 ( // @[RegFile.scala 66:20:@46200.4]
    .clock(regs_308_clock),
    .reset(regs_308_reset),
    .io_in(regs_308_io_in),
    .io_reset(regs_308_io_reset),
    .io_out(regs_308_io_out),
    .io_enable(regs_308_io_enable)
  );
  FringeFF regs_309 ( // @[RegFile.scala 66:20:@46214.4]
    .clock(regs_309_clock),
    .reset(regs_309_reset),
    .io_in(regs_309_io_in),
    .io_reset(regs_309_io_reset),
    .io_out(regs_309_io_out),
    .io_enable(regs_309_io_enable)
  );
  FringeFF regs_310 ( // @[RegFile.scala 66:20:@46228.4]
    .clock(regs_310_clock),
    .reset(regs_310_reset),
    .io_in(regs_310_io_in),
    .io_reset(regs_310_io_reset),
    .io_out(regs_310_io_out),
    .io_enable(regs_310_io_enable)
  );
  FringeFF regs_311 ( // @[RegFile.scala 66:20:@46242.4]
    .clock(regs_311_clock),
    .reset(regs_311_reset),
    .io_in(regs_311_io_in),
    .io_reset(regs_311_io_reset),
    .io_out(regs_311_io_out),
    .io_enable(regs_311_io_enable)
  );
  FringeFF regs_312 ( // @[RegFile.scala 66:20:@46256.4]
    .clock(regs_312_clock),
    .reset(regs_312_reset),
    .io_in(regs_312_io_in),
    .io_reset(regs_312_io_reset),
    .io_out(regs_312_io_out),
    .io_enable(regs_312_io_enable)
  );
  FringeFF regs_313 ( // @[RegFile.scala 66:20:@46270.4]
    .clock(regs_313_clock),
    .reset(regs_313_reset),
    .io_in(regs_313_io_in),
    .io_reset(regs_313_io_reset),
    .io_out(regs_313_io_out),
    .io_enable(regs_313_io_enable)
  );
  FringeFF regs_314 ( // @[RegFile.scala 66:20:@46284.4]
    .clock(regs_314_clock),
    .reset(regs_314_reset),
    .io_in(regs_314_io_in),
    .io_reset(regs_314_io_reset),
    .io_out(regs_314_io_out),
    .io_enable(regs_314_io_enable)
  );
  FringeFF regs_315 ( // @[RegFile.scala 66:20:@46298.4]
    .clock(regs_315_clock),
    .reset(regs_315_reset),
    .io_in(regs_315_io_in),
    .io_reset(regs_315_io_reset),
    .io_out(regs_315_io_out),
    .io_enable(regs_315_io_enable)
  );
  FringeFF regs_316 ( // @[RegFile.scala 66:20:@46312.4]
    .clock(regs_316_clock),
    .reset(regs_316_reset),
    .io_in(regs_316_io_in),
    .io_reset(regs_316_io_reset),
    .io_out(regs_316_io_out),
    .io_enable(regs_316_io_enable)
  );
  FringeFF regs_317 ( // @[RegFile.scala 66:20:@46326.4]
    .clock(regs_317_clock),
    .reset(regs_317_reset),
    .io_in(regs_317_io_in),
    .io_reset(regs_317_io_reset),
    .io_out(regs_317_io_out),
    .io_enable(regs_317_io_enable)
  );
  FringeFF regs_318 ( // @[RegFile.scala 66:20:@46340.4]
    .clock(regs_318_clock),
    .reset(regs_318_reset),
    .io_in(regs_318_io_in),
    .io_reset(regs_318_io_reset),
    .io_out(regs_318_io_out),
    .io_enable(regs_318_io_enable)
  );
  FringeFF regs_319 ( // @[RegFile.scala 66:20:@46354.4]
    .clock(regs_319_clock),
    .reset(regs_319_reset),
    .io_in(regs_319_io_in),
    .io_reset(regs_319_io_reset),
    .io_out(regs_319_io_out),
    .io_enable(regs_319_io_enable)
  );
  FringeFF regs_320 ( // @[RegFile.scala 66:20:@46368.4]
    .clock(regs_320_clock),
    .reset(regs_320_reset),
    .io_in(regs_320_io_in),
    .io_reset(regs_320_io_reset),
    .io_out(regs_320_io_out),
    .io_enable(regs_320_io_enable)
  );
  FringeFF regs_321 ( // @[RegFile.scala 66:20:@46382.4]
    .clock(regs_321_clock),
    .reset(regs_321_reset),
    .io_in(regs_321_io_in),
    .io_reset(regs_321_io_reset),
    .io_out(regs_321_io_out),
    .io_enable(regs_321_io_enable)
  );
  FringeFF regs_322 ( // @[RegFile.scala 66:20:@46396.4]
    .clock(regs_322_clock),
    .reset(regs_322_reset),
    .io_in(regs_322_io_in),
    .io_reset(regs_322_io_reset),
    .io_out(regs_322_io_out),
    .io_enable(regs_322_io_enable)
  );
  FringeFF regs_323 ( // @[RegFile.scala 66:20:@46410.4]
    .clock(regs_323_clock),
    .reset(regs_323_reset),
    .io_in(regs_323_io_in),
    .io_reset(regs_323_io_reset),
    .io_out(regs_323_io_out),
    .io_enable(regs_323_io_enable)
  );
  FringeFF regs_324 ( // @[RegFile.scala 66:20:@46424.4]
    .clock(regs_324_clock),
    .reset(regs_324_reset),
    .io_in(regs_324_io_in),
    .io_reset(regs_324_io_reset),
    .io_out(regs_324_io_out),
    .io_enable(regs_324_io_enable)
  );
  FringeFF regs_325 ( // @[RegFile.scala 66:20:@46438.4]
    .clock(regs_325_clock),
    .reset(regs_325_reset),
    .io_in(regs_325_io_in),
    .io_reset(regs_325_io_reset),
    .io_out(regs_325_io_out),
    .io_enable(regs_325_io_enable)
  );
  FringeFF regs_326 ( // @[RegFile.scala 66:20:@46452.4]
    .clock(regs_326_clock),
    .reset(regs_326_reset),
    .io_in(regs_326_io_in),
    .io_reset(regs_326_io_reset),
    .io_out(regs_326_io_out),
    .io_enable(regs_326_io_enable)
  );
  FringeFF regs_327 ( // @[RegFile.scala 66:20:@46466.4]
    .clock(regs_327_clock),
    .reset(regs_327_reset),
    .io_in(regs_327_io_in),
    .io_reset(regs_327_io_reset),
    .io_out(regs_327_io_out),
    .io_enable(regs_327_io_enable)
  );
  FringeFF regs_328 ( // @[RegFile.scala 66:20:@46480.4]
    .clock(regs_328_clock),
    .reset(regs_328_reset),
    .io_in(regs_328_io_in),
    .io_reset(regs_328_io_reset),
    .io_out(regs_328_io_out),
    .io_enable(regs_328_io_enable)
  );
  FringeFF regs_329 ( // @[RegFile.scala 66:20:@46494.4]
    .clock(regs_329_clock),
    .reset(regs_329_reset),
    .io_in(regs_329_io_in),
    .io_reset(regs_329_io_reset),
    .io_out(regs_329_io_out),
    .io_enable(regs_329_io_enable)
  );
  FringeFF regs_330 ( // @[RegFile.scala 66:20:@46508.4]
    .clock(regs_330_clock),
    .reset(regs_330_reset),
    .io_in(regs_330_io_in),
    .io_reset(regs_330_io_reset),
    .io_out(regs_330_io_out),
    .io_enable(regs_330_io_enable)
  );
  FringeFF regs_331 ( // @[RegFile.scala 66:20:@46522.4]
    .clock(regs_331_clock),
    .reset(regs_331_reset),
    .io_in(regs_331_io_in),
    .io_reset(regs_331_io_reset),
    .io_out(regs_331_io_out),
    .io_enable(regs_331_io_enable)
  );
  FringeFF regs_332 ( // @[RegFile.scala 66:20:@46536.4]
    .clock(regs_332_clock),
    .reset(regs_332_reset),
    .io_in(regs_332_io_in),
    .io_reset(regs_332_io_reset),
    .io_out(regs_332_io_out),
    .io_enable(regs_332_io_enable)
  );
  FringeFF regs_333 ( // @[RegFile.scala 66:20:@46550.4]
    .clock(regs_333_clock),
    .reset(regs_333_reset),
    .io_in(regs_333_io_in),
    .io_reset(regs_333_io_reset),
    .io_out(regs_333_io_out),
    .io_enable(regs_333_io_enable)
  );
  FringeFF regs_334 ( // @[RegFile.scala 66:20:@46564.4]
    .clock(regs_334_clock),
    .reset(regs_334_reset),
    .io_in(regs_334_io_in),
    .io_reset(regs_334_io_reset),
    .io_out(regs_334_io_out),
    .io_enable(regs_334_io_enable)
  );
  FringeFF regs_335 ( // @[RegFile.scala 66:20:@46578.4]
    .clock(regs_335_clock),
    .reset(regs_335_reset),
    .io_in(regs_335_io_in),
    .io_reset(regs_335_io_reset),
    .io_out(regs_335_io_out),
    .io_enable(regs_335_io_enable)
  );
  FringeFF regs_336 ( // @[RegFile.scala 66:20:@46592.4]
    .clock(regs_336_clock),
    .reset(regs_336_reset),
    .io_in(regs_336_io_in),
    .io_reset(regs_336_io_reset),
    .io_out(regs_336_io_out),
    .io_enable(regs_336_io_enable)
  );
  FringeFF regs_337 ( // @[RegFile.scala 66:20:@46606.4]
    .clock(regs_337_clock),
    .reset(regs_337_reset),
    .io_in(regs_337_io_in),
    .io_reset(regs_337_io_reset),
    .io_out(regs_337_io_out),
    .io_enable(regs_337_io_enable)
  );
  FringeFF regs_338 ( // @[RegFile.scala 66:20:@46620.4]
    .clock(regs_338_clock),
    .reset(regs_338_reset),
    .io_in(regs_338_io_in),
    .io_reset(regs_338_io_reset),
    .io_out(regs_338_io_out),
    .io_enable(regs_338_io_enable)
  );
  FringeFF regs_339 ( // @[RegFile.scala 66:20:@46634.4]
    .clock(regs_339_clock),
    .reset(regs_339_reset),
    .io_in(regs_339_io_in),
    .io_reset(regs_339_io_reset),
    .io_out(regs_339_io_out),
    .io_enable(regs_339_io_enable)
  );
  FringeFF regs_340 ( // @[RegFile.scala 66:20:@46648.4]
    .clock(regs_340_clock),
    .reset(regs_340_reset),
    .io_in(regs_340_io_in),
    .io_reset(regs_340_io_reset),
    .io_out(regs_340_io_out),
    .io_enable(regs_340_io_enable)
  );
  FringeFF regs_341 ( // @[RegFile.scala 66:20:@46662.4]
    .clock(regs_341_clock),
    .reset(regs_341_reset),
    .io_in(regs_341_io_in),
    .io_reset(regs_341_io_reset),
    .io_out(regs_341_io_out),
    .io_enable(regs_341_io_enable)
  );
  FringeFF regs_342 ( // @[RegFile.scala 66:20:@46676.4]
    .clock(regs_342_clock),
    .reset(regs_342_reset),
    .io_in(regs_342_io_in),
    .io_reset(regs_342_io_reset),
    .io_out(regs_342_io_out),
    .io_enable(regs_342_io_enable)
  );
  FringeFF regs_343 ( // @[RegFile.scala 66:20:@46690.4]
    .clock(regs_343_clock),
    .reset(regs_343_reset),
    .io_in(regs_343_io_in),
    .io_reset(regs_343_io_reset),
    .io_out(regs_343_io_out),
    .io_enable(regs_343_io_enable)
  );
  FringeFF regs_344 ( // @[RegFile.scala 66:20:@46704.4]
    .clock(regs_344_clock),
    .reset(regs_344_reset),
    .io_in(regs_344_io_in),
    .io_reset(regs_344_io_reset),
    .io_out(regs_344_io_out),
    .io_enable(regs_344_io_enable)
  );
  FringeFF regs_345 ( // @[RegFile.scala 66:20:@46718.4]
    .clock(regs_345_clock),
    .reset(regs_345_reset),
    .io_in(regs_345_io_in),
    .io_reset(regs_345_io_reset),
    .io_out(regs_345_io_out),
    .io_enable(regs_345_io_enable)
  );
  FringeFF regs_346 ( // @[RegFile.scala 66:20:@46732.4]
    .clock(regs_346_clock),
    .reset(regs_346_reset),
    .io_in(regs_346_io_in),
    .io_reset(regs_346_io_reset),
    .io_out(regs_346_io_out),
    .io_enable(regs_346_io_enable)
  );
  FringeFF regs_347 ( // @[RegFile.scala 66:20:@46746.4]
    .clock(regs_347_clock),
    .reset(regs_347_reset),
    .io_in(regs_347_io_in),
    .io_reset(regs_347_io_reset),
    .io_out(regs_347_io_out),
    .io_enable(regs_347_io_enable)
  );
  FringeFF regs_348 ( // @[RegFile.scala 66:20:@46760.4]
    .clock(regs_348_clock),
    .reset(regs_348_reset),
    .io_in(regs_348_io_in),
    .io_reset(regs_348_io_reset),
    .io_out(regs_348_io_out),
    .io_enable(regs_348_io_enable)
  );
  FringeFF regs_349 ( // @[RegFile.scala 66:20:@46774.4]
    .clock(regs_349_clock),
    .reset(regs_349_reset),
    .io_in(regs_349_io_in),
    .io_reset(regs_349_io_reset),
    .io_out(regs_349_io_out),
    .io_enable(regs_349_io_enable)
  );
  FringeFF regs_350 ( // @[RegFile.scala 66:20:@46788.4]
    .clock(regs_350_clock),
    .reset(regs_350_reset),
    .io_in(regs_350_io_in),
    .io_reset(regs_350_io_reset),
    .io_out(regs_350_io_out),
    .io_enable(regs_350_io_enable)
  );
  FringeFF regs_351 ( // @[RegFile.scala 66:20:@46802.4]
    .clock(regs_351_clock),
    .reset(regs_351_reset),
    .io_in(regs_351_io_in),
    .io_reset(regs_351_io_reset),
    .io_out(regs_351_io_out),
    .io_enable(regs_351_io_enable)
  );
  FringeFF regs_352 ( // @[RegFile.scala 66:20:@46816.4]
    .clock(regs_352_clock),
    .reset(regs_352_reset),
    .io_in(regs_352_io_in),
    .io_reset(regs_352_io_reset),
    .io_out(regs_352_io_out),
    .io_enable(regs_352_io_enable)
  );
  FringeFF regs_353 ( // @[RegFile.scala 66:20:@46830.4]
    .clock(regs_353_clock),
    .reset(regs_353_reset),
    .io_in(regs_353_io_in),
    .io_reset(regs_353_io_reset),
    .io_out(regs_353_io_out),
    .io_enable(regs_353_io_enable)
  );
  FringeFF regs_354 ( // @[RegFile.scala 66:20:@46844.4]
    .clock(regs_354_clock),
    .reset(regs_354_reset),
    .io_in(regs_354_io_in),
    .io_reset(regs_354_io_reset),
    .io_out(regs_354_io_out),
    .io_enable(regs_354_io_enable)
  );
  FringeFF regs_355 ( // @[RegFile.scala 66:20:@46858.4]
    .clock(regs_355_clock),
    .reset(regs_355_reset),
    .io_in(regs_355_io_in),
    .io_reset(regs_355_io_reset),
    .io_out(regs_355_io_out),
    .io_enable(regs_355_io_enable)
  );
  FringeFF regs_356 ( // @[RegFile.scala 66:20:@46872.4]
    .clock(regs_356_clock),
    .reset(regs_356_reset),
    .io_in(regs_356_io_in),
    .io_reset(regs_356_io_reset),
    .io_out(regs_356_io_out),
    .io_enable(regs_356_io_enable)
  );
  FringeFF regs_357 ( // @[RegFile.scala 66:20:@46886.4]
    .clock(regs_357_clock),
    .reset(regs_357_reset),
    .io_in(regs_357_io_in),
    .io_reset(regs_357_io_reset),
    .io_out(regs_357_io_out),
    .io_enable(regs_357_io_enable)
  );
  FringeFF regs_358 ( // @[RegFile.scala 66:20:@46900.4]
    .clock(regs_358_clock),
    .reset(regs_358_reset),
    .io_in(regs_358_io_in),
    .io_reset(regs_358_io_reset),
    .io_out(regs_358_io_out),
    .io_enable(regs_358_io_enable)
  );
  FringeFF regs_359 ( // @[RegFile.scala 66:20:@46914.4]
    .clock(regs_359_clock),
    .reset(regs_359_reset),
    .io_in(regs_359_io_in),
    .io_reset(regs_359_io_reset),
    .io_out(regs_359_io_out),
    .io_enable(regs_359_io_enable)
  );
  FringeFF regs_360 ( // @[RegFile.scala 66:20:@46928.4]
    .clock(regs_360_clock),
    .reset(regs_360_reset),
    .io_in(regs_360_io_in),
    .io_reset(regs_360_io_reset),
    .io_out(regs_360_io_out),
    .io_enable(regs_360_io_enable)
  );
  FringeFF regs_361 ( // @[RegFile.scala 66:20:@46942.4]
    .clock(regs_361_clock),
    .reset(regs_361_reset),
    .io_in(regs_361_io_in),
    .io_reset(regs_361_io_reset),
    .io_out(regs_361_io_out),
    .io_enable(regs_361_io_enable)
  );
  FringeFF regs_362 ( // @[RegFile.scala 66:20:@46956.4]
    .clock(regs_362_clock),
    .reset(regs_362_reset),
    .io_in(regs_362_io_in),
    .io_reset(regs_362_io_reset),
    .io_out(regs_362_io_out),
    .io_enable(regs_362_io_enable)
  );
  FringeFF regs_363 ( // @[RegFile.scala 66:20:@46970.4]
    .clock(regs_363_clock),
    .reset(regs_363_reset),
    .io_in(regs_363_io_in),
    .io_reset(regs_363_io_reset),
    .io_out(regs_363_io_out),
    .io_enable(regs_363_io_enable)
  );
  FringeFF regs_364 ( // @[RegFile.scala 66:20:@46984.4]
    .clock(regs_364_clock),
    .reset(regs_364_reset),
    .io_in(regs_364_io_in),
    .io_reset(regs_364_io_reset),
    .io_out(regs_364_io_out),
    .io_enable(regs_364_io_enable)
  );
  FringeFF regs_365 ( // @[RegFile.scala 66:20:@46998.4]
    .clock(regs_365_clock),
    .reset(regs_365_reset),
    .io_in(regs_365_io_in),
    .io_reset(regs_365_io_reset),
    .io_out(regs_365_io_out),
    .io_enable(regs_365_io_enable)
  );
  FringeFF regs_366 ( // @[RegFile.scala 66:20:@47012.4]
    .clock(regs_366_clock),
    .reset(regs_366_reset),
    .io_in(regs_366_io_in),
    .io_reset(regs_366_io_reset),
    .io_out(regs_366_io_out),
    .io_enable(regs_366_io_enable)
  );
  FringeFF regs_367 ( // @[RegFile.scala 66:20:@47026.4]
    .clock(regs_367_clock),
    .reset(regs_367_reset),
    .io_in(regs_367_io_in),
    .io_reset(regs_367_io_reset),
    .io_out(regs_367_io_out),
    .io_enable(regs_367_io_enable)
  );
  FringeFF regs_368 ( // @[RegFile.scala 66:20:@47040.4]
    .clock(regs_368_clock),
    .reset(regs_368_reset),
    .io_in(regs_368_io_in),
    .io_reset(regs_368_io_reset),
    .io_out(regs_368_io_out),
    .io_enable(regs_368_io_enable)
  );
  FringeFF regs_369 ( // @[RegFile.scala 66:20:@47054.4]
    .clock(regs_369_clock),
    .reset(regs_369_reset),
    .io_in(regs_369_io_in),
    .io_reset(regs_369_io_reset),
    .io_out(regs_369_io_out),
    .io_enable(regs_369_io_enable)
  );
  FringeFF regs_370 ( // @[RegFile.scala 66:20:@47068.4]
    .clock(regs_370_clock),
    .reset(regs_370_reset),
    .io_in(regs_370_io_in),
    .io_reset(regs_370_io_reset),
    .io_out(regs_370_io_out),
    .io_enable(regs_370_io_enable)
  );
  FringeFF regs_371 ( // @[RegFile.scala 66:20:@47082.4]
    .clock(regs_371_clock),
    .reset(regs_371_reset),
    .io_in(regs_371_io_in),
    .io_reset(regs_371_io_reset),
    .io_out(regs_371_io_out),
    .io_enable(regs_371_io_enable)
  );
  FringeFF regs_372 ( // @[RegFile.scala 66:20:@47096.4]
    .clock(regs_372_clock),
    .reset(regs_372_reset),
    .io_in(regs_372_io_in),
    .io_reset(regs_372_io_reset),
    .io_out(regs_372_io_out),
    .io_enable(regs_372_io_enable)
  );
  FringeFF regs_373 ( // @[RegFile.scala 66:20:@47110.4]
    .clock(regs_373_clock),
    .reset(regs_373_reset),
    .io_in(regs_373_io_in),
    .io_reset(regs_373_io_reset),
    .io_out(regs_373_io_out),
    .io_enable(regs_373_io_enable)
  );
  FringeFF regs_374 ( // @[RegFile.scala 66:20:@47124.4]
    .clock(regs_374_clock),
    .reset(regs_374_reset),
    .io_in(regs_374_io_in),
    .io_reset(regs_374_io_reset),
    .io_out(regs_374_io_out),
    .io_enable(regs_374_io_enable)
  );
  FringeFF regs_375 ( // @[RegFile.scala 66:20:@47138.4]
    .clock(regs_375_clock),
    .reset(regs_375_reset),
    .io_in(regs_375_io_in),
    .io_reset(regs_375_io_reset),
    .io_out(regs_375_io_out),
    .io_enable(regs_375_io_enable)
  );
  FringeFF regs_376 ( // @[RegFile.scala 66:20:@47152.4]
    .clock(regs_376_clock),
    .reset(regs_376_reset),
    .io_in(regs_376_io_in),
    .io_reset(regs_376_io_reset),
    .io_out(regs_376_io_out),
    .io_enable(regs_376_io_enable)
  );
  FringeFF regs_377 ( // @[RegFile.scala 66:20:@47166.4]
    .clock(regs_377_clock),
    .reset(regs_377_reset),
    .io_in(regs_377_io_in),
    .io_reset(regs_377_io_reset),
    .io_out(regs_377_io_out),
    .io_enable(regs_377_io_enable)
  );
  FringeFF regs_378 ( // @[RegFile.scala 66:20:@47180.4]
    .clock(regs_378_clock),
    .reset(regs_378_reset),
    .io_in(regs_378_io_in),
    .io_reset(regs_378_io_reset),
    .io_out(regs_378_io_out),
    .io_enable(regs_378_io_enable)
  );
  FringeFF regs_379 ( // @[RegFile.scala 66:20:@47194.4]
    .clock(regs_379_clock),
    .reset(regs_379_reset),
    .io_in(regs_379_io_in),
    .io_reset(regs_379_io_reset),
    .io_out(regs_379_io_out),
    .io_enable(regs_379_io_enable)
  );
  FringeFF regs_380 ( // @[RegFile.scala 66:20:@47208.4]
    .clock(regs_380_clock),
    .reset(regs_380_reset),
    .io_in(regs_380_io_in),
    .io_reset(regs_380_io_reset),
    .io_out(regs_380_io_out),
    .io_enable(regs_380_io_enable)
  );
  FringeFF regs_381 ( // @[RegFile.scala 66:20:@47222.4]
    .clock(regs_381_clock),
    .reset(regs_381_reset),
    .io_in(regs_381_io_in),
    .io_reset(regs_381_io_reset),
    .io_out(regs_381_io_out),
    .io_enable(regs_381_io_enable)
  );
  FringeFF regs_382 ( // @[RegFile.scala 66:20:@47236.4]
    .clock(regs_382_clock),
    .reset(regs_382_reset),
    .io_in(regs_382_io_in),
    .io_reset(regs_382_io_reset),
    .io_out(regs_382_io_out),
    .io_enable(regs_382_io_enable)
  );
  FringeFF regs_383 ( // @[RegFile.scala 66:20:@47250.4]
    .clock(regs_383_clock),
    .reset(regs_383_reset),
    .io_in(regs_383_io_in),
    .io_reset(regs_383_io_reset),
    .io_out(regs_383_io_out),
    .io_enable(regs_383_io_enable)
  );
  FringeFF regs_384 ( // @[RegFile.scala 66:20:@47264.4]
    .clock(regs_384_clock),
    .reset(regs_384_reset),
    .io_in(regs_384_io_in),
    .io_reset(regs_384_io_reset),
    .io_out(regs_384_io_out),
    .io_enable(regs_384_io_enable)
  );
  FringeFF regs_385 ( // @[RegFile.scala 66:20:@47278.4]
    .clock(regs_385_clock),
    .reset(regs_385_reset),
    .io_in(regs_385_io_in),
    .io_reset(regs_385_io_reset),
    .io_out(regs_385_io_out),
    .io_enable(regs_385_io_enable)
  );
  FringeFF regs_386 ( // @[RegFile.scala 66:20:@47292.4]
    .clock(regs_386_clock),
    .reset(regs_386_reset),
    .io_in(regs_386_io_in),
    .io_reset(regs_386_io_reset),
    .io_out(regs_386_io_out),
    .io_enable(regs_386_io_enable)
  );
  FringeFF regs_387 ( // @[RegFile.scala 66:20:@47306.4]
    .clock(regs_387_clock),
    .reset(regs_387_reset),
    .io_in(regs_387_io_in),
    .io_reset(regs_387_io_reset),
    .io_out(regs_387_io_out),
    .io_enable(regs_387_io_enable)
  );
  FringeFF regs_388 ( // @[RegFile.scala 66:20:@47320.4]
    .clock(regs_388_clock),
    .reset(regs_388_reset),
    .io_in(regs_388_io_in),
    .io_reset(regs_388_io_reset),
    .io_out(regs_388_io_out),
    .io_enable(regs_388_io_enable)
  );
  FringeFF regs_389 ( // @[RegFile.scala 66:20:@47334.4]
    .clock(regs_389_clock),
    .reset(regs_389_reset),
    .io_in(regs_389_io_in),
    .io_reset(regs_389_io_reset),
    .io_out(regs_389_io_out),
    .io_enable(regs_389_io_enable)
  );
  FringeFF regs_390 ( // @[RegFile.scala 66:20:@47348.4]
    .clock(regs_390_clock),
    .reset(regs_390_reset),
    .io_in(regs_390_io_in),
    .io_reset(regs_390_io_reset),
    .io_out(regs_390_io_out),
    .io_enable(regs_390_io_enable)
  );
  FringeFF regs_391 ( // @[RegFile.scala 66:20:@47362.4]
    .clock(regs_391_clock),
    .reset(regs_391_reset),
    .io_in(regs_391_io_in),
    .io_reset(regs_391_io_reset),
    .io_out(regs_391_io_out),
    .io_enable(regs_391_io_enable)
  );
  FringeFF regs_392 ( // @[RegFile.scala 66:20:@47376.4]
    .clock(regs_392_clock),
    .reset(regs_392_reset),
    .io_in(regs_392_io_in),
    .io_reset(regs_392_io_reset),
    .io_out(regs_392_io_out),
    .io_enable(regs_392_io_enable)
  );
  FringeFF regs_393 ( // @[RegFile.scala 66:20:@47390.4]
    .clock(regs_393_clock),
    .reset(regs_393_reset),
    .io_in(regs_393_io_in),
    .io_reset(regs_393_io_reset),
    .io_out(regs_393_io_out),
    .io_enable(regs_393_io_enable)
  );
  FringeFF regs_394 ( // @[RegFile.scala 66:20:@47404.4]
    .clock(regs_394_clock),
    .reset(regs_394_reset),
    .io_in(regs_394_io_in),
    .io_reset(regs_394_io_reset),
    .io_out(regs_394_io_out),
    .io_enable(regs_394_io_enable)
  );
  FringeFF regs_395 ( // @[RegFile.scala 66:20:@47418.4]
    .clock(regs_395_clock),
    .reset(regs_395_reset),
    .io_in(regs_395_io_in),
    .io_reset(regs_395_io_reset),
    .io_out(regs_395_io_out),
    .io_enable(regs_395_io_enable)
  );
  FringeFF regs_396 ( // @[RegFile.scala 66:20:@47432.4]
    .clock(regs_396_clock),
    .reset(regs_396_reset),
    .io_in(regs_396_io_in),
    .io_reset(regs_396_io_reset),
    .io_out(regs_396_io_out),
    .io_enable(regs_396_io_enable)
  );
  FringeFF regs_397 ( // @[RegFile.scala 66:20:@47446.4]
    .clock(regs_397_clock),
    .reset(regs_397_reset),
    .io_in(regs_397_io_in),
    .io_reset(regs_397_io_reset),
    .io_out(regs_397_io_out),
    .io_enable(regs_397_io_enable)
  );
  FringeFF regs_398 ( // @[RegFile.scala 66:20:@47460.4]
    .clock(regs_398_clock),
    .reset(regs_398_reset),
    .io_in(regs_398_io_in),
    .io_reset(regs_398_io_reset),
    .io_out(regs_398_io_out),
    .io_enable(regs_398_io_enable)
  );
  FringeFF regs_399 ( // @[RegFile.scala 66:20:@47474.4]
    .clock(regs_399_clock),
    .reset(regs_399_reset),
    .io_in(regs_399_io_in),
    .io_reset(regs_399_io_reset),
    .io_out(regs_399_io_out),
    .io_enable(regs_399_io_enable)
  );
  FringeFF regs_400 ( // @[RegFile.scala 66:20:@47488.4]
    .clock(regs_400_clock),
    .reset(regs_400_reset),
    .io_in(regs_400_io_in),
    .io_reset(regs_400_io_reset),
    .io_out(regs_400_io_out),
    .io_enable(regs_400_io_enable)
  );
  FringeFF regs_401 ( // @[RegFile.scala 66:20:@47502.4]
    .clock(regs_401_clock),
    .reset(regs_401_reset),
    .io_in(regs_401_io_in),
    .io_reset(regs_401_io_reset),
    .io_out(regs_401_io_out),
    .io_enable(regs_401_io_enable)
  );
  FringeFF regs_402 ( // @[RegFile.scala 66:20:@47516.4]
    .clock(regs_402_clock),
    .reset(regs_402_reset),
    .io_in(regs_402_io_in),
    .io_reset(regs_402_io_reset),
    .io_out(regs_402_io_out),
    .io_enable(regs_402_io_enable)
  );
  FringeFF regs_403 ( // @[RegFile.scala 66:20:@47530.4]
    .clock(regs_403_clock),
    .reset(regs_403_reset),
    .io_in(regs_403_io_in),
    .io_reset(regs_403_io_reset),
    .io_out(regs_403_io_out),
    .io_enable(regs_403_io_enable)
  );
  FringeFF regs_404 ( // @[RegFile.scala 66:20:@47544.4]
    .clock(regs_404_clock),
    .reset(regs_404_reset),
    .io_in(regs_404_io_in),
    .io_reset(regs_404_io_reset),
    .io_out(regs_404_io_out),
    .io_enable(regs_404_io_enable)
  );
  FringeFF regs_405 ( // @[RegFile.scala 66:20:@47558.4]
    .clock(regs_405_clock),
    .reset(regs_405_reset),
    .io_in(regs_405_io_in),
    .io_reset(regs_405_io_reset),
    .io_out(regs_405_io_out),
    .io_enable(regs_405_io_enable)
  );
  FringeFF regs_406 ( // @[RegFile.scala 66:20:@47572.4]
    .clock(regs_406_clock),
    .reset(regs_406_reset),
    .io_in(regs_406_io_in),
    .io_reset(regs_406_io_reset),
    .io_out(regs_406_io_out),
    .io_enable(regs_406_io_enable)
  );
  FringeFF regs_407 ( // @[RegFile.scala 66:20:@47586.4]
    .clock(regs_407_clock),
    .reset(regs_407_reset),
    .io_in(regs_407_io_in),
    .io_reset(regs_407_io_reset),
    .io_out(regs_407_io_out),
    .io_enable(regs_407_io_enable)
  );
  FringeFF regs_408 ( // @[RegFile.scala 66:20:@47600.4]
    .clock(regs_408_clock),
    .reset(regs_408_reset),
    .io_in(regs_408_io_in),
    .io_reset(regs_408_io_reset),
    .io_out(regs_408_io_out),
    .io_enable(regs_408_io_enable)
  );
  FringeFF regs_409 ( // @[RegFile.scala 66:20:@47614.4]
    .clock(regs_409_clock),
    .reset(regs_409_reset),
    .io_in(regs_409_io_in),
    .io_reset(regs_409_io_reset),
    .io_out(regs_409_io_out),
    .io_enable(regs_409_io_enable)
  );
  FringeFF regs_410 ( // @[RegFile.scala 66:20:@47628.4]
    .clock(regs_410_clock),
    .reset(regs_410_reset),
    .io_in(regs_410_io_in),
    .io_reset(regs_410_io_reset),
    .io_out(regs_410_io_out),
    .io_enable(regs_410_io_enable)
  );
  FringeFF regs_411 ( // @[RegFile.scala 66:20:@47642.4]
    .clock(regs_411_clock),
    .reset(regs_411_reset),
    .io_in(regs_411_io_in),
    .io_reset(regs_411_io_reset),
    .io_out(regs_411_io_out),
    .io_enable(regs_411_io_enable)
  );
  FringeFF regs_412 ( // @[RegFile.scala 66:20:@47656.4]
    .clock(regs_412_clock),
    .reset(regs_412_reset),
    .io_in(regs_412_io_in),
    .io_reset(regs_412_io_reset),
    .io_out(regs_412_io_out),
    .io_enable(regs_412_io_enable)
  );
  FringeFF regs_413 ( // @[RegFile.scala 66:20:@47670.4]
    .clock(regs_413_clock),
    .reset(regs_413_reset),
    .io_in(regs_413_io_in),
    .io_reset(regs_413_io_reset),
    .io_out(regs_413_io_out),
    .io_enable(regs_413_io_enable)
  );
  FringeFF regs_414 ( // @[RegFile.scala 66:20:@47684.4]
    .clock(regs_414_clock),
    .reset(regs_414_reset),
    .io_in(regs_414_io_in),
    .io_reset(regs_414_io_reset),
    .io_out(regs_414_io_out),
    .io_enable(regs_414_io_enable)
  );
  FringeFF regs_415 ( // @[RegFile.scala 66:20:@47698.4]
    .clock(regs_415_clock),
    .reset(regs_415_reset),
    .io_in(regs_415_io_in),
    .io_reset(regs_415_io_reset),
    .io_out(regs_415_io_out),
    .io_enable(regs_415_io_enable)
  );
  FringeFF regs_416 ( // @[RegFile.scala 66:20:@47712.4]
    .clock(regs_416_clock),
    .reset(regs_416_reset),
    .io_in(regs_416_io_in),
    .io_reset(regs_416_io_reset),
    .io_out(regs_416_io_out),
    .io_enable(regs_416_io_enable)
  );
  FringeFF regs_417 ( // @[RegFile.scala 66:20:@47726.4]
    .clock(regs_417_clock),
    .reset(regs_417_reset),
    .io_in(regs_417_io_in),
    .io_reset(regs_417_io_reset),
    .io_out(regs_417_io_out),
    .io_enable(regs_417_io_enable)
  );
  FringeFF regs_418 ( // @[RegFile.scala 66:20:@47740.4]
    .clock(regs_418_clock),
    .reset(regs_418_reset),
    .io_in(regs_418_io_in),
    .io_reset(regs_418_io_reset),
    .io_out(regs_418_io_out),
    .io_enable(regs_418_io_enable)
  );
  FringeFF regs_419 ( // @[RegFile.scala 66:20:@47754.4]
    .clock(regs_419_clock),
    .reset(regs_419_reset),
    .io_in(regs_419_io_in),
    .io_reset(regs_419_io_reset),
    .io_out(regs_419_io_out),
    .io_enable(regs_419_io_enable)
  );
  FringeFF regs_420 ( // @[RegFile.scala 66:20:@47768.4]
    .clock(regs_420_clock),
    .reset(regs_420_reset),
    .io_in(regs_420_io_in),
    .io_reset(regs_420_io_reset),
    .io_out(regs_420_io_out),
    .io_enable(regs_420_io_enable)
  );
  FringeFF regs_421 ( // @[RegFile.scala 66:20:@47782.4]
    .clock(regs_421_clock),
    .reset(regs_421_reset),
    .io_in(regs_421_io_in),
    .io_reset(regs_421_io_reset),
    .io_out(regs_421_io_out),
    .io_enable(regs_421_io_enable)
  );
  FringeFF regs_422 ( // @[RegFile.scala 66:20:@47796.4]
    .clock(regs_422_clock),
    .reset(regs_422_reset),
    .io_in(regs_422_io_in),
    .io_reset(regs_422_io_reset),
    .io_out(regs_422_io_out),
    .io_enable(regs_422_io_enable)
  );
  FringeFF regs_423 ( // @[RegFile.scala 66:20:@47810.4]
    .clock(regs_423_clock),
    .reset(regs_423_reset),
    .io_in(regs_423_io_in),
    .io_reset(regs_423_io_reset),
    .io_out(regs_423_io_out),
    .io_enable(regs_423_io_enable)
  );
  FringeFF regs_424 ( // @[RegFile.scala 66:20:@47824.4]
    .clock(regs_424_clock),
    .reset(regs_424_reset),
    .io_in(regs_424_io_in),
    .io_reset(regs_424_io_reset),
    .io_out(regs_424_io_out),
    .io_enable(regs_424_io_enable)
  );
  FringeFF regs_425 ( // @[RegFile.scala 66:20:@47838.4]
    .clock(regs_425_clock),
    .reset(regs_425_reset),
    .io_in(regs_425_io_in),
    .io_reset(regs_425_io_reset),
    .io_out(regs_425_io_out),
    .io_enable(regs_425_io_enable)
  );
  FringeFF regs_426 ( // @[RegFile.scala 66:20:@47852.4]
    .clock(regs_426_clock),
    .reset(regs_426_reset),
    .io_in(regs_426_io_in),
    .io_reset(regs_426_io_reset),
    .io_out(regs_426_io_out),
    .io_enable(regs_426_io_enable)
  );
  FringeFF regs_427 ( // @[RegFile.scala 66:20:@47866.4]
    .clock(regs_427_clock),
    .reset(regs_427_reset),
    .io_in(regs_427_io_in),
    .io_reset(regs_427_io_reset),
    .io_out(regs_427_io_out),
    .io_enable(regs_427_io_enable)
  );
  FringeFF regs_428 ( // @[RegFile.scala 66:20:@47880.4]
    .clock(regs_428_clock),
    .reset(regs_428_reset),
    .io_in(regs_428_io_in),
    .io_reset(regs_428_io_reset),
    .io_out(regs_428_io_out),
    .io_enable(regs_428_io_enable)
  );
  FringeFF regs_429 ( // @[RegFile.scala 66:20:@47894.4]
    .clock(regs_429_clock),
    .reset(regs_429_reset),
    .io_in(regs_429_io_in),
    .io_reset(regs_429_io_reset),
    .io_out(regs_429_io_out),
    .io_enable(regs_429_io_enable)
  );
  FringeFF regs_430 ( // @[RegFile.scala 66:20:@47908.4]
    .clock(regs_430_clock),
    .reset(regs_430_reset),
    .io_in(regs_430_io_in),
    .io_reset(regs_430_io_reset),
    .io_out(regs_430_io_out),
    .io_enable(regs_430_io_enable)
  );
  FringeFF regs_431 ( // @[RegFile.scala 66:20:@47922.4]
    .clock(regs_431_clock),
    .reset(regs_431_reset),
    .io_in(regs_431_io_in),
    .io_reset(regs_431_io_reset),
    .io_out(regs_431_io_out),
    .io_enable(regs_431_io_enable)
  );
  FringeFF regs_432 ( // @[RegFile.scala 66:20:@47936.4]
    .clock(regs_432_clock),
    .reset(regs_432_reset),
    .io_in(regs_432_io_in),
    .io_reset(regs_432_io_reset),
    .io_out(regs_432_io_out),
    .io_enable(regs_432_io_enable)
  );
  FringeFF regs_433 ( // @[RegFile.scala 66:20:@47950.4]
    .clock(regs_433_clock),
    .reset(regs_433_reset),
    .io_in(regs_433_io_in),
    .io_reset(regs_433_io_reset),
    .io_out(regs_433_io_out),
    .io_enable(regs_433_io_enable)
  );
  FringeFF regs_434 ( // @[RegFile.scala 66:20:@47964.4]
    .clock(regs_434_clock),
    .reset(regs_434_reset),
    .io_in(regs_434_io_in),
    .io_reset(regs_434_io_reset),
    .io_out(regs_434_io_out),
    .io_enable(regs_434_io_enable)
  );
  FringeFF regs_435 ( // @[RegFile.scala 66:20:@47978.4]
    .clock(regs_435_clock),
    .reset(regs_435_reset),
    .io_in(regs_435_io_in),
    .io_reset(regs_435_io_reset),
    .io_out(regs_435_io_out),
    .io_enable(regs_435_io_enable)
  );
  FringeFF regs_436 ( // @[RegFile.scala 66:20:@47992.4]
    .clock(regs_436_clock),
    .reset(regs_436_reset),
    .io_in(regs_436_io_in),
    .io_reset(regs_436_io_reset),
    .io_out(regs_436_io_out),
    .io_enable(regs_436_io_enable)
  );
  FringeFF regs_437 ( // @[RegFile.scala 66:20:@48006.4]
    .clock(regs_437_clock),
    .reset(regs_437_reset),
    .io_in(regs_437_io_in),
    .io_reset(regs_437_io_reset),
    .io_out(regs_437_io_out),
    .io_enable(regs_437_io_enable)
  );
  FringeFF regs_438 ( // @[RegFile.scala 66:20:@48020.4]
    .clock(regs_438_clock),
    .reset(regs_438_reset),
    .io_in(regs_438_io_in),
    .io_reset(regs_438_io_reset),
    .io_out(regs_438_io_out),
    .io_enable(regs_438_io_enable)
  );
  FringeFF regs_439 ( // @[RegFile.scala 66:20:@48034.4]
    .clock(regs_439_clock),
    .reset(regs_439_reset),
    .io_in(regs_439_io_in),
    .io_reset(regs_439_io_reset),
    .io_out(regs_439_io_out),
    .io_enable(regs_439_io_enable)
  );
  FringeFF regs_440 ( // @[RegFile.scala 66:20:@48048.4]
    .clock(regs_440_clock),
    .reset(regs_440_reset),
    .io_in(regs_440_io_in),
    .io_reset(regs_440_io_reset),
    .io_out(regs_440_io_out),
    .io_enable(regs_440_io_enable)
  );
  FringeFF regs_441 ( // @[RegFile.scala 66:20:@48062.4]
    .clock(regs_441_clock),
    .reset(regs_441_reset),
    .io_in(regs_441_io_in),
    .io_reset(regs_441_io_reset),
    .io_out(regs_441_io_out),
    .io_enable(regs_441_io_enable)
  );
  FringeFF regs_442 ( // @[RegFile.scala 66:20:@48076.4]
    .clock(regs_442_clock),
    .reset(regs_442_reset),
    .io_in(regs_442_io_in),
    .io_reset(regs_442_io_reset),
    .io_out(regs_442_io_out),
    .io_enable(regs_442_io_enable)
  );
  FringeFF regs_443 ( // @[RegFile.scala 66:20:@48090.4]
    .clock(regs_443_clock),
    .reset(regs_443_reset),
    .io_in(regs_443_io_in),
    .io_reset(regs_443_io_reset),
    .io_out(regs_443_io_out),
    .io_enable(regs_443_io_enable)
  );
  FringeFF regs_444 ( // @[RegFile.scala 66:20:@48104.4]
    .clock(regs_444_clock),
    .reset(regs_444_reset),
    .io_in(regs_444_io_in),
    .io_reset(regs_444_io_reset),
    .io_out(regs_444_io_out),
    .io_enable(regs_444_io_enable)
  );
  FringeFF regs_445 ( // @[RegFile.scala 66:20:@48118.4]
    .clock(regs_445_clock),
    .reset(regs_445_reset),
    .io_in(regs_445_io_in),
    .io_reset(regs_445_io_reset),
    .io_out(regs_445_io_out),
    .io_enable(regs_445_io_enable)
  );
  FringeFF regs_446 ( // @[RegFile.scala 66:20:@48132.4]
    .clock(regs_446_clock),
    .reset(regs_446_reset),
    .io_in(regs_446_io_in),
    .io_reset(regs_446_io_reset),
    .io_out(regs_446_io_out),
    .io_enable(regs_446_io_enable)
  );
  FringeFF regs_447 ( // @[RegFile.scala 66:20:@48146.4]
    .clock(regs_447_clock),
    .reset(regs_447_reset),
    .io_in(regs_447_io_in),
    .io_reset(regs_447_io_reset),
    .io_out(regs_447_io_out),
    .io_enable(regs_447_io_enable)
  );
  FringeFF regs_448 ( // @[RegFile.scala 66:20:@48160.4]
    .clock(regs_448_clock),
    .reset(regs_448_reset),
    .io_in(regs_448_io_in),
    .io_reset(regs_448_io_reset),
    .io_out(regs_448_io_out),
    .io_enable(regs_448_io_enable)
  );
  FringeFF regs_449 ( // @[RegFile.scala 66:20:@48174.4]
    .clock(regs_449_clock),
    .reset(regs_449_reset),
    .io_in(regs_449_io_in),
    .io_reset(regs_449_io_reset),
    .io_out(regs_449_io_out),
    .io_enable(regs_449_io_enable)
  );
  FringeFF regs_450 ( // @[RegFile.scala 66:20:@48188.4]
    .clock(regs_450_clock),
    .reset(regs_450_reset),
    .io_in(regs_450_io_in),
    .io_reset(regs_450_io_reset),
    .io_out(regs_450_io_out),
    .io_enable(regs_450_io_enable)
  );
  FringeFF regs_451 ( // @[RegFile.scala 66:20:@48202.4]
    .clock(regs_451_clock),
    .reset(regs_451_reset),
    .io_in(regs_451_io_in),
    .io_reset(regs_451_io_reset),
    .io_out(regs_451_io_out),
    .io_enable(regs_451_io_enable)
  );
  FringeFF regs_452 ( // @[RegFile.scala 66:20:@48216.4]
    .clock(regs_452_clock),
    .reset(regs_452_reset),
    .io_in(regs_452_io_in),
    .io_reset(regs_452_io_reset),
    .io_out(regs_452_io_out),
    .io_enable(regs_452_io_enable)
  );
  FringeFF regs_453 ( // @[RegFile.scala 66:20:@48230.4]
    .clock(regs_453_clock),
    .reset(regs_453_reset),
    .io_in(regs_453_io_in),
    .io_reset(regs_453_io_reset),
    .io_out(regs_453_io_out),
    .io_enable(regs_453_io_enable)
  );
  FringeFF regs_454 ( // @[RegFile.scala 66:20:@48244.4]
    .clock(regs_454_clock),
    .reset(regs_454_reset),
    .io_in(regs_454_io_in),
    .io_reset(regs_454_io_reset),
    .io_out(regs_454_io_out),
    .io_enable(regs_454_io_enable)
  );
  FringeFF regs_455 ( // @[RegFile.scala 66:20:@48258.4]
    .clock(regs_455_clock),
    .reset(regs_455_reset),
    .io_in(regs_455_io_in),
    .io_reset(regs_455_io_reset),
    .io_out(regs_455_io_out),
    .io_enable(regs_455_io_enable)
  );
  FringeFF regs_456 ( // @[RegFile.scala 66:20:@48272.4]
    .clock(regs_456_clock),
    .reset(regs_456_reset),
    .io_in(regs_456_io_in),
    .io_reset(regs_456_io_reset),
    .io_out(regs_456_io_out),
    .io_enable(regs_456_io_enable)
  );
  FringeFF regs_457 ( // @[RegFile.scala 66:20:@48286.4]
    .clock(regs_457_clock),
    .reset(regs_457_reset),
    .io_in(regs_457_io_in),
    .io_reset(regs_457_io_reset),
    .io_out(regs_457_io_out),
    .io_enable(regs_457_io_enable)
  );
  FringeFF regs_458 ( // @[RegFile.scala 66:20:@48300.4]
    .clock(regs_458_clock),
    .reset(regs_458_reset),
    .io_in(regs_458_io_in),
    .io_reset(regs_458_io_reset),
    .io_out(regs_458_io_out),
    .io_enable(regs_458_io_enable)
  );
  FringeFF regs_459 ( // @[RegFile.scala 66:20:@48314.4]
    .clock(regs_459_clock),
    .reset(regs_459_reset),
    .io_in(regs_459_io_in),
    .io_reset(regs_459_io_reset),
    .io_out(regs_459_io_out),
    .io_enable(regs_459_io_enable)
  );
  FringeFF regs_460 ( // @[RegFile.scala 66:20:@48328.4]
    .clock(regs_460_clock),
    .reset(regs_460_reset),
    .io_in(regs_460_io_in),
    .io_reset(regs_460_io_reset),
    .io_out(regs_460_io_out),
    .io_enable(regs_460_io_enable)
  );
  FringeFF regs_461 ( // @[RegFile.scala 66:20:@48342.4]
    .clock(regs_461_clock),
    .reset(regs_461_reset),
    .io_in(regs_461_io_in),
    .io_reset(regs_461_io_reset),
    .io_out(regs_461_io_out),
    .io_enable(regs_461_io_enable)
  );
  FringeFF regs_462 ( // @[RegFile.scala 66:20:@48356.4]
    .clock(regs_462_clock),
    .reset(regs_462_reset),
    .io_in(regs_462_io_in),
    .io_reset(regs_462_io_reset),
    .io_out(regs_462_io_out),
    .io_enable(regs_462_io_enable)
  );
  FringeFF regs_463 ( // @[RegFile.scala 66:20:@48370.4]
    .clock(regs_463_clock),
    .reset(regs_463_reset),
    .io_in(regs_463_io_in),
    .io_reset(regs_463_io_reset),
    .io_out(regs_463_io_out),
    .io_enable(regs_463_io_enable)
  );
  FringeFF regs_464 ( // @[RegFile.scala 66:20:@48384.4]
    .clock(regs_464_clock),
    .reset(regs_464_reset),
    .io_in(regs_464_io_in),
    .io_reset(regs_464_io_reset),
    .io_out(regs_464_io_out),
    .io_enable(regs_464_io_enable)
  );
  FringeFF regs_465 ( // @[RegFile.scala 66:20:@48398.4]
    .clock(regs_465_clock),
    .reset(regs_465_reset),
    .io_in(regs_465_io_in),
    .io_reset(regs_465_io_reset),
    .io_out(regs_465_io_out),
    .io_enable(regs_465_io_enable)
  );
  FringeFF regs_466 ( // @[RegFile.scala 66:20:@48412.4]
    .clock(regs_466_clock),
    .reset(regs_466_reset),
    .io_in(regs_466_io_in),
    .io_reset(regs_466_io_reset),
    .io_out(regs_466_io_out),
    .io_enable(regs_466_io_enable)
  );
  FringeFF regs_467 ( // @[RegFile.scala 66:20:@48426.4]
    .clock(regs_467_clock),
    .reset(regs_467_reset),
    .io_in(regs_467_io_in),
    .io_reset(regs_467_io_reset),
    .io_out(regs_467_io_out),
    .io_enable(regs_467_io_enable)
  );
  FringeFF regs_468 ( // @[RegFile.scala 66:20:@48440.4]
    .clock(regs_468_clock),
    .reset(regs_468_reset),
    .io_in(regs_468_io_in),
    .io_reset(regs_468_io_reset),
    .io_out(regs_468_io_out),
    .io_enable(regs_468_io_enable)
  );
  FringeFF regs_469 ( // @[RegFile.scala 66:20:@48454.4]
    .clock(regs_469_clock),
    .reset(regs_469_reset),
    .io_in(regs_469_io_in),
    .io_reset(regs_469_io_reset),
    .io_out(regs_469_io_out),
    .io_enable(regs_469_io_enable)
  );
  FringeFF regs_470 ( // @[RegFile.scala 66:20:@48468.4]
    .clock(regs_470_clock),
    .reset(regs_470_reset),
    .io_in(regs_470_io_in),
    .io_reset(regs_470_io_reset),
    .io_out(regs_470_io_out),
    .io_enable(regs_470_io_enable)
  );
  FringeFF regs_471 ( // @[RegFile.scala 66:20:@48482.4]
    .clock(regs_471_clock),
    .reset(regs_471_reset),
    .io_in(regs_471_io_in),
    .io_reset(regs_471_io_reset),
    .io_out(regs_471_io_out),
    .io_enable(regs_471_io_enable)
  );
  FringeFF regs_472 ( // @[RegFile.scala 66:20:@48496.4]
    .clock(regs_472_clock),
    .reset(regs_472_reset),
    .io_in(regs_472_io_in),
    .io_reset(regs_472_io_reset),
    .io_out(regs_472_io_out),
    .io_enable(regs_472_io_enable)
  );
  FringeFF regs_473 ( // @[RegFile.scala 66:20:@48510.4]
    .clock(regs_473_clock),
    .reset(regs_473_reset),
    .io_in(regs_473_io_in),
    .io_reset(regs_473_io_reset),
    .io_out(regs_473_io_out),
    .io_enable(regs_473_io_enable)
  );
  FringeFF regs_474 ( // @[RegFile.scala 66:20:@48524.4]
    .clock(regs_474_clock),
    .reset(regs_474_reset),
    .io_in(regs_474_io_in),
    .io_reset(regs_474_io_reset),
    .io_out(regs_474_io_out),
    .io_enable(regs_474_io_enable)
  );
  FringeFF regs_475 ( // @[RegFile.scala 66:20:@48538.4]
    .clock(regs_475_clock),
    .reset(regs_475_reset),
    .io_in(regs_475_io_in),
    .io_reset(regs_475_io_reset),
    .io_out(regs_475_io_out),
    .io_enable(regs_475_io_enable)
  );
  FringeFF regs_476 ( // @[RegFile.scala 66:20:@48552.4]
    .clock(regs_476_clock),
    .reset(regs_476_reset),
    .io_in(regs_476_io_in),
    .io_reset(regs_476_io_reset),
    .io_out(regs_476_io_out),
    .io_enable(regs_476_io_enable)
  );
  FringeFF regs_477 ( // @[RegFile.scala 66:20:@48566.4]
    .clock(regs_477_clock),
    .reset(regs_477_reset),
    .io_in(regs_477_io_in),
    .io_reset(regs_477_io_reset),
    .io_out(regs_477_io_out),
    .io_enable(regs_477_io_enable)
  );
  FringeFF regs_478 ( // @[RegFile.scala 66:20:@48580.4]
    .clock(regs_478_clock),
    .reset(regs_478_reset),
    .io_in(regs_478_io_in),
    .io_reset(regs_478_io_reset),
    .io_out(regs_478_io_out),
    .io_enable(regs_478_io_enable)
  );
  FringeFF regs_479 ( // @[RegFile.scala 66:20:@48594.4]
    .clock(regs_479_clock),
    .reset(regs_479_reset),
    .io_in(regs_479_io_in),
    .io_reset(regs_479_io_reset),
    .io_out(regs_479_io_out),
    .io_enable(regs_479_io_enable)
  );
  FringeFF regs_480 ( // @[RegFile.scala 66:20:@48608.4]
    .clock(regs_480_clock),
    .reset(regs_480_reset),
    .io_in(regs_480_io_in),
    .io_reset(regs_480_io_reset),
    .io_out(regs_480_io_out),
    .io_enable(regs_480_io_enable)
  );
  FringeFF regs_481 ( // @[RegFile.scala 66:20:@48622.4]
    .clock(regs_481_clock),
    .reset(regs_481_reset),
    .io_in(regs_481_io_in),
    .io_reset(regs_481_io_reset),
    .io_out(regs_481_io_out),
    .io_enable(regs_481_io_enable)
  );
  FringeFF regs_482 ( // @[RegFile.scala 66:20:@48636.4]
    .clock(regs_482_clock),
    .reset(regs_482_reset),
    .io_in(regs_482_io_in),
    .io_reset(regs_482_io_reset),
    .io_out(regs_482_io_out),
    .io_enable(regs_482_io_enable)
  );
  FringeFF regs_483 ( // @[RegFile.scala 66:20:@48650.4]
    .clock(regs_483_clock),
    .reset(regs_483_reset),
    .io_in(regs_483_io_in),
    .io_reset(regs_483_io_reset),
    .io_out(regs_483_io_out),
    .io_enable(regs_483_io_enable)
  );
  FringeFF regs_484 ( // @[RegFile.scala 66:20:@48664.4]
    .clock(regs_484_clock),
    .reset(regs_484_reset),
    .io_in(regs_484_io_in),
    .io_reset(regs_484_io_reset),
    .io_out(regs_484_io_out),
    .io_enable(regs_484_io_enable)
  );
  FringeFF regs_485 ( // @[RegFile.scala 66:20:@48678.4]
    .clock(regs_485_clock),
    .reset(regs_485_reset),
    .io_in(regs_485_io_in),
    .io_reset(regs_485_io_reset),
    .io_out(regs_485_io_out),
    .io_enable(regs_485_io_enable)
  );
  FringeFF regs_486 ( // @[RegFile.scala 66:20:@48692.4]
    .clock(regs_486_clock),
    .reset(regs_486_reset),
    .io_in(regs_486_io_in),
    .io_reset(regs_486_io_reset),
    .io_out(regs_486_io_out),
    .io_enable(regs_486_io_enable)
  );
  FringeFF regs_487 ( // @[RegFile.scala 66:20:@48706.4]
    .clock(regs_487_clock),
    .reset(regs_487_reset),
    .io_in(regs_487_io_in),
    .io_reset(regs_487_io_reset),
    .io_out(regs_487_io_out),
    .io_enable(regs_487_io_enable)
  );
  FringeFF regs_488 ( // @[RegFile.scala 66:20:@48720.4]
    .clock(regs_488_clock),
    .reset(regs_488_reset),
    .io_in(regs_488_io_in),
    .io_reset(regs_488_io_reset),
    .io_out(regs_488_io_out),
    .io_enable(regs_488_io_enable)
  );
  FringeFF regs_489 ( // @[RegFile.scala 66:20:@48734.4]
    .clock(regs_489_clock),
    .reset(regs_489_reset),
    .io_in(regs_489_io_in),
    .io_reset(regs_489_io_reset),
    .io_out(regs_489_io_out),
    .io_enable(regs_489_io_enable)
  );
  FringeFF regs_490 ( // @[RegFile.scala 66:20:@48748.4]
    .clock(regs_490_clock),
    .reset(regs_490_reset),
    .io_in(regs_490_io_in),
    .io_reset(regs_490_io_reset),
    .io_out(regs_490_io_out),
    .io_enable(regs_490_io_enable)
  );
  FringeFF regs_491 ( // @[RegFile.scala 66:20:@48762.4]
    .clock(regs_491_clock),
    .reset(regs_491_reset),
    .io_in(regs_491_io_in),
    .io_reset(regs_491_io_reset),
    .io_out(regs_491_io_out),
    .io_enable(regs_491_io_enable)
  );
  FringeFF regs_492 ( // @[RegFile.scala 66:20:@48776.4]
    .clock(regs_492_clock),
    .reset(regs_492_reset),
    .io_in(regs_492_io_in),
    .io_reset(regs_492_io_reset),
    .io_out(regs_492_io_out),
    .io_enable(regs_492_io_enable)
  );
  FringeFF regs_493 ( // @[RegFile.scala 66:20:@48790.4]
    .clock(regs_493_clock),
    .reset(regs_493_reset),
    .io_in(regs_493_io_in),
    .io_reset(regs_493_io_reset),
    .io_out(regs_493_io_out),
    .io_enable(regs_493_io_enable)
  );
  FringeFF regs_494 ( // @[RegFile.scala 66:20:@48804.4]
    .clock(regs_494_clock),
    .reset(regs_494_reset),
    .io_in(regs_494_io_in),
    .io_reset(regs_494_io_reset),
    .io_out(regs_494_io_out),
    .io_enable(regs_494_io_enable)
  );
  FringeFF regs_495 ( // @[RegFile.scala 66:20:@48818.4]
    .clock(regs_495_clock),
    .reset(regs_495_reset),
    .io_in(regs_495_io_in),
    .io_reset(regs_495_io_reset),
    .io_out(regs_495_io_out),
    .io_enable(regs_495_io_enable)
  );
  FringeFF regs_496 ( // @[RegFile.scala 66:20:@48832.4]
    .clock(regs_496_clock),
    .reset(regs_496_reset),
    .io_in(regs_496_io_in),
    .io_reset(regs_496_io_reset),
    .io_out(regs_496_io_out),
    .io_enable(regs_496_io_enable)
  );
  FringeFF regs_497 ( // @[RegFile.scala 66:20:@48846.4]
    .clock(regs_497_clock),
    .reset(regs_497_reset),
    .io_in(regs_497_io_in),
    .io_reset(regs_497_io_reset),
    .io_out(regs_497_io_out),
    .io_enable(regs_497_io_enable)
  );
  FringeFF regs_498 ( // @[RegFile.scala 66:20:@48860.4]
    .clock(regs_498_clock),
    .reset(regs_498_reset),
    .io_in(regs_498_io_in),
    .io_reset(regs_498_io_reset),
    .io_out(regs_498_io_out),
    .io_enable(regs_498_io_enable)
  );
  FringeFF regs_499 ( // @[RegFile.scala 66:20:@48874.4]
    .clock(regs_499_clock),
    .reset(regs_499_reset),
    .io_in(regs_499_io_in),
    .io_reset(regs_499_io_reset),
    .io_out(regs_499_io_out),
    .io_enable(regs_499_io_enable)
  );
  FringeFF regs_500 ( // @[RegFile.scala 66:20:@48888.4]
    .clock(regs_500_clock),
    .reset(regs_500_reset),
    .io_in(regs_500_io_in),
    .io_reset(regs_500_io_reset),
    .io_out(regs_500_io_out),
    .io_enable(regs_500_io_enable)
  );
  FringeFF regs_501 ( // @[RegFile.scala 66:20:@48902.4]
    .clock(regs_501_clock),
    .reset(regs_501_reset),
    .io_in(regs_501_io_in),
    .io_reset(regs_501_io_reset),
    .io_out(regs_501_io_out),
    .io_enable(regs_501_io_enable)
  );
  FringeFF regs_502 ( // @[RegFile.scala 66:20:@48916.4]
    .clock(regs_502_clock),
    .reset(regs_502_reset),
    .io_in(regs_502_io_in),
    .io_reset(regs_502_io_reset),
    .io_out(regs_502_io_out),
    .io_enable(regs_502_io_enable)
  );
  FringeFF regs_503 ( // @[RegFile.scala 66:20:@48930.4]
    .clock(regs_503_clock),
    .reset(regs_503_reset),
    .io_in(regs_503_io_in),
    .io_reset(regs_503_io_reset),
    .io_out(regs_503_io_out),
    .io_enable(regs_503_io_enable)
  );
  FringeFF regs_504 ( // @[RegFile.scala 66:20:@48944.4]
    .clock(regs_504_clock),
    .reset(regs_504_reset),
    .io_in(regs_504_io_in),
    .io_reset(regs_504_io_reset),
    .io_out(regs_504_io_out),
    .io_enable(regs_504_io_enable)
  );
  FringeFF regs_505 ( // @[RegFile.scala 66:20:@48958.4]
    .clock(regs_505_clock),
    .reset(regs_505_reset),
    .io_in(regs_505_io_in),
    .io_reset(regs_505_io_reset),
    .io_out(regs_505_io_out),
    .io_enable(regs_505_io_enable)
  );
  FringeFF regs_506 ( // @[RegFile.scala 66:20:@48972.4]
    .clock(regs_506_clock),
    .reset(regs_506_reset),
    .io_in(regs_506_io_in),
    .io_reset(regs_506_io_reset),
    .io_out(regs_506_io_out),
    .io_enable(regs_506_io_enable)
  );
  FringeFF regs_507 ( // @[RegFile.scala 66:20:@48986.4]
    .clock(regs_507_clock),
    .reset(regs_507_reset),
    .io_in(regs_507_io_in),
    .io_reset(regs_507_io_reset),
    .io_out(regs_507_io_out),
    .io_enable(regs_507_io_enable)
  );
  FringeFF regs_508 ( // @[RegFile.scala 66:20:@49000.4]
    .clock(regs_508_clock),
    .reset(regs_508_reset),
    .io_in(regs_508_io_in),
    .io_reset(regs_508_io_reset),
    .io_out(regs_508_io_out),
    .io_enable(regs_508_io_enable)
  );
  FringeFF regs_509 ( // @[RegFile.scala 66:20:@49014.4]
    .clock(regs_509_clock),
    .reset(regs_509_reset),
    .io_in(regs_509_io_in),
    .io_reset(regs_509_io_reset),
    .io_out(regs_509_io_out),
    .io_enable(regs_509_io_enable)
  );
  FringeFF regs_510 ( // @[RegFile.scala 66:20:@49028.4]
    .clock(regs_510_clock),
    .reset(regs_510_reset),
    .io_in(regs_510_io_in),
    .io_reset(regs_510_io_reset),
    .io_out(regs_510_io_out),
    .io_enable(regs_510_io_enable)
  );
  FringeFF regs_511 ( // @[RegFile.scala 66:20:@49042.4]
    .clock(regs_511_clock),
    .reset(regs_511_reset),
    .io_in(regs_511_io_in),
    .io_reset(regs_511_io_reset),
    .io_out(regs_511_io_out),
    .io_enable(regs_511_io_enable)
  );
  FringeFF regs_512 ( // @[RegFile.scala 66:20:@49056.4]
    .clock(regs_512_clock),
    .reset(regs_512_reset),
    .io_in(regs_512_io_in),
    .io_reset(regs_512_io_reset),
    .io_out(regs_512_io_out),
    .io_enable(regs_512_io_enable)
  );
  FringeFF regs_513 ( // @[RegFile.scala 66:20:@49070.4]
    .clock(regs_513_clock),
    .reset(regs_513_reset),
    .io_in(regs_513_io_in),
    .io_reset(regs_513_io_reset),
    .io_out(regs_513_io_out),
    .io_enable(regs_513_io_enable)
  );
  FringeFF regs_514 ( // @[RegFile.scala 66:20:@49084.4]
    .clock(regs_514_clock),
    .reset(regs_514_reset),
    .io_in(regs_514_io_in),
    .io_reset(regs_514_io_reset),
    .io_out(regs_514_io_out),
    .io_enable(regs_514_io_enable)
  );
  FringeFF regs_515 ( // @[RegFile.scala 66:20:@49098.4]
    .clock(regs_515_clock),
    .reset(regs_515_reset),
    .io_in(regs_515_io_in),
    .io_reset(regs_515_io_reset),
    .io_out(regs_515_io_out),
    .io_enable(regs_515_io_enable)
  );
  FringeFF regs_516 ( // @[RegFile.scala 66:20:@49112.4]
    .clock(regs_516_clock),
    .reset(regs_516_reset),
    .io_in(regs_516_io_in),
    .io_reset(regs_516_io_reset),
    .io_out(regs_516_io_out),
    .io_enable(regs_516_io_enable)
  );
  FringeFF regs_517 ( // @[RegFile.scala 66:20:@49126.4]
    .clock(regs_517_clock),
    .reset(regs_517_reset),
    .io_in(regs_517_io_in),
    .io_reset(regs_517_io_reset),
    .io_out(regs_517_io_out),
    .io_enable(regs_517_io_enable)
  );
  FringeFF regs_518 ( // @[RegFile.scala 66:20:@49140.4]
    .clock(regs_518_clock),
    .reset(regs_518_reset),
    .io_in(regs_518_io_in),
    .io_reset(regs_518_io_reset),
    .io_out(regs_518_io_out),
    .io_enable(regs_518_io_enable)
  );
  FringeFF regs_519 ( // @[RegFile.scala 66:20:@49154.4]
    .clock(regs_519_clock),
    .reset(regs_519_reset),
    .io_in(regs_519_io_in),
    .io_reset(regs_519_io_reset),
    .io_out(regs_519_io_out),
    .io_enable(regs_519_io_enable)
  );
  FringeFF regs_520 ( // @[RegFile.scala 66:20:@49168.4]
    .clock(regs_520_clock),
    .reset(regs_520_reset),
    .io_in(regs_520_io_in),
    .io_reset(regs_520_io_reset),
    .io_out(regs_520_io_out),
    .io_enable(regs_520_io_enable)
  );
  FringeFF regs_521 ( // @[RegFile.scala 66:20:@49182.4]
    .clock(regs_521_clock),
    .reset(regs_521_reset),
    .io_in(regs_521_io_in),
    .io_reset(regs_521_io_reset),
    .io_out(regs_521_io_out),
    .io_enable(regs_521_io_enable)
  );
  MuxN rport ( // @[RegFile.scala 95:21:@49196.4]
    .io_ins_0(rport_io_ins_0),
    .io_ins_1(rport_io_ins_1),
    .io_ins_2(rport_io_ins_2),
    .io_ins_3(rport_io_ins_3),
    .io_ins_4(rport_io_ins_4),
    .io_ins_5(rport_io_ins_5),
    .io_ins_6(rport_io_ins_6),
    .io_ins_7(rport_io_ins_7),
    .io_ins_8(rport_io_ins_8),
    .io_ins_9(rport_io_ins_9),
    .io_ins_10(rport_io_ins_10),
    .io_ins_11(rport_io_ins_11),
    .io_ins_12(rport_io_ins_12),
    .io_ins_13(rport_io_ins_13),
    .io_ins_14(rport_io_ins_14),
    .io_ins_15(rport_io_ins_15),
    .io_ins_16(rport_io_ins_16),
    .io_ins_17(rport_io_ins_17),
    .io_ins_18(rport_io_ins_18),
    .io_ins_19(rport_io_ins_19),
    .io_ins_20(rport_io_ins_20),
    .io_ins_21(rport_io_ins_21),
    .io_ins_22(rport_io_ins_22),
    .io_ins_23(rport_io_ins_23),
    .io_ins_24(rport_io_ins_24),
    .io_ins_25(rport_io_ins_25),
    .io_ins_26(rport_io_ins_26),
    .io_ins_27(rport_io_ins_27),
    .io_ins_28(rport_io_ins_28),
    .io_ins_29(rport_io_ins_29),
    .io_ins_30(rport_io_ins_30),
    .io_ins_31(rport_io_ins_31),
    .io_ins_32(rport_io_ins_32),
    .io_ins_33(rport_io_ins_33),
    .io_ins_34(rport_io_ins_34),
    .io_ins_35(rport_io_ins_35),
    .io_ins_36(rport_io_ins_36),
    .io_ins_37(rport_io_ins_37),
    .io_ins_38(rport_io_ins_38),
    .io_ins_39(rport_io_ins_39),
    .io_ins_40(rport_io_ins_40),
    .io_ins_41(rport_io_ins_41),
    .io_ins_42(rport_io_ins_42),
    .io_ins_43(rport_io_ins_43),
    .io_ins_44(rport_io_ins_44),
    .io_ins_45(rport_io_ins_45),
    .io_ins_46(rport_io_ins_46),
    .io_ins_47(rport_io_ins_47),
    .io_ins_48(rport_io_ins_48),
    .io_ins_49(rport_io_ins_49),
    .io_ins_50(rport_io_ins_50),
    .io_ins_51(rport_io_ins_51),
    .io_ins_52(rport_io_ins_52),
    .io_ins_53(rport_io_ins_53),
    .io_ins_54(rport_io_ins_54),
    .io_ins_55(rport_io_ins_55),
    .io_ins_56(rport_io_ins_56),
    .io_ins_57(rport_io_ins_57),
    .io_ins_58(rport_io_ins_58),
    .io_ins_59(rport_io_ins_59),
    .io_ins_60(rport_io_ins_60),
    .io_ins_61(rport_io_ins_61),
    .io_ins_62(rport_io_ins_62),
    .io_ins_63(rport_io_ins_63),
    .io_ins_64(rport_io_ins_64),
    .io_ins_65(rport_io_ins_65),
    .io_ins_66(rport_io_ins_66),
    .io_ins_67(rport_io_ins_67),
    .io_ins_68(rport_io_ins_68),
    .io_ins_69(rport_io_ins_69),
    .io_ins_70(rport_io_ins_70),
    .io_ins_71(rport_io_ins_71),
    .io_ins_72(rport_io_ins_72),
    .io_ins_73(rport_io_ins_73),
    .io_ins_74(rport_io_ins_74),
    .io_ins_75(rport_io_ins_75),
    .io_ins_76(rport_io_ins_76),
    .io_ins_77(rport_io_ins_77),
    .io_ins_78(rport_io_ins_78),
    .io_ins_79(rport_io_ins_79),
    .io_ins_80(rport_io_ins_80),
    .io_ins_81(rport_io_ins_81),
    .io_ins_82(rport_io_ins_82),
    .io_ins_83(rport_io_ins_83),
    .io_ins_84(rport_io_ins_84),
    .io_ins_85(rport_io_ins_85),
    .io_ins_86(rport_io_ins_86),
    .io_ins_87(rport_io_ins_87),
    .io_ins_88(rport_io_ins_88),
    .io_ins_89(rport_io_ins_89),
    .io_ins_90(rport_io_ins_90),
    .io_ins_91(rport_io_ins_91),
    .io_ins_92(rport_io_ins_92),
    .io_ins_93(rport_io_ins_93),
    .io_ins_94(rport_io_ins_94),
    .io_ins_95(rport_io_ins_95),
    .io_ins_96(rport_io_ins_96),
    .io_ins_97(rport_io_ins_97),
    .io_ins_98(rport_io_ins_98),
    .io_ins_99(rport_io_ins_99),
    .io_ins_100(rport_io_ins_100),
    .io_ins_101(rport_io_ins_101),
    .io_ins_102(rport_io_ins_102),
    .io_ins_103(rport_io_ins_103),
    .io_ins_104(rport_io_ins_104),
    .io_ins_105(rport_io_ins_105),
    .io_ins_106(rport_io_ins_106),
    .io_ins_107(rport_io_ins_107),
    .io_ins_108(rport_io_ins_108),
    .io_ins_109(rport_io_ins_109),
    .io_ins_110(rport_io_ins_110),
    .io_ins_111(rport_io_ins_111),
    .io_ins_112(rport_io_ins_112),
    .io_ins_113(rport_io_ins_113),
    .io_ins_114(rport_io_ins_114),
    .io_ins_115(rport_io_ins_115),
    .io_ins_116(rport_io_ins_116),
    .io_ins_117(rport_io_ins_117),
    .io_ins_118(rport_io_ins_118),
    .io_ins_119(rport_io_ins_119),
    .io_ins_120(rport_io_ins_120),
    .io_ins_121(rport_io_ins_121),
    .io_ins_122(rport_io_ins_122),
    .io_ins_123(rport_io_ins_123),
    .io_ins_124(rport_io_ins_124),
    .io_ins_125(rport_io_ins_125),
    .io_ins_126(rport_io_ins_126),
    .io_ins_127(rport_io_ins_127),
    .io_ins_128(rport_io_ins_128),
    .io_ins_129(rport_io_ins_129),
    .io_ins_130(rport_io_ins_130),
    .io_ins_131(rport_io_ins_131),
    .io_ins_132(rport_io_ins_132),
    .io_ins_133(rport_io_ins_133),
    .io_ins_134(rport_io_ins_134),
    .io_ins_135(rport_io_ins_135),
    .io_ins_136(rport_io_ins_136),
    .io_ins_137(rport_io_ins_137),
    .io_ins_138(rport_io_ins_138),
    .io_ins_139(rport_io_ins_139),
    .io_ins_140(rport_io_ins_140),
    .io_ins_141(rport_io_ins_141),
    .io_ins_142(rport_io_ins_142),
    .io_ins_143(rport_io_ins_143),
    .io_ins_144(rport_io_ins_144),
    .io_ins_145(rport_io_ins_145),
    .io_ins_146(rport_io_ins_146),
    .io_ins_147(rport_io_ins_147),
    .io_ins_148(rport_io_ins_148),
    .io_ins_149(rport_io_ins_149),
    .io_ins_150(rport_io_ins_150),
    .io_ins_151(rport_io_ins_151),
    .io_ins_152(rport_io_ins_152),
    .io_ins_153(rport_io_ins_153),
    .io_ins_154(rport_io_ins_154),
    .io_ins_155(rport_io_ins_155),
    .io_ins_156(rport_io_ins_156),
    .io_ins_157(rport_io_ins_157),
    .io_ins_158(rport_io_ins_158),
    .io_ins_159(rport_io_ins_159),
    .io_ins_160(rport_io_ins_160),
    .io_ins_161(rport_io_ins_161),
    .io_ins_162(rport_io_ins_162),
    .io_ins_163(rport_io_ins_163),
    .io_ins_164(rport_io_ins_164),
    .io_ins_165(rport_io_ins_165),
    .io_ins_166(rport_io_ins_166),
    .io_ins_167(rport_io_ins_167),
    .io_ins_168(rport_io_ins_168),
    .io_ins_169(rport_io_ins_169),
    .io_ins_170(rport_io_ins_170),
    .io_ins_171(rport_io_ins_171),
    .io_ins_172(rport_io_ins_172),
    .io_ins_173(rport_io_ins_173),
    .io_ins_174(rport_io_ins_174),
    .io_ins_175(rport_io_ins_175),
    .io_ins_176(rport_io_ins_176),
    .io_ins_177(rport_io_ins_177),
    .io_ins_178(rport_io_ins_178),
    .io_ins_179(rport_io_ins_179),
    .io_ins_180(rport_io_ins_180),
    .io_ins_181(rport_io_ins_181),
    .io_ins_182(rport_io_ins_182),
    .io_ins_183(rport_io_ins_183),
    .io_ins_184(rport_io_ins_184),
    .io_ins_185(rport_io_ins_185),
    .io_ins_186(rport_io_ins_186),
    .io_ins_187(rport_io_ins_187),
    .io_ins_188(rport_io_ins_188),
    .io_ins_189(rport_io_ins_189),
    .io_ins_190(rport_io_ins_190),
    .io_ins_191(rport_io_ins_191),
    .io_ins_192(rport_io_ins_192),
    .io_ins_193(rport_io_ins_193),
    .io_ins_194(rport_io_ins_194),
    .io_ins_195(rport_io_ins_195),
    .io_ins_196(rport_io_ins_196),
    .io_ins_197(rport_io_ins_197),
    .io_ins_198(rport_io_ins_198),
    .io_ins_199(rport_io_ins_199),
    .io_ins_200(rport_io_ins_200),
    .io_ins_201(rport_io_ins_201),
    .io_ins_202(rport_io_ins_202),
    .io_ins_203(rport_io_ins_203),
    .io_ins_204(rport_io_ins_204),
    .io_ins_205(rport_io_ins_205),
    .io_ins_206(rport_io_ins_206),
    .io_ins_207(rport_io_ins_207),
    .io_ins_208(rport_io_ins_208),
    .io_ins_209(rport_io_ins_209),
    .io_ins_210(rport_io_ins_210),
    .io_ins_211(rport_io_ins_211),
    .io_ins_212(rport_io_ins_212),
    .io_ins_213(rport_io_ins_213),
    .io_ins_214(rport_io_ins_214),
    .io_ins_215(rport_io_ins_215),
    .io_ins_216(rport_io_ins_216),
    .io_ins_217(rport_io_ins_217),
    .io_ins_218(rport_io_ins_218),
    .io_ins_219(rport_io_ins_219),
    .io_ins_220(rport_io_ins_220),
    .io_ins_221(rport_io_ins_221),
    .io_ins_222(rport_io_ins_222),
    .io_ins_223(rport_io_ins_223),
    .io_ins_224(rport_io_ins_224),
    .io_ins_225(rport_io_ins_225),
    .io_ins_226(rport_io_ins_226),
    .io_ins_227(rport_io_ins_227),
    .io_ins_228(rport_io_ins_228),
    .io_ins_229(rport_io_ins_229),
    .io_ins_230(rport_io_ins_230),
    .io_ins_231(rport_io_ins_231),
    .io_ins_232(rport_io_ins_232),
    .io_ins_233(rport_io_ins_233),
    .io_ins_234(rport_io_ins_234),
    .io_ins_235(rport_io_ins_235),
    .io_ins_236(rport_io_ins_236),
    .io_ins_237(rport_io_ins_237),
    .io_ins_238(rport_io_ins_238),
    .io_ins_239(rport_io_ins_239),
    .io_ins_240(rport_io_ins_240),
    .io_ins_241(rport_io_ins_241),
    .io_ins_242(rport_io_ins_242),
    .io_ins_243(rport_io_ins_243),
    .io_ins_244(rport_io_ins_244),
    .io_ins_245(rport_io_ins_245),
    .io_ins_246(rport_io_ins_246),
    .io_ins_247(rport_io_ins_247),
    .io_ins_248(rport_io_ins_248),
    .io_ins_249(rport_io_ins_249),
    .io_ins_250(rport_io_ins_250),
    .io_ins_251(rport_io_ins_251),
    .io_ins_252(rport_io_ins_252),
    .io_ins_253(rport_io_ins_253),
    .io_ins_254(rport_io_ins_254),
    .io_ins_255(rport_io_ins_255),
    .io_ins_256(rport_io_ins_256),
    .io_ins_257(rport_io_ins_257),
    .io_ins_258(rport_io_ins_258),
    .io_ins_259(rport_io_ins_259),
    .io_ins_260(rport_io_ins_260),
    .io_ins_261(rport_io_ins_261),
    .io_ins_262(rport_io_ins_262),
    .io_ins_263(rport_io_ins_263),
    .io_ins_264(rport_io_ins_264),
    .io_ins_265(rport_io_ins_265),
    .io_ins_266(rport_io_ins_266),
    .io_ins_267(rport_io_ins_267),
    .io_ins_268(rport_io_ins_268),
    .io_ins_269(rport_io_ins_269),
    .io_ins_270(rport_io_ins_270),
    .io_ins_271(rport_io_ins_271),
    .io_ins_272(rport_io_ins_272),
    .io_ins_273(rport_io_ins_273),
    .io_ins_274(rport_io_ins_274),
    .io_ins_275(rport_io_ins_275),
    .io_ins_276(rport_io_ins_276),
    .io_ins_277(rport_io_ins_277),
    .io_ins_278(rport_io_ins_278),
    .io_ins_279(rport_io_ins_279),
    .io_ins_280(rport_io_ins_280),
    .io_ins_281(rport_io_ins_281),
    .io_ins_282(rport_io_ins_282),
    .io_ins_283(rport_io_ins_283),
    .io_ins_284(rport_io_ins_284),
    .io_ins_285(rport_io_ins_285),
    .io_ins_286(rport_io_ins_286),
    .io_ins_287(rport_io_ins_287),
    .io_ins_288(rport_io_ins_288),
    .io_ins_289(rport_io_ins_289),
    .io_ins_290(rport_io_ins_290),
    .io_ins_291(rport_io_ins_291),
    .io_ins_292(rport_io_ins_292),
    .io_ins_293(rport_io_ins_293),
    .io_ins_294(rport_io_ins_294),
    .io_ins_295(rport_io_ins_295),
    .io_ins_296(rport_io_ins_296),
    .io_ins_297(rport_io_ins_297),
    .io_ins_298(rport_io_ins_298),
    .io_ins_299(rport_io_ins_299),
    .io_ins_300(rport_io_ins_300),
    .io_ins_301(rport_io_ins_301),
    .io_ins_302(rport_io_ins_302),
    .io_ins_303(rport_io_ins_303),
    .io_ins_304(rport_io_ins_304),
    .io_ins_305(rport_io_ins_305),
    .io_ins_306(rport_io_ins_306),
    .io_ins_307(rport_io_ins_307),
    .io_ins_308(rport_io_ins_308),
    .io_ins_309(rport_io_ins_309),
    .io_ins_310(rport_io_ins_310),
    .io_ins_311(rport_io_ins_311),
    .io_ins_312(rport_io_ins_312),
    .io_ins_313(rport_io_ins_313),
    .io_ins_314(rport_io_ins_314),
    .io_ins_315(rport_io_ins_315),
    .io_ins_316(rport_io_ins_316),
    .io_ins_317(rport_io_ins_317),
    .io_ins_318(rport_io_ins_318),
    .io_ins_319(rport_io_ins_319),
    .io_ins_320(rport_io_ins_320),
    .io_ins_321(rport_io_ins_321),
    .io_ins_322(rport_io_ins_322),
    .io_ins_323(rport_io_ins_323),
    .io_ins_324(rport_io_ins_324),
    .io_ins_325(rport_io_ins_325),
    .io_ins_326(rport_io_ins_326),
    .io_ins_327(rport_io_ins_327),
    .io_ins_328(rport_io_ins_328),
    .io_ins_329(rport_io_ins_329),
    .io_ins_330(rport_io_ins_330),
    .io_ins_331(rport_io_ins_331),
    .io_ins_332(rport_io_ins_332),
    .io_ins_333(rport_io_ins_333),
    .io_ins_334(rport_io_ins_334),
    .io_ins_335(rport_io_ins_335),
    .io_ins_336(rport_io_ins_336),
    .io_ins_337(rport_io_ins_337),
    .io_ins_338(rport_io_ins_338),
    .io_ins_339(rport_io_ins_339),
    .io_ins_340(rport_io_ins_340),
    .io_ins_341(rport_io_ins_341),
    .io_ins_342(rport_io_ins_342),
    .io_ins_343(rport_io_ins_343),
    .io_ins_344(rport_io_ins_344),
    .io_ins_345(rport_io_ins_345),
    .io_ins_346(rport_io_ins_346),
    .io_ins_347(rport_io_ins_347),
    .io_ins_348(rport_io_ins_348),
    .io_ins_349(rport_io_ins_349),
    .io_ins_350(rport_io_ins_350),
    .io_ins_351(rport_io_ins_351),
    .io_ins_352(rport_io_ins_352),
    .io_ins_353(rport_io_ins_353),
    .io_ins_354(rport_io_ins_354),
    .io_ins_355(rport_io_ins_355),
    .io_ins_356(rport_io_ins_356),
    .io_ins_357(rport_io_ins_357),
    .io_ins_358(rport_io_ins_358),
    .io_ins_359(rport_io_ins_359),
    .io_ins_360(rport_io_ins_360),
    .io_ins_361(rport_io_ins_361),
    .io_ins_362(rport_io_ins_362),
    .io_ins_363(rport_io_ins_363),
    .io_ins_364(rport_io_ins_364),
    .io_ins_365(rport_io_ins_365),
    .io_ins_366(rport_io_ins_366),
    .io_ins_367(rport_io_ins_367),
    .io_ins_368(rport_io_ins_368),
    .io_ins_369(rport_io_ins_369),
    .io_ins_370(rport_io_ins_370),
    .io_ins_371(rport_io_ins_371),
    .io_ins_372(rport_io_ins_372),
    .io_ins_373(rport_io_ins_373),
    .io_ins_374(rport_io_ins_374),
    .io_ins_375(rport_io_ins_375),
    .io_ins_376(rport_io_ins_376),
    .io_ins_377(rport_io_ins_377),
    .io_ins_378(rport_io_ins_378),
    .io_ins_379(rport_io_ins_379),
    .io_ins_380(rport_io_ins_380),
    .io_ins_381(rport_io_ins_381),
    .io_ins_382(rport_io_ins_382),
    .io_ins_383(rport_io_ins_383),
    .io_ins_384(rport_io_ins_384),
    .io_ins_385(rport_io_ins_385),
    .io_ins_386(rport_io_ins_386),
    .io_ins_387(rport_io_ins_387),
    .io_ins_388(rport_io_ins_388),
    .io_ins_389(rport_io_ins_389),
    .io_ins_390(rport_io_ins_390),
    .io_ins_391(rport_io_ins_391),
    .io_ins_392(rport_io_ins_392),
    .io_ins_393(rport_io_ins_393),
    .io_ins_394(rport_io_ins_394),
    .io_ins_395(rport_io_ins_395),
    .io_ins_396(rport_io_ins_396),
    .io_ins_397(rport_io_ins_397),
    .io_ins_398(rport_io_ins_398),
    .io_ins_399(rport_io_ins_399),
    .io_ins_400(rport_io_ins_400),
    .io_ins_401(rport_io_ins_401),
    .io_ins_402(rport_io_ins_402),
    .io_ins_403(rport_io_ins_403),
    .io_ins_404(rport_io_ins_404),
    .io_ins_405(rport_io_ins_405),
    .io_ins_406(rport_io_ins_406),
    .io_ins_407(rport_io_ins_407),
    .io_ins_408(rport_io_ins_408),
    .io_ins_409(rport_io_ins_409),
    .io_ins_410(rport_io_ins_410),
    .io_ins_411(rport_io_ins_411),
    .io_ins_412(rport_io_ins_412),
    .io_ins_413(rport_io_ins_413),
    .io_ins_414(rport_io_ins_414),
    .io_ins_415(rport_io_ins_415),
    .io_ins_416(rport_io_ins_416),
    .io_ins_417(rport_io_ins_417),
    .io_ins_418(rport_io_ins_418),
    .io_ins_419(rport_io_ins_419),
    .io_ins_420(rport_io_ins_420),
    .io_ins_421(rport_io_ins_421),
    .io_ins_422(rport_io_ins_422),
    .io_ins_423(rport_io_ins_423),
    .io_ins_424(rport_io_ins_424),
    .io_ins_425(rport_io_ins_425),
    .io_ins_426(rport_io_ins_426),
    .io_ins_427(rport_io_ins_427),
    .io_ins_428(rport_io_ins_428),
    .io_ins_429(rport_io_ins_429),
    .io_ins_430(rport_io_ins_430),
    .io_ins_431(rport_io_ins_431),
    .io_ins_432(rport_io_ins_432),
    .io_ins_433(rport_io_ins_433),
    .io_ins_434(rport_io_ins_434),
    .io_ins_435(rport_io_ins_435),
    .io_ins_436(rport_io_ins_436),
    .io_ins_437(rport_io_ins_437),
    .io_ins_438(rport_io_ins_438),
    .io_ins_439(rport_io_ins_439),
    .io_ins_440(rport_io_ins_440),
    .io_ins_441(rport_io_ins_441),
    .io_ins_442(rport_io_ins_442),
    .io_ins_443(rport_io_ins_443),
    .io_ins_444(rport_io_ins_444),
    .io_ins_445(rport_io_ins_445),
    .io_ins_446(rport_io_ins_446),
    .io_ins_447(rport_io_ins_447),
    .io_ins_448(rport_io_ins_448),
    .io_ins_449(rport_io_ins_449),
    .io_ins_450(rport_io_ins_450),
    .io_ins_451(rport_io_ins_451),
    .io_ins_452(rport_io_ins_452),
    .io_ins_453(rport_io_ins_453),
    .io_ins_454(rport_io_ins_454),
    .io_ins_455(rport_io_ins_455),
    .io_ins_456(rport_io_ins_456),
    .io_ins_457(rport_io_ins_457),
    .io_ins_458(rport_io_ins_458),
    .io_ins_459(rport_io_ins_459),
    .io_ins_460(rport_io_ins_460),
    .io_ins_461(rport_io_ins_461),
    .io_ins_462(rport_io_ins_462),
    .io_ins_463(rport_io_ins_463),
    .io_ins_464(rport_io_ins_464),
    .io_ins_465(rport_io_ins_465),
    .io_ins_466(rport_io_ins_466),
    .io_ins_467(rport_io_ins_467),
    .io_ins_468(rport_io_ins_468),
    .io_ins_469(rport_io_ins_469),
    .io_ins_470(rport_io_ins_470),
    .io_ins_471(rport_io_ins_471),
    .io_ins_472(rport_io_ins_472),
    .io_ins_473(rport_io_ins_473),
    .io_ins_474(rport_io_ins_474),
    .io_ins_475(rport_io_ins_475),
    .io_ins_476(rport_io_ins_476),
    .io_ins_477(rport_io_ins_477),
    .io_ins_478(rport_io_ins_478),
    .io_ins_479(rport_io_ins_479),
    .io_ins_480(rport_io_ins_480),
    .io_ins_481(rport_io_ins_481),
    .io_ins_482(rport_io_ins_482),
    .io_ins_483(rport_io_ins_483),
    .io_ins_484(rport_io_ins_484),
    .io_ins_485(rport_io_ins_485),
    .io_ins_486(rport_io_ins_486),
    .io_ins_487(rport_io_ins_487),
    .io_ins_488(rport_io_ins_488),
    .io_ins_489(rport_io_ins_489),
    .io_ins_490(rport_io_ins_490),
    .io_ins_491(rport_io_ins_491),
    .io_ins_492(rport_io_ins_492),
    .io_ins_493(rport_io_ins_493),
    .io_ins_494(rport_io_ins_494),
    .io_ins_495(rport_io_ins_495),
    .io_ins_496(rport_io_ins_496),
    .io_ins_497(rport_io_ins_497),
    .io_ins_498(rport_io_ins_498),
    .io_ins_499(rport_io_ins_499),
    .io_ins_500(rport_io_ins_500),
    .io_ins_501(rport_io_ins_501),
    .io_ins_502(rport_io_ins_502),
    .io_ins_503(rport_io_ins_503),
    .io_ins_504(rport_io_ins_504),
    .io_ins_505(rport_io_ins_505),
    .io_ins_506(rport_io_ins_506),
    .io_ins_507(rport_io_ins_507),
    .io_ins_508(rport_io_ins_508),
    .io_ins_509(rport_io_ins_509),
    .io_ins_510(rport_io_ins_510),
    .io_ins_511(rport_io_ins_511),
    .io_ins_512(rport_io_ins_512),
    .io_ins_513(rport_io_ins_513),
    .io_ins_514(rport_io_ins_514),
    .io_ins_515(rport_io_ins_515),
    .io_ins_516(rport_io_ins_516),
    .io_ins_517(rport_io_ins_517),
    .io_ins_518(rport_io_ins_518),
    .io_ins_519(rport_io_ins_519),
    .io_ins_520(rport_io_ins_520),
    .io_ins_521(rport_io_ins_521),
    .io_sel(rport_io_sel),
    .io_out(rport_io_out)
  );
  assign _T_3190 = io_waddr == 32'h0; // @[RegFile.scala 80:42:@41890.4]
  assign _T_3196 = io_waddr == 32'h1; // @[RegFile.scala 68:46:@41902.4]
  assign _T_3197 = io_wen & _T_3196; // @[RegFile.scala 68:34:@41903.4]
  assign _T_3210 = io_waddr == 32'h2; // @[RegFile.scala 80:42:@41921.4]
  assign _T_3216 = io_waddr == 32'h3; // @[RegFile.scala 74:80:@41933.4]
  assign _T_3217 = io_wen & _T_3216; // @[RegFile.scala 74:68:@41934.4]
  assign _T_3223 = io_waddr == 32'h4; // @[RegFile.scala 74:80:@41947.4]
  assign _T_3224 = io_wen & _T_3223; // @[RegFile.scala 74:68:@41948.4]
  assign _T_3230 = io_waddr == 32'h5; // @[RegFile.scala 74:80:@41961.4]
  assign _T_3231 = io_wen & _T_3230; // @[RegFile.scala 74:68:@41962.4]
  assign _T_3237 = io_waddr == 32'h6; // @[RegFile.scala 74:80:@41975.4]
  assign _T_3238 = io_wen & _T_3237; // @[RegFile.scala 74:68:@41976.4]
  assign _T_3244 = io_waddr == 32'h7; // @[RegFile.scala 74:80:@41989.4]
  assign _T_3245 = io_wen & _T_3244; // @[RegFile.scala 74:68:@41990.4]
  assign _T_3251 = io_waddr == 32'h8; // @[RegFile.scala 74:80:@42003.4]
  assign _T_3252 = io_wen & _T_3251; // @[RegFile.scala 74:68:@42004.4]
  assign _T_3258 = io_waddr == 32'h9; // @[RegFile.scala 74:80:@42017.4]
  assign _T_3259 = io_wen & _T_3258; // @[RegFile.scala 74:68:@42018.4]
  assign _T_3265 = io_waddr == 32'ha; // @[RegFile.scala 74:80:@42031.4]
  assign _T_3266 = io_wen & _T_3265; // @[RegFile.scala 74:68:@42032.4]
  assign _T_3272 = io_waddr == 32'hb; // @[RegFile.scala 74:80:@42045.4]
  assign _T_3273 = io_wen & _T_3272; // @[RegFile.scala 74:68:@42046.4]
  assign _T_3279 = io_waddr == 32'hc; // @[RegFile.scala 74:80:@42059.4]
  assign _T_3280 = io_wen & _T_3279; // @[RegFile.scala 74:68:@42060.4]
  assign _T_3286 = io_waddr == 32'hd; // @[RegFile.scala 74:80:@42073.4]
  assign _T_3287 = io_wen & _T_3286; // @[RegFile.scala 74:68:@42074.4]
  assign _T_3293 = io_waddr == 32'he; // @[RegFile.scala 74:80:@42087.4]
  assign _T_3294 = io_wen & _T_3293; // @[RegFile.scala 74:68:@42088.4]
  assign _T_3300 = io_waddr == 32'hf; // @[RegFile.scala 74:80:@42101.4]
  assign _T_3301 = io_wen & _T_3300; // @[RegFile.scala 74:68:@42102.4]
  assign _T_3307 = io_waddr == 32'h10; // @[RegFile.scala 74:80:@42115.4]
  assign _T_3308 = io_wen & _T_3307; // @[RegFile.scala 74:68:@42116.4]
  assign _T_3314 = io_waddr == 32'h11; // @[RegFile.scala 74:80:@42129.4]
  assign _T_3315 = io_wen & _T_3314; // @[RegFile.scala 74:68:@42130.4]
  assign _T_3321 = io_waddr == 32'h12; // @[RegFile.scala 74:80:@42143.4]
  assign _T_3322 = io_wen & _T_3321; // @[RegFile.scala 74:68:@42144.4]
  assign _T_3328 = io_waddr == 32'h13; // @[RegFile.scala 74:80:@42157.4]
  assign _T_3329 = io_wen & _T_3328; // @[RegFile.scala 74:68:@42158.4]
  assign _T_3335 = io_waddr == 32'h14; // @[RegFile.scala 74:80:@42171.4]
  assign _T_3336 = io_wen & _T_3335; // @[RegFile.scala 74:68:@42172.4]
  assign _T_3342 = io_waddr == 32'h15; // @[RegFile.scala 74:80:@42185.4]
  assign _T_3343 = io_wen & _T_3342; // @[RegFile.scala 74:68:@42186.4]
  assign _T_3349 = io_waddr == 32'h16; // @[RegFile.scala 74:80:@42199.4]
  assign _T_3350 = io_wen & _T_3349; // @[RegFile.scala 74:68:@42200.4]
  assign io_rdata = rport_io_out; // @[RegFile.scala 107:14:@50245.4]
  assign io_argIns_0 = regs_0_io_out; // @[RegFile.scala 111:13:@50250.4]
  assign io_argIns_1 = regs_1_io_out; // @[RegFile.scala 111:13:@50251.4]
  assign io_argIns_2 = regs_2_io_out; // @[RegFile.scala 111:13:@50252.4]
  assign regs_0_clock = clock; // @[:@41888.4]
  assign regs_0_reset = reset; // @[:@41889.4 RegFile.scala 82:16:@41895.4]
  assign regs_0_io_in = io_wdata; // @[RegFile.scala 81:16:@41893.4]
  assign regs_0_io_reset = reset; // @[RegFile.scala 83:19:@41897.4]
  assign regs_0_io_enable = io_wen & _T_3190; // @[RegFile.scala 80:20:@41892.4]
  assign regs_1_clock = clock; // @[:@41900.4]
  assign regs_1_reset = reset; // @[:@41901.4 RegFile.scala 70:16:@41913.4]
  assign regs_1_io_in = _T_3197 ? io_wdata : io_argOuts_0_bits; // @[RegFile.scala 69:16:@41911.4]
  assign regs_1_io_reset = reset; // @[RegFile.scala 72:19:@41916.4]
  assign regs_1_io_enable = _T_3197 ? _T_3197 : io_argOuts_0_valid; // @[RegFile.scala 68:20:@41907.4]
  assign regs_2_clock = clock; // @[:@41919.4]
  assign regs_2_reset = reset; // @[:@41920.4 RegFile.scala 82:16:@41926.4]
  assign regs_2_io_in = io_wdata; // @[RegFile.scala 81:16:@41924.4]
  assign regs_2_io_reset = reset; // @[RegFile.scala 83:19:@41928.4]
  assign regs_2_io_enable = io_wen & _T_3210; // @[RegFile.scala 80:20:@41923.4]
  assign regs_3_clock = clock; // @[:@41931.4]
  assign regs_3_reset = io_reset; // @[:@41932.4 RegFile.scala 76:16:@41939.4]
  assign regs_3_io_in = io_argOuts_1_valid ? io_argOuts_1_bits : io_wdata; // @[RegFile.scala 75:16:@41938.4]
  assign regs_3_io_reset = reset; // @[RegFile.scala 78:19:@41942.4]
  assign regs_3_io_enable = io_argOuts_1_valid | _T_3217; // @[RegFile.scala 74:20:@41936.4]
  assign regs_4_clock = clock; // @[:@41945.4]
  assign regs_4_reset = io_reset; // @[:@41946.4 RegFile.scala 76:16:@41953.4]
  assign regs_4_io_in = io_argOuts_2_valid ? io_argOuts_2_bits : io_wdata; // @[RegFile.scala 75:16:@41952.4]
  assign regs_4_io_reset = reset; // @[RegFile.scala 78:19:@41956.4]
  assign regs_4_io_enable = io_argOuts_2_valid | _T_3224; // @[RegFile.scala 74:20:@41950.4]
  assign regs_5_clock = clock; // @[:@41959.4]
  assign regs_5_reset = io_reset; // @[:@41960.4 RegFile.scala 76:16:@41967.4]
  assign regs_5_io_in = io_argOuts_3_valid ? io_argOuts_3_bits : io_wdata; // @[RegFile.scala 75:16:@41966.4]
  assign regs_5_io_reset = reset; // @[RegFile.scala 78:19:@41970.4]
  assign regs_5_io_enable = io_argOuts_3_valid | _T_3231; // @[RegFile.scala 74:20:@41964.4]
  assign regs_6_clock = clock; // @[:@41973.4]
  assign regs_6_reset = io_reset; // @[:@41974.4 RegFile.scala 76:16:@41981.4]
  assign regs_6_io_in = io_argOuts_4_valid ? io_argOuts_4_bits : io_wdata; // @[RegFile.scala 75:16:@41980.4]
  assign regs_6_io_reset = reset; // @[RegFile.scala 78:19:@41984.4]
  assign regs_6_io_enable = io_argOuts_4_valid | _T_3238; // @[RegFile.scala 74:20:@41978.4]
  assign regs_7_clock = clock; // @[:@41987.4]
  assign regs_7_reset = io_reset; // @[:@41988.4 RegFile.scala 76:16:@41995.4]
  assign regs_7_io_in = io_argOuts_5_valid ? io_argOuts_5_bits : io_wdata; // @[RegFile.scala 75:16:@41994.4]
  assign regs_7_io_reset = reset; // @[RegFile.scala 78:19:@41998.4]
  assign regs_7_io_enable = io_argOuts_5_valid | _T_3245; // @[RegFile.scala 74:20:@41992.4]
  assign regs_8_clock = clock; // @[:@42001.4]
  assign regs_8_reset = io_reset; // @[:@42002.4 RegFile.scala 76:16:@42009.4]
  assign regs_8_io_in = io_argOuts_6_valid ? io_argOuts_6_bits : io_wdata; // @[RegFile.scala 75:16:@42008.4]
  assign regs_8_io_reset = reset; // @[RegFile.scala 78:19:@42012.4]
  assign regs_8_io_enable = io_argOuts_6_valid | _T_3252; // @[RegFile.scala 74:20:@42006.4]
  assign regs_9_clock = clock; // @[:@42015.4]
  assign regs_9_reset = io_reset; // @[:@42016.4 RegFile.scala 76:16:@42023.4]
  assign regs_9_io_in = io_argOuts_7_valid ? io_argOuts_7_bits : io_wdata; // @[RegFile.scala 75:16:@42022.4]
  assign regs_9_io_reset = reset; // @[RegFile.scala 78:19:@42026.4]
  assign regs_9_io_enable = io_argOuts_7_valid | _T_3259; // @[RegFile.scala 74:20:@42020.4]
  assign regs_10_clock = clock; // @[:@42029.4]
  assign regs_10_reset = io_reset; // @[:@42030.4 RegFile.scala 76:16:@42037.4]
  assign regs_10_io_in = io_argOuts_8_valid ? io_argOuts_8_bits : io_wdata; // @[RegFile.scala 75:16:@42036.4]
  assign regs_10_io_reset = reset; // @[RegFile.scala 78:19:@42040.4]
  assign regs_10_io_enable = io_argOuts_8_valid | _T_3266; // @[RegFile.scala 74:20:@42034.4]
  assign regs_11_clock = clock; // @[:@42043.4]
  assign regs_11_reset = io_reset; // @[:@42044.4 RegFile.scala 76:16:@42051.4]
  assign regs_11_io_in = io_argOuts_9_valid ? io_argOuts_9_bits : io_wdata; // @[RegFile.scala 75:16:@42050.4]
  assign regs_11_io_reset = reset; // @[RegFile.scala 78:19:@42054.4]
  assign regs_11_io_enable = io_argOuts_9_valid | _T_3273; // @[RegFile.scala 74:20:@42048.4]
  assign regs_12_clock = clock; // @[:@42057.4]
  assign regs_12_reset = io_reset; // @[:@42058.4 RegFile.scala 76:16:@42065.4]
  assign regs_12_io_in = io_argOuts_10_valid ? io_argOuts_10_bits : io_wdata; // @[RegFile.scala 75:16:@42064.4]
  assign regs_12_io_reset = reset; // @[RegFile.scala 78:19:@42068.4]
  assign regs_12_io_enable = io_argOuts_10_valid | _T_3280; // @[RegFile.scala 74:20:@42062.4]
  assign regs_13_clock = clock; // @[:@42071.4]
  assign regs_13_reset = io_reset; // @[:@42072.4 RegFile.scala 76:16:@42079.4]
  assign regs_13_io_in = io_argOuts_11_valid ? io_argOuts_11_bits : io_wdata; // @[RegFile.scala 75:16:@42078.4]
  assign regs_13_io_reset = reset; // @[RegFile.scala 78:19:@42082.4]
  assign regs_13_io_enable = io_argOuts_11_valid | _T_3287; // @[RegFile.scala 74:20:@42076.4]
  assign regs_14_clock = clock; // @[:@42085.4]
  assign regs_14_reset = io_reset; // @[:@42086.4 RegFile.scala 76:16:@42093.4]
  assign regs_14_io_in = io_argOuts_12_valid ? io_argOuts_12_bits : io_wdata; // @[RegFile.scala 75:16:@42092.4]
  assign regs_14_io_reset = reset; // @[RegFile.scala 78:19:@42096.4]
  assign regs_14_io_enable = io_argOuts_12_valid | _T_3294; // @[RegFile.scala 74:20:@42090.4]
  assign regs_15_clock = clock; // @[:@42099.4]
  assign regs_15_reset = io_reset; // @[:@42100.4 RegFile.scala 76:16:@42107.4]
  assign regs_15_io_in = io_argOuts_13_valid ? io_argOuts_13_bits : io_wdata; // @[RegFile.scala 75:16:@42106.4]
  assign regs_15_io_reset = reset; // @[RegFile.scala 78:19:@42110.4]
  assign regs_15_io_enable = io_argOuts_13_valid | _T_3301; // @[RegFile.scala 74:20:@42104.4]
  assign regs_16_clock = clock; // @[:@42113.4]
  assign regs_16_reset = io_reset; // @[:@42114.4 RegFile.scala 76:16:@42121.4]
  assign regs_16_io_in = io_argOuts_14_valid ? io_argOuts_14_bits : io_wdata; // @[RegFile.scala 75:16:@42120.4]
  assign regs_16_io_reset = reset; // @[RegFile.scala 78:19:@42124.4]
  assign regs_16_io_enable = io_argOuts_14_valid | _T_3308; // @[RegFile.scala 74:20:@42118.4]
  assign regs_17_clock = clock; // @[:@42127.4]
  assign regs_17_reset = io_reset; // @[:@42128.4 RegFile.scala 76:16:@42135.4]
  assign regs_17_io_in = io_argOuts_15_valid ? io_argOuts_15_bits : io_wdata; // @[RegFile.scala 75:16:@42134.4]
  assign regs_17_io_reset = reset; // @[RegFile.scala 78:19:@42138.4]
  assign regs_17_io_enable = io_argOuts_15_valid | _T_3315; // @[RegFile.scala 74:20:@42132.4]
  assign regs_18_clock = clock; // @[:@42141.4]
  assign regs_18_reset = io_reset; // @[:@42142.4 RegFile.scala 76:16:@42149.4]
  assign regs_18_io_in = io_argOuts_16_valid ? io_argOuts_16_bits : io_wdata; // @[RegFile.scala 75:16:@42148.4]
  assign regs_18_io_reset = reset; // @[RegFile.scala 78:19:@42152.4]
  assign regs_18_io_enable = io_argOuts_16_valid | _T_3322; // @[RegFile.scala 74:20:@42146.4]
  assign regs_19_clock = clock; // @[:@42155.4]
  assign regs_19_reset = io_reset; // @[:@42156.4 RegFile.scala 76:16:@42163.4]
  assign regs_19_io_in = io_argOuts_17_valid ? io_argOuts_17_bits : io_wdata; // @[RegFile.scala 75:16:@42162.4]
  assign regs_19_io_reset = reset; // @[RegFile.scala 78:19:@42166.4]
  assign regs_19_io_enable = io_argOuts_17_valid | _T_3329; // @[RegFile.scala 74:20:@42160.4]
  assign regs_20_clock = clock; // @[:@42169.4]
  assign regs_20_reset = io_reset; // @[:@42170.4 RegFile.scala 76:16:@42177.4]
  assign regs_20_io_in = io_argOuts_18_valid ? io_argOuts_18_bits : io_wdata; // @[RegFile.scala 75:16:@42176.4]
  assign regs_20_io_reset = reset; // @[RegFile.scala 78:19:@42180.4]
  assign regs_20_io_enable = io_argOuts_18_valid | _T_3336; // @[RegFile.scala 74:20:@42174.4]
  assign regs_21_clock = clock; // @[:@42183.4]
  assign regs_21_reset = io_reset; // @[:@42184.4 RegFile.scala 76:16:@42191.4]
  assign regs_21_io_in = io_argOuts_19_valid ? io_argOuts_19_bits : io_wdata; // @[RegFile.scala 75:16:@42190.4]
  assign regs_21_io_reset = reset; // @[RegFile.scala 78:19:@42194.4]
  assign regs_21_io_enable = io_argOuts_19_valid | _T_3343; // @[RegFile.scala 74:20:@42188.4]
  assign regs_22_clock = clock; // @[:@42197.4]
  assign regs_22_reset = io_reset; // @[:@42198.4 RegFile.scala 76:16:@42205.4]
  assign regs_22_io_in = io_argOuts_20_valid ? io_argOuts_20_bits : io_wdata; // @[RegFile.scala 75:16:@42204.4]
  assign regs_22_io_reset = reset; // @[RegFile.scala 78:19:@42208.4]
  assign regs_22_io_enable = io_argOuts_20_valid | _T_3350; // @[RegFile.scala 74:20:@42202.4]
  assign regs_23_clock = clock; // @[:@42211.4]
  assign regs_23_reset = io_reset; // @[:@42212.4 RegFile.scala 76:16:@42219.4]
  assign regs_23_io_in = 64'h0; // @[RegFile.scala 75:16:@42218.4]
  assign regs_23_io_reset = reset; // @[RegFile.scala 78:19:@42222.4]
  assign regs_23_io_enable = 1'h1; // @[RegFile.scala 74:20:@42216.4]
  assign regs_24_clock = clock; // @[:@42225.4]
  assign regs_24_reset = io_reset; // @[:@42226.4 RegFile.scala 76:16:@42233.4]
  assign regs_24_io_in = 64'h0; // @[RegFile.scala 75:16:@42232.4]
  assign regs_24_io_reset = reset; // @[RegFile.scala 78:19:@42236.4]
  assign regs_24_io_enable = 1'h1; // @[RegFile.scala 74:20:@42230.4]
  assign regs_25_clock = clock; // @[:@42239.4]
  assign regs_25_reset = io_reset; // @[:@42240.4 RegFile.scala 76:16:@42247.4]
  assign regs_25_io_in = 64'h0; // @[RegFile.scala 75:16:@42246.4]
  assign regs_25_io_reset = reset; // @[RegFile.scala 78:19:@42250.4]
  assign regs_25_io_enable = 1'h1; // @[RegFile.scala 74:20:@42244.4]
  assign regs_26_clock = clock; // @[:@42253.4]
  assign regs_26_reset = io_reset; // @[:@42254.4 RegFile.scala 76:16:@42261.4]
  assign regs_26_io_in = 64'h0; // @[RegFile.scala 75:16:@42260.4]
  assign regs_26_io_reset = reset; // @[RegFile.scala 78:19:@42264.4]
  assign regs_26_io_enable = 1'h1; // @[RegFile.scala 74:20:@42258.4]
  assign regs_27_clock = clock; // @[:@42267.4]
  assign regs_27_reset = io_reset; // @[:@42268.4 RegFile.scala 76:16:@42275.4]
  assign regs_27_io_in = 64'h0; // @[RegFile.scala 75:16:@42274.4]
  assign regs_27_io_reset = reset; // @[RegFile.scala 78:19:@42278.4]
  assign regs_27_io_enable = 1'h1; // @[RegFile.scala 74:20:@42272.4]
  assign regs_28_clock = clock; // @[:@42281.4]
  assign regs_28_reset = io_reset; // @[:@42282.4 RegFile.scala 76:16:@42289.4]
  assign regs_28_io_in = 64'h0; // @[RegFile.scala 75:16:@42288.4]
  assign regs_28_io_reset = reset; // @[RegFile.scala 78:19:@42292.4]
  assign regs_28_io_enable = 1'h1; // @[RegFile.scala 74:20:@42286.4]
  assign regs_29_clock = clock; // @[:@42295.4]
  assign regs_29_reset = io_reset; // @[:@42296.4 RegFile.scala 76:16:@42303.4]
  assign regs_29_io_in = 64'h0; // @[RegFile.scala 75:16:@42302.4]
  assign regs_29_io_reset = reset; // @[RegFile.scala 78:19:@42306.4]
  assign regs_29_io_enable = 1'h1; // @[RegFile.scala 74:20:@42300.4]
  assign regs_30_clock = clock; // @[:@42309.4]
  assign regs_30_reset = io_reset; // @[:@42310.4 RegFile.scala 76:16:@42317.4]
  assign regs_30_io_in = 64'h0; // @[RegFile.scala 75:16:@42316.4]
  assign regs_30_io_reset = reset; // @[RegFile.scala 78:19:@42320.4]
  assign regs_30_io_enable = 1'h1; // @[RegFile.scala 74:20:@42314.4]
  assign regs_31_clock = clock; // @[:@42323.4]
  assign regs_31_reset = io_reset; // @[:@42324.4 RegFile.scala 76:16:@42331.4]
  assign regs_31_io_in = 64'h0; // @[RegFile.scala 75:16:@42330.4]
  assign regs_31_io_reset = reset; // @[RegFile.scala 78:19:@42334.4]
  assign regs_31_io_enable = 1'h1; // @[RegFile.scala 74:20:@42328.4]
  assign regs_32_clock = clock; // @[:@42337.4]
  assign regs_32_reset = io_reset; // @[:@42338.4 RegFile.scala 76:16:@42345.4]
  assign regs_32_io_in = 64'h0; // @[RegFile.scala 75:16:@42344.4]
  assign regs_32_io_reset = reset; // @[RegFile.scala 78:19:@42348.4]
  assign regs_32_io_enable = 1'h1; // @[RegFile.scala 74:20:@42342.4]
  assign regs_33_clock = clock; // @[:@42351.4]
  assign regs_33_reset = io_reset; // @[:@42352.4 RegFile.scala 76:16:@42359.4]
  assign regs_33_io_in = 64'h0; // @[RegFile.scala 75:16:@42358.4]
  assign regs_33_io_reset = reset; // @[RegFile.scala 78:19:@42362.4]
  assign regs_33_io_enable = 1'h1; // @[RegFile.scala 74:20:@42356.4]
  assign regs_34_clock = clock; // @[:@42365.4]
  assign regs_34_reset = io_reset; // @[:@42366.4 RegFile.scala 76:16:@42373.4]
  assign regs_34_io_in = 64'h0; // @[RegFile.scala 75:16:@42372.4]
  assign regs_34_io_reset = reset; // @[RegFile.scala 78:19:@42376.4]
  assign regs_34_io_enable = 1'h1; // @[RegFile.scala 74:20:@42370.4]
  assign regs_35_clock = clock; // @[:@42379.4]
  assign regs_35_reset = io_reset; // @[:@42380.4 RegFile.scala 76:16:@42387.4]
  assign regs_35_io_in = 64'h0; // @[RegFile.scala 75:16:@42386.4]
  assign regs_35_io_reset = reset; // @[RegFile.scala 78:19:@42390.4]
  assign regs_35_io_enable = 1'h1; // @[RegFile.scala 74:20:@42384.4]
  assign regs_36_clock = clock; // @[:@42393.4]
  assign regs_36_reset = io_reset; // @[:@42394.4 RegFile.scala 76:16:@42401.4]
  assign regs_36_io_in = 64'h0; // @[RegFile.scala 75:16:@42400.4]
  assign regs_36_io_reset = reset; // @[RegFile.scala 78:19:@42404.4]
  assign regs_36_io_enable = 1'h1; // @[RegFile.scala 74:20:@42398.4]
  assign regs_37_clock = clock; // @[:@42407.4]
  assign regs_37_reset = io_reset; // @[:@42408.4 RegFile.scala 76:16:@42415.4]
  assign regs_37_io_in = 64'h0; // @[RegFile.scala 75:16:@42414.4]
  assign regs_37_io_reset = reset; // @[RegFile.scala 78:19:@42418.4]
  assign regs_37_io_enable = 1'h1; // @[RegFile.scala 74:20:@42412.4]
  assign regs_38_clock = clock; // @[:@42421.4]
  assign regs_38_reset = io_reset; // @[:@42422.4 RegFile.scala 76:16:@42429.4]
  assign regs_38_io_in = 64'h0; // @[RegFile.scala 75:16:@42428.4]
  assign regs_38_io_reset = reset; // @[RegFile.scala 78:19:@42432.4]
  assign regs_38_io_enable = 1'h1; // @[RegFile.scala 74:20:@42426.4]
  assign regs_39_clock = clock; // @[:@42435.4]
  assign regs_39_reset = io_reset; // @[:@42436.4 RegFile.scala 76:16:@42443.4]
  assign regs_39_io_in = 64'h0; // @[RegFile.scala 75:16:@42442.4]
  assign regs_39_io_reset = reset; // @[RegFile.scala 78:19:@42446.4]
  assign regs_39_io_enable = 1'h1; // @[RegFile.scala 74:20:@42440.4]
  assign regs_40_clock = clock; // @[:@42449.4]
  assign regs_40_reset = io_reset; // @[:@42450.4 RegFile.scala 76:16:@42457.4]
  assign regs_40_io_in = 64'h0; // @[RegFile.scala 75:16:@42456.4]
  assign regs_40_io_reset = reset; // @[RegFile.scala 78:19:@42460.4]
  assign regs_40_io_enable = 1'h1; // @[RegFile.scala 74:20:@42454.4]
  assign regs_41_clock = clock; // @[:@42463.4]
  assign regs_41_reset = io_reset; // @[:@42464.4 RegFile.scala 76:16:@42471.4]
  assign regs_41_io_in = 64'h0; // @[RegFile.scala 75:16:@42470.4]
  assign regs_41_io_reset = reset; // @[RegFile.scala 78:19:@42474.4]
  assign regs_41_io_enable = 1'h1; // @[RegFile.scala 74:20:@42468.4]
  assign regs_42_clock = clock; // @[:@42477.4]
  assign regs_42_reset = io_reset; // @[:@42478.4 RegFile.scala 76:16:@42485.4]
  assign regs_42_io_in = 64'h0; // @[RegFile.scala 75:16:@42484.4]
  assign regs_42_io_reset = reset; // @[RegFile.scala 78:19:@42488.4]
  assign regs_42_io_enable = 1'h1; // @[RegFile.scala 74:20:@42482.4]
  assign regs_43_clock = clock; // @[:@42491.4]
  assign regs_43_reset = io_reset; // @[:@42492.4 RegFile.scala 76:16:@42499.4]
  assign regs_43_io_in = 64'h0; // @[RegFile.scala 75:16:@42498.4]
  assign regs_43_io_reset = reset; // @[RegFile.scala 78:19:@42502.4]
  assign regs_43_io_enable = 1'h1; // @[RegFile.scala 74:20:@42496.4]
  assign regs_44_clock = clock; // @[:@42505.4]
  assign regs_44_reset = io_reset; // @[:@42506.4 RegFile.scala 76:16:@42513.4]
  assign regs_44_io_in = 64'h0; // @[RegFile.scala 75:16:@42512.4]
  assign regs_44_io_reset = reset; // @[RegFile.scala 78:19:@42516.4]
  assign regs_44_io_enable = 1'h1; // @[RegFile.scala 74:20:@42510.4]
  assign regs_45_clock = clock; // @[:@42519.4]
  assign regs_45_reset = io_reset; // @[:@42520.4 RegFile.scala 76:16:@42527.4]
  assign regs_45_io_in = 64'h0; // @[RegFile.scala 75:16:@42526.4]
  assign regs_45_io_reset = reset; // @[RegFile.scala 78:19:@42530.4]
  assign regs_45_io_enable = 1'h1; // @[RegFile.scala 74:20:@42524.4]
  assign regs_46_clock = clock; // @[:@42533.4]
  assign regs_46_reset = io_reset; // @[:@42534.4 RegFile.scala 76:16:@42541.4]
  assign regs_46_io_in = 64'h0; // @[RegFile.scala 75:16:@42540.4]
  assign regs_46_io_reset = reset; // @[RegFile.scala 78:19:@42544.4]
  assign regs_46_io_enable = 1'h1; // @[RegFile.scala 74:20:@42538.4]
  assign regs_47_clock = clock; // @[:@42547.4]
  assign regs_47_reset = io_reset; // @[:@42548.4 RegFile.scala 76:16:@42555.4]
  assign regs_47_io_in = 64'h0; // @[RegFile.scala 75:16:@42554.4]
  assign regs_47_io_reset = reset; // @[RegFile.scala 78:19:@42558.4]
  assign regs_47_io_enable = 1'h1; // @[RegFile.scala 74:20:@42552.4]
  assign regs_48_clock = clock; // @[:@42561.4]
  assign regs_48_reset = io_reset; // @[:@42562.4 RegFile.scala 76:16:@42569.4]
  assign regs_48_io_in = 64'h0; // @[RegFile.scala 75:16:@42568.4]
  assign regs_48_io_reset = reset; // @[RegFile.scala 78:19:@42572.4]
  assign regs_48_io_enable = 1'h1; // @[RegFile.scala 74:20:@42566.4]
  assign regs_49_clock = clock; // @[:@42575.4]
  assign regs_49_reset = io_reset; // @[:@42576.4 RegFile.scala 76:16:@42583.4]
  assign regs_49_io_in = 64'h0; // @[RegFile.scala 75:16:@42582.4]
  assign regs_49_io_reset = reset; // @[RegFile.scala 78:19:@42586.4]
  assign regs_49_io_enable = 1'h1; // @[RegFile.scala 74:20:@42580.4]
  assign regs_50_clock = clock; // @[:@42589.4]
  assign regs_50_reset = io_reset; // @[:@42590.4 RegFile.scala 76:16:@42597.4]
  assign regs_50_io_in = 64'h0; // @[RegFile.scala 75:16:@42596.4]
  assign regs_50_io_reset = reset; // @[RegFile.scala 78:19:@42600.4]
  assign regs_50_io_enable = 1'h1; // @[RegFile.scala 74:20:@42594.4]
  assign regs_51_clock = clock; // @[:@42603.4]
  assign regs_51_reset = io_reset; // @[:@42604.4 RegFile.scala 76:16:@42611.4]
  assign regs_51_io_in = 64'h0; // @[RegFile.scala 75:16:@42610.4]
  assign regs_51_io_reset = reset; // @[RegFile.scala 78:19:@42614.4]
  assign regs_51_io_enable = 1'h1; // @[RegFile.scala 74:20:@42608.4]
  assign regs_52_clock = clock; // @[:@42617.4]
  assign regs_52_reset = io_reset; // @[:@42618.4 RegFile.scala 76:16:@42625.4]
  assign regs_52_io_in = 64'h0; // @[RegFile.scala 75:16:@42624.4]
  assign regs_52_io_reset = reset; // @[RegFile.scala 78:19:@42628.4]
  assign regs_52_io_enable = 1'h1; // @[RegFile.scala 74:20:@42622.4]
  assign regs_53_clock = clock; // @[:@42631.4]
  assign regs_53_reset = io_reset; // @[:@42632.4 RegFile.scala 76:16:@42639.4]
  assign regs_53_io_in = 64'h0; // @[RegFile.scala 75:16:@42638.4]
  assign regs_53_io_reset = reset; // @[RegFile.scala 78:19:@42642.4]
  assign regs_53_io_enable = 1'h1; // @[RegFile.scala 74:20:@42636.4]
  assign regs_54_clock = clock; // @[:@42645.4]
  assign regs_54_reset = io_reset; // @[:@42646.4 RegFile.scala 76:16:@42653.4]
  assign regs_54_io_in = 64'h0; // @[RegFile.scala 75:16:@42652.4]
  assign regs_54_io_reset = reset; // @[RegFile.scala 78:19:@42656.4]
  assign regs_54_io_enable = 1'h1; // @[RegFile.scala 74:20:@42650.4]
  assign regs_55_clock = clock; // @[:@42659.4]
  assign regs_55_reset = io_reset; // @[:@42660.4 RegFile.scala 76:16:@42667.4]
  assign regs_55_io_in = 64'h0; // @[RegFile.scala 75:16:@42666.4]
  assign regs_55_io_reset = reset; // @[RegFile.scala 78:19:@42670.4]
  assign regs_55_io_enable = 1'h1; // @[RegFile.scala 74:20:@42664.4]
  assign regs_56_clock = clock; // @[:@42673.4]
  assign regs_56_reset = io_reset; // @[:@42674.4 RegFile.scala 76:16:@42681.4]
  assign regs_56_io_in = 64'h0; // @[RegFile.scala 75:16:@42680.4]
  assign regs_56_io_reset = reset; // @[RegFile.scala 78:19:@42684.4]
  assign regs_56_io_enable = 1'h1; // @[RegFile.scala 74:20:@42678.4]
  assign regs_57_clock = clock; // @[:@42687.4]
  assign regs_57_reset = io_reset; // @[:@42688.4 RegFile.scala 76:16:@42695.4]
  assign regs_57_io_in = 64'h0; // @[RegFile.scala 75:16:@42694.4]
  assign regs_57_io_reset = reset; // @[RegFile.scala 78:19:@42698.4]
  assign regs_57_io_enable = 1'h1; // @[RegFile.scala 74:20:@42692.4]
  assign regs_58_clock = clock; // @[:@42701.4]
  assign regs_58_reset = io_reset; // @[:@42702.4 RegFile.scala 76:16:@42709.4]
  assign regs_58_io_in = 64'h0; // @[RegFile.scala 75:16:@42708.4]
  assign regs_58_io_reset = reset; // @[RegFile.scala 78:19:@42712.4]
  assign regs_58_io_enable = 1'h1; // @[RegFile.scala 74:20:@42706.4]
  assign regs_59_clock = clock; // @[:@42715.4]
  assign regs_59_reset = io_reset; // @[:@42716.4 RegFile.scala 76:16:@42723.4]
  assign regs_59_io_in = 64'h0; // @[RegFile.scala 75:16:@42722.4]
  assign regs_59_io_reset = reset; // @[RegFile.scala 78:19:@42726.4]
  assign regs_59_io_enable = 1'h1; // @[RegFile.scala 74:20:@42720.4]
  assign regs_60_clock = clock; // @[:@42729.4]
  assign regs_60_reset = io_reset; // @[:@42730.4 RegFile.scala 76:16:@42737.4]
  assign regs_60_io_in = 64'h0; // @[RegFile.scala 75:16:@42736.4]
  assign regs_60_io_reset = reset; // @[RegFile.scala 78:19:@42740.4]
  assign regs_60_io_enable = 1'h1; // @[RegFile.scala 74:20:@42734.4]
  assign regs_61_clock = clock; // @[:@42743.4]
  assign regs_61_reset = io_reset; // @[:@42744.4 RegFile.scala 76:16:@42751.4]
  assign regs_61_io_in = 64'h0; // @[RegFile.scala 75:16:@42750.4]
  assign regs_61_io_reset = reset; // @[RegFile.scala 78:19:@42754.4]
  assign regs_61_io_enable = 1'h1; // @[RegFile.scala 74:20:@42748.4]
  assign regs_62_clock = clock; // @[:@42757.4]
  assign regs_62_reset = io_reset; // @[:@42758.4 RegFile.scala 76:16:@42765.4]
  assign regs_62_io_in = 64'h0; // @[RegFile.scala 75:16:@42764.4]
  assign regs_62_io_reset = reset; // @[RegFile.scala 78:19:@42768.4]
  assign regs_62_io_enable = 1'h1; // @[RegFile.scala 74:20:@42762.4]
  assign regs_63_clock = clock; // @[:@42771.4]
  assign regs_63_reset = io_reset; // @[:@42772.4 RegFile.scala 76:16:@42779.4]
  assign regs_63_io_in = 64'h0; // @[RegFile.scala 75:16:@42778.4]
  assign regs_63_io_reset = reset; // @[RegFile.scala 78:19:@42782.4]
  assign regs_63_io_enable = 1'h1; // @[RegFile.scala 74:20:@42776.4]
  assign regs_64_clock = clock; // @[:@42785.4]
  assign regs_64_reset = io_reset; // @[:@42786.4 RegFile.scala 76:16:@42793.4]
  assign regs_64_io_in = 64'h0; // @[RegFile.scala 75:16:@42792.4]
  assign regs_64_io_reset = reset; // @[RegFile.scala 78:19:@42796.4]
  assign regs_64_io_enable = 1'h1; // @[RegFile.scala 74:20:@42790.4]
  assign regs_65_clock = clock; // @[:@42799.4]
  assign regs_65_reset = io_reset; // @[:@42800.4 RegFile.scala 76:16:@42807.4]
  assign regs_65_io_in = 64'h0; // @[RegFile.scala 75:16:@42806.4]
  assign regs_65_io_reset = reset; // @[RegFile.scala 78:19:@42810.4]
  assign regs_65_io_enable = 1'h1; // @[RegFile.scala 74:20:@42804.4]
  assign regs_66_clock = clock; // @[:@42813.4]
  assign regs_66_reset = io_reset; // @[:@42814.4 RegFile.scala 76:16:@42821.4]
  assign regs_66_io_in = 64'h0; // @[RegFile.scala 75:16:@42820.4]
  assign regs_66_io_reset = reset; // @[RegFile.scala 78:19:@42824.4]
  assign regs_66_io_enable = 1'h1; // @[RegFile.scala 74:20:@42818.4]
  assign regs_67_clock = clock; // @[:@42827.4]
  assign regs_67_reset = io_reset; // @[:@42828.4 RegFile.scala 76:16:@42835.4]
  assign regs_67_io_in = 64'h0; // @[RegFile.scala 75:16:@42834.4]
  assign regs_67_io_reset = reset; // @[RegFile.scala 78:19:@42838.4]
  assign regs_67_io_enable = 1'h1; // @[RegFile.scala 74:20:@42832.4]
  assign regs_68_clock = clock; // @[:@42841.4]
  assign regs_68_reset = io_reset; // @[:@42842.4 RegFile.scala 76:16:@42849.4]
  assign regs_68_io_in = 64'h0; // @[RegFile.scala 75:16:@42848.4]
  assign regs_68_io_reset = reset; // @[RegFile.scala 78:19:@42852.4]
  assign regs_68_io_enable = 1'h1; // @[RegFile.scala 74:20:@42846.4]
  assign regs_69_clock = clock; // @[:@42855.4]
  assign regs_69_reset = io_reset; // @[:@42856.4 RegFile.scala 76:16:@42863.4]
  assign regs_69_io_in = 64'h0; // @[RegFile.scala 75:16:@42862.4]
  assign regs_69_io_reset = reset; // @[RegFile.scala 78:19:@42866.4]
  assign regs_69_io_enable = 1'h1; // @[RegFile.scala 74:20:@42860.4]
  assign regs_70_clock = clock; // @[:@42869.4]
  assign regs_70_reset = io_reset; // @[:@42870.4 RegFile.scala 76:16:@42877.4]
  assign regs_70_io_in = 64'h0; // @[RegFile.scala 75:16:@42876.4]
  assign regs_70_io_reset = reset; // @[RegFile.scala 78:19:@42880.4]
  assign regs_70_io_enable = 1'h1; // @[RegFile.scala 74:20:@42874.4]
  assign regs_71_clock = clock; // @[:@42883.4]
  assign regs_71_reset = io_reset; // @[:@42884.4 RegFile.scala 76:16:@42891.4]
  assign regs_71_io_in = 64'h0; // @[RegFile.scala 75:16:@42890.4]
  assign regs_71_io_reset = reset; // @[RegFile.scala 78:19:@42894.4]
  assign regs_71_io_enable = 1'h1; // @[RegFile.scala 74:20:@42888.4]
  assign regs_72_clock = clock; // @[:@42897.4]
  assign regs_72_reset = io_reset; // @[:@42898.4 RegFile.scala 76:16:@42905.4]
  assign regs_72_io_in = 64'h0; // @[RegFile.scala 75:16:@42904.4]
  assign regs_72_io_reset = reset; // @[RegFile.scala 78:19:@42908.4]
  assign regs_72_io_enable = 1'h1; // @[RegFile.scala 74:20:@42902.4]
  assign regs_73_clock = clock; // @[:@42911.4]
  assign regs_73_reset = io_reset; // @[:@42912.4 RegFile.scala 76:16:@42919.4]
  assign regs_73_io_in = 64'h0; // @[RegFile.scala 75:16:@42918.4]
  assign regs_73_io_reset = reset; // @[RegFile.scala 78:19:@42922.4]
  assign regs_73_io_enable = 1'h1; // @[RegFile.scala 74:20:@42916.4]
  assign regs_74_clock = clock; // @[:@42925.4]
  assign regs_74_reset = io_reset; // @[:@42926.4 RegFile.scala 76:16:@42933.4]
  assign regs_74_io_in = 64'h0; // @[RegFile.scala 75:16:@42932.4]
  assign regs_74_io_reset = reset; // @[RegFile.scala 78:19:@42936.4]
  assign regs_74_io_enable = 1'h1; // @[RegFile.scala 74:20:@42930.4]
  assign regs_75_clock = clock; // @[:@42939.4]
  assign regs_75_reset = io_reset; // @[:@42940.4 RegFile.scala 76:16:@42947.4]
  assign regs_75_io_in = 64'h0; // @[RegFile.scala 75:16:@42946.4]
  assign regs_75_io_reset = reset; // @[RegFile.scala 78:19:@42950.4]
  assign regs_75_io_enable = 1'h1; // @[RegFile.scala 74:20:@42944.4]
  assign regs_76_clock = clock; // @[:@42953.4]
  assign regs_76_reset = io_reset; // @[:@42954.4 RegFile.scala 76:16:@42961.4]
  assign regs_76_io_in = 64'h0; // @[RegFile.scala 75:16:@42960.4]
  assign regs_76_io_reset = reset; // @[RegFile.scala 78:19:@42964.4]
  assign regs_76_io_enable = 1'h1; // @[RegFile.scala 74:20:@42958.4]
  assign regs_77_clock = clock; // @[:@42967.4]
  assign regs_77_reset = io_reset; // @[:@42968.4 RegFile.scala 76:16:@42975.4]
  assign regs_77_io_in = 64'h0; // @[RegFile.scala 75:16:@42974.4]
  assign regs_77_io_reset = reset; // @[RegFile.scala 78:19:@42978.4]
  assign regs_77_io_enable = 1'h1; // @[RegFile.scala 74:20:@42972.4]
  assign regs_78_clock = clock; // @[:@42981.4]
  assign regs_78_reset = io_reset; // @[:@42982.4 RegFile.scala 76:16:@42989.4]
  assign regs_78_io_in = 64'h0; // @[RegFile.scala 75:16:@42988.4]
  assign regs_78_io_reset = reset; // @[RegFile.scala 78:19:@42992.4]
  assign regs_78_io_enable = 1'h1; // @[RegFile.scala 74:20:@42986.4]
  assign regs_79_clock = clock; // @[:@42995.4]
  assign regs_79_reset = io_reset; // @[:@42996.4 RegFile.scala 76:16:@43003.4]
  assign regs_79_io_in = 64'h0; // @[RegFile.scala 75:16:@43002.4]
  assign regs_79_io_reset = reset; // @[RegFile.scala 78:19:@43006.4]
  assign regs_79_io_enable = 1'h1; // @[RegFile.scala 74:20:@43000.4]
  assign regs_80_clock = clock; // @[:@43009.4]
  assign regs_80_reset = io_reset; // @[:@43010.4 RegFile.scala 76:16:@43017.4]
  assign regs_80_io_in = 64'h0; // @[RegFile.scala 75:16:@43016.4]
  assign regs_80_io_reset = reset; // @[RegFile.scala 78:19:@43020.4]
  assign regs_80_io_enable = 1'h1; // @[RegFile.scala 74:20:@43014.4]
  assign regs_81_clock = clock; // @[:@43023.4]
  assign regs_81_reset = io_reset; // @[:@43024.4 RegFile.scala 76:16:@43031.4]
  assign regs_81_io_in = 64'h0; // @[RegFile.scala 75:16:@43030.4]
  assign regs_81_io_reset = reset; // @[RegFile.scala 78:19:@43034.4]
  assign regs_81_io_enable = 1'h1; // @[RegFile.scala 74:20:@43028.4]
  assign regs_82_clock = clock; // @[:@43037.4]
  assign regs_82_reset = io_reset; // @[:@43038.4 RegFile.scala 76:16:@43045.4]
  assign regs_82_io_in = 64'h0; // @[RegFile.scala 75:16:@43044.4]
  assign regs_82_io_reset = reset; // @[RegFile.scala 78:19:@43048.4]
  assign regs_82_io_enable = 1'h1; // @[RegFile.scala 74:20:@43042.4]
  assign regs_83_clock = clock; // @[:@43051.4]
  assign regs_83_reset = io_reset; // @[:@43052.4 RegFile.scala 76:16:@43059.4]
  assign regs_83_io_in = 64'h0; // @[RegFile.scala 75:16:@43058.4]
  assign regs_83_io_reset = reset; // @[RegFile.scala 78:19:@43062.4]
  assign regs_83_io_enable = 1'h1; // @[RegFile.scala 74:20:@43056.4]
  assign regs_84_clock = clock; // @[:@43065.4]
  assign regs_84_reset = io_reset; // @[:@43066.4 RegFile.scala 76:16:@43073.4]
  assign regs_84_io_in = 64'h0; // @[RegFile.scala 75:16:@43072.4]
  assign regs_84_io_reset = reset; // @[RegFile.scala 78:19:@43076.4]
  assign regs_84_io_enable = 1'h1; // @[RegFile.scala 74:20:@43070.4]
  assign regs_85_clock = clock; // @[:@43079.4]
  assign regs_85_reset = io_reset; // @[:@43080.4 RegFile.scala 76:16:@43087.4]
  assign regs_85_io_in = 64'h0; // @[RegFile.scala 75:16:@43086.4]
  assign regs_85_io_reset = reset; // @[RegFile.scala 78:19:@43090.4]
  assign regs_85_io_enable = 1'h1; // @[RegFile.scala 74:20:@43084.4]
  assign regs_86_clock = clock; // @[:@43093.4]
  assign regs_86_reset = io_reset; // @[:@43094.4 RegFile.scala 76:16:@43101.4]
  assign regs_86_io_in = 64'h0; // @[RegFile.scala 75:16:@43100.4]
  assign regs_86_io_reset = reset; // @[RegFile.scala 78:19:@43104.4]
  assign regs_86_io_enable = 1'h1; // @[RegFile.scala 74:20:@43098.4]
  assign regs_87_clock = clock; // @[:@43107.4]
  assign regs_87_reset = io_reset; // @[:@43108.4 RegFile.scala 76:16:@43115.4]
  assign regs_87_io_in = 64'h0; // @[RegFile.scala 75:16:@43114.4]
  assign regs_87_io_reset = reset; // @[RegFile.scala 78:19:@43118.4]
  assign regs_87_io_enable = 1'h1; // @[RegFile.scala 74:20:@43112.4]
  assign regs_88_clock = clock; // @[:@43121.4]
  assign regs_88_reset = io_reset; // @[:@43122.4 RegFile.scala 76:16:@43129.4]
  assign regs_88_io_in = 64'h0; // @[RegFile.scala 75:16:@43128.4]
  assign regs_88_io_reset = reset; // @[RegFile.scala 78:19:@43132.4]
  assign regs_88_io_enable = 1'h1; // @[RegFile.scala 74:20:@43126.4]
  assign regs_89_clock = clock; // @[:@43135.4]
  assign regs_89_reset = io_reset; // @[:@43136.4 RegFile.scala 76:16:@43143.4]
  assign regs_89_io_in = 64'h0; // @[RegFile.scala 75:16:@43142.4]
  assign regs_89_io_reset = reset; // @[RegFile.scala 78:19:@43146.4]
  assign regs_89_io_enable = 1'h1; // @[RegFile.scala 74:20:@43140.4]
  assign regs_90_clock = clock; // @[:@43149.4]
  assign regs_90_reset = io_reset; // @[:@43150.4 RegFile.scala 76:16:@43157.4]
  assign regs_90_io_in = 64'h0; // @[RegFile.scala 75:16:@43156.4]
  assign regs_90_io_reset = reset; // @[RegFile.scala 78:19:@43160.4]
  assign regs_90_io_enable = 1'h1; // @[RegFile.scala 74:20:@43154.4]
  assign regs_91_clock = clock; // @[:@43163.4]
  assign regs_91_reset = io_reset; // @[:@43164.4 RegFile.scala 76:16:@43171.4]
  assign regs_91_io_in = 64'h0; // @[RegFile.scala 75:16:@43170.4]
  assign regs_91_io_reset = reset; // @[RegFile.scala 78:19:@43174.4]
  assign regs_91_io_enable = 1'h1; // @[RegFile.scala 74:20:@43168.4]
  assign regs_92_clock = clock; // @[:@43177.4]
  assign regs_92_reset = io_reset; // @[:@43178.4 RegFile.scala 76:16:@43185.4]
  assign regs_92_io_in = 64'h0; // @[RegFile.scala 75:16:@43184.4]
  assign regs_92_io_reset = reset; // @[RegFile.scala 78:19:@43188.4]
  assign regs_92_io_enable = 1'h1; // @[RegFile.scala 74:20:@43182.4]
  assign regs_93_clock = clock; // @[:@43191.4]
  assign regs_93_reset = io_reset; // @[:@43192.4 RegFile.scala 76:16:@43199.4]
  assign regs_93_io_in = 64'h0; // @[RegFile.scala 75:16:@43198.4]
  assign regs_93_io_reset = reset; // @[RegFile.scala 78:19:@43202.4]
  assign regs_93_io_enable = 1'h1; // @[RegFile.scala 74:20:@43196.4]
  assign regs_94_clock = clock; // @[:@43205.4]
  assign regs_94_reset = io_reset; // @[:@43206.4 RegFile.scala 76:16:@43213.4]
  assign regs_94_io_in = 64'h0; // @[RegFile.scala 75:16:@43212.4]
  assign regs_94_io_reset = reset; // @[RegFile.scala 78:19:@43216.4]
  assign regs_94_io_enable = 1'h1; // @[RegFile.scala 74:20:@43210.4]
  assign regs_95_clock = clock; // @[:@43219.4]
  assign regs_95_reset = io_reset; // @[:@43220.4 RegFile.scala 76:16:@43227.4]
  assign regs_95_io_in = 64'h0; // @[RegFile.scala 75:16:@43226.4]
  assign regs_95_io_reset = reset; // @[RegFile.scala 78:19:@43230.4]
  assign regs_95_io_enable = 1'h1; // @[RegFile.scala 74:20:@43224.4]
  assign regs_96_clock = clock; // @[:@43233.4]
  assign regs_96_reset = io_reset; // @[:@43234.4 RegFile.scala 76:16:@43241.4]
  assign regs_96_io_in = 64'h0; // @[RegFile.scala 75:16:@43240.4]
  assign regs_96_io_reset = reset; // @[RegFile.scala 78:19:@43244.4]
  assign regs_96_io_enable = 1'h1; // @[RegFile.scala 74:20:@43238.4]
  assign regs_97_clock = clock; // @[:@43247.4]
  assign regs_97_reset = io_reset; // @[:@43248.4 RegFile.scala 76:16:@43255.4]
  assign regs_97_io_in = 64'h0; // @[RegFile.scala 75:16:@43254.4]
  assign regs_97_io_reset = reset; // @[RegFile.scala 78:19:@43258.4]
  assign regs_97_io_enable = 1'h1; // @[RegFile.scala 74:20:@43252.4]
  assign regs_98_clock = clock; // @[:@43261.4]
  assign regs_98_reset = io_reset; // @[:@43262.4 RegFile.scala 76:16:@43269.4]
  assign regs_98_io_in = 64'h0; // @[RegFile.scala 75:16:@43268.4]
  assign regs_98_io_reset = reset; // @[RegFile.scala 78:19:@43272.4]
  assign regs_98_io_enable = 1'h1; // @[RegFile.scala 74:20:@43266.4]
  assign regs_99_clock = clock; // @[:@43275.4]
  assign regs_99_reset = io_reset; // @[:@43276.4 RegFile.scala 76:16:@43283.4]
  assign regs_99_io_in = 64'h0; // @[RegFile.scala 75:16:@43282.4]
  assign regs_99_io_reset = reset; // @[RegFile.scala 78:19:@43286.4]
  assign regs_99_io_enable = 1'h1; // @[RegFile.scala 74:20:@43280.4]
  assign regs_100_clock = clock; // @[:@43289.4]
  assign regs_100_reset = io_reset; // @[:@43290.4 RegFile.scala 76:16:@43297.4]
  assign regs_100_io_in = 64'h0; // @[RegFile.scala 75:16:@43296.4]
  assign regs_100_io_reset = reset; // @[RegFile.scala 78:19:@43300.4]
  assign regs_100_io_enable = 1'h1; // @[RegFile.scala 74:20:@43294.4]
  assign regs_101_clock = clock; // @[:@43303.4]
  assign regs_101_reset = io_reset; // @[:@43304.4 RegFile.scala 76:16:@43311.4]
  assign regs_101_io_in = 64'h0; // @[RegFile.scala 75:16:@43310.4]
  assign regs_101_io_reset = reset; // @[RegFile.scala 78:19:@43314.4]
  assign regs_101_io_enable = 1'h1; // @[RegFile.scala 74:20:@43308.4]
  assign regs_102_clock = clock; // @[:@43317.4]
  assign regs_102_reset = io_reset; // @[:@43318.4 RegFile.scala 76:16:@43325.4]
  assign regs_102_io_in = 64'h0; // @[RegFile.scala 75:16:@43324.4]
  assign regs_102_io_reset = reset; // @[RegFile.scala 78:19:@43328.4]
  assign regs_102_io_enable = 1'h1; // @[RegFile.scala 74:20:@43322.4]
  assign regs_103_clock = clock; // @[:@43331.4]
  assign regs_103_reset = io_reset; // @[:@43332.4 RegFile.scala 76:16:@43339.4]
  assign regs_103_io_in = 64'h0; // @[RegFile.scala 75:16:@43338.4]
  assign regs_103_io_reset = reset; // @[RegFile.scala 78:19:@43342.4]
  assign regs_103_io_enable = 1'h1; // @[RegFile.scala 74:20:@43336.4]
  assign regs_104_clock = clock; // @[:@43345.4]
  assign regs_104_reset = io_reset; // @[:@43346.4 RegFile.scala 76:16:@43353.4]
  assign regs_104_io_in = 64'h0; // @[RegFile.scala 75:16:@43352.4]
  assign regs_104_io_reset = reset; // @[RegFile.scala 78:19:@43356.4]
  assign regs_104_io_enable = 1'h1; // @[RegFile.scala 74:20:@43350.4]
  assign regs_105_clock = clock; // @[:@43359.4]
  assign regs_105_reset = io_reset; // @[:@43360.4 RegFile.scala 76:16:@43367.4]
  assign regs_105_io_in = 64'h0; // @[RegFile.scala 75:16:@43366.4]
  assign regs_105_io_reset = reset; // @[RegFile.scala 78:19:@43370.4]
  assign regs_105_io_enable = 1'h1; // @[RegFile.scala 74:20:@43364.4]
  assign regs_106_clock = clock; // @[:@43373.4]
  assign regs_106_reset = io_reset; // @[:@43374.4 RegFile.scala 76:16:@43381.4]
  assign regs_106_io_in = 64'h0; // @[RegFile.scala 75:16:@43380.4]
  assign regs_106_io_reset = reset; // @[RegFile.scala 78:19:@43384.4]
  assign regs_106_io_enable = 1'h1; // @[RegFile.scala 74:20:@43378.4]
  assign regs_107_clock = clock; // @[:@43387.4]
  assign regs_107_reset = io_reset; // @[:@43388.4 RegFile.scala 76:16:@43395.4]
  assign regs_107_io_in = 64'h0; // @[RegFile.scala 75:16:@43394.4]
  assign regs_107_io_reset = reset; // @[RegFile.scala 78:19:@43398.4]
  assign regs_107_io_enable = 1'h1; // @[RegFile.scala 74:20:@43392.4]
  assign regs_108_clock = clock; // @[:@43401.4]
  assign regs_108_reset = io_reset; // @[:@43402.4 RegFile.scala 76:16:@43409.4]
  assign regs_108_io_in = 64'h0; // @[RegFile.scala 75:16:@43408.4]
  assign regs_108_io_reset = reset; // @[RegFile.scala 78:19:@43412.4]
  assign regs_108_io_enable = 1'h1; // @[RegFile.scala 74:20:@43406.4]
  assign regs_109_clock = clock; // @[:@43415.4]
  assign regs_109_reset = io_reset; // @[:@43416.4 RegFile.scala 76:16:@43423.4]
  assign regs_109_io_in = 64'h0; // @[RegFile.scala 75:16:@43422.4]
  assign regs_109_io_reset = reset; // @[RegFile.scala 78:19:@43426.4]
  assign regs_109_io_enable = 1'h1; // @[RegFile.scala 74:20:@43420.4]
  assign regs_110_clock = clock; // @[:@43429.4]
  assign regs_110_reset = io_reset; // @[:@43430.4 RegFile.scala 76:16:@43437.4]
  assign regs_110_io_in = 64'h0; // @[RegFile.scala 75:16:@43436.4]
  assign regs_110_io_reset = reset; // @[RegFile.scala 78:19:@43440.4]
  assign regs_110_io_enable = 1'h1; // @[RegFile.scala 74:20:@43434.4]
  assign regs_111_clock = clock; // @[:@43443.4]
  assign regs_111_reset = io_reset; // @[:@43444.4 RegFile.scala 76:16:@43451.4]
  assign regs_111_io_in = 64'h0; // @[RegFile.scala 75:16:@43450.4]
  assign regs_111_io_reset = reset; // @[RegFile.scala 78:19:@43454.4]
  assign regs_111_io_enable = 1'h1; // @[RegFile.scala 74:20:@43448.4]
  assign regs_112_clock = clock; // @[:@43457.4]
  assign regs_112_reset = io_reset; // @[:@43458.4 RegFile.scala 76:16:@43465.4]
  assign regs_112_io_in = 64'h0; // @[RegFile.scala 75:16:@43464.4]
  assign regs_112_io_reset = reset; // @[RegFile.scala 78:19:@43468.4]
  assign regs_112_io_enable = 1'h1; // @[RegFile.scala 74:20:@43462.4]
  assign regs_113_clock = clock; // @[:@43471.4]
  assign regs_113_reset = io_reset; // @[:@43472.4 RegFile.scala 76:16:@43479.4]
  assign regs_113_io_in = 64'h0; // @[RegFile.scala 75:16:@43478.4]
  assign regs_113_io_reset = reset; // @[RegFile.scala 78:19:@43482.4]
  assign regs_113_io_enable = 1'h1; // @[RegFile.scala 74:20:@43476.4]
  assign regs_114_clock = clock; // @[:@43485.4]
  assign regs_114_reset = io_reset; // @[:@43486.4 RegFile.scala 76:16:@43493.4]
  assign regs_114_io_in = 64'h0; // @[RegFile.scala 75:16:@43492.4]
  assign regs_114_io_reset = reset; // @[RegFile.scala 78:19:@43496.4]
  assign regs_114_io_enable = 1'h1; // @[RegFile.scala 74:20:@43490.4]
  assign regs_115_clock = clock; // @[:@43499.4]
  assign regs_115_reset = io_reset; // @[:@43500.4 RegFile.scala 76:16:@43507.4]
  assign regs_115_io_in = 64'h0; // @[RegFile.scala 75:16:@43506.4]
  assign regs_115_io_reset = reset; // @[RegFile.scala 78:19:@43510.4]
  assign regs_115_io_enable = 1'h1; // @[RegFile.scala 74:20:@43504.4]
  assign regs_116_clock = clock; // @[:@43513.4]
  assign regs_116_reset = io_reset; // @[:@43514.4 RegFile.scala 76:16:@43521.4]
  assign regs_116_io_in = 64'h0; // @[RegFile.scala 75:16:@43520.4]
  assign regs_116_io_reset = reset; // @[RegFile.scala 78:19:@43524.4]
  assign regs_116_io_enable = 1'h1; // @[RegFile.scala 74:20:@43518.4]
  assign regs_117_clock = clock; // @[:@43527.4]
  assign regs_117_reset = io_reset; // @[:@43528.4 RegFile.scala 76:16:@43535.4]
  assign regs_117_io_in = 64'h0; // @[RegFile.scala 75:16:@43534.4]
  assign regs_117_io_reset = reset; // @[RegFile.scala 78:19:@43538.4]
  assign regs_117_io_enable = 1'h1; // @[RegFile.scala 74:20:@43532.4]
  assign regs_118_clock = clock; // @[:@43541.4]
  assign regs_118_reset = io_reset; // @[:@43542.4 RegFile.scala 76:16:@43549.4]
  assign regs_118_io_in = 64'h0; // @[RegFile.scala 75:16:@43548.4]
  assign regs_118_io_reset = reset; // @[RegFile.scala 78:19:@43552.4]
  assign regs_118_io_enable = 1'h1; // @[RegFile.scala 74:20:@43546.4]
  assign regs_119_clock = clock; // @[:@43555.4]
  assign regs_119_reset = io_reset; // @[:@43556.4 RegFile.scala 76:16:@43563.4]
  assign regs_119_io_in = 64'h0; // @[RegFile.scala 75:16:@43562.4]
  assign regs_119_io_reset = reset; // @[RegFile.scala 78:19:@43566.4]
  assign regs_119_io_enable = 1'h1; // @[RegFile.scala 74:20:@43560.4]
  assign regs_120_clock = clock; // @[:@43569.4]
  assign regs_120_reset = io_reset; // @[:@43570.4 RegFile.scala 76:16:@43577.4]
  assign regs_120_io_in = 64'h0; // @[RegFile.scala 75:16:@43576.4]
  assign regs_120_io_reset = reset; // @[RegFile.scala 78:19:@43580.4]
  assign regs_120_io_enable = 1'h1; // @[RegFile.scala 74:20:@43574.4]
  assign regs_121_clock = clock; // @[:@43583.4]
  assign regs_121_reset = io_reset; // @[:@43584.4 RegFile.scala 76:16:@43591.4]
  assign regs_121_io_in = 64'h0; // @[RegFile.scala 75:16:@43590.4]
  assign regs_121_io_reset = reset; // @[RegFile.scala 78:19:@43594.4]
  assign regs_121_io_enable = 1'h1; // @[RegFile.scala 74:20:@43588.4]
  assign regs_122_clock = clock; // @[:@43597.4]
  assign regs_122_reset = io_reset; // @[:@43598.4 RegFile.scala 76:16:@43605.4]
  assign regs_122_io_in = 64'h0; // @[RegFile.scala 75:16:@43604.4]
  assign regs_122_io_reset = reset; // @[RegFile.scala 78:19:@43608.4]
  assign regs_122_io_enable = 1'h1; // @[RegFile.scala 74:20:@43602.4]
  assign regs_123_clock = clock; // @[:@43611.4]
  assign regs_123_reset = io_reset; // @[:@43612.4 RegFile.scala 76:16:@43619.4]
  assign regs_123_io_in = 64'h0; // @[RegFile.scala 75:16:@43618.4]
  assign regs_123_io_reset = reset; // @[RegFile.scala 78:19:@43622.4]
  assign regs_123_io_enable = 1'h1; // @[RegFile.scala 74:20:@43616.4]
  assign regs_124_clock = clock; // @[:@43625.4]
  assign regs_124_reset = io_reset; // @[:@43626.4 RegFile.scala 76:16:@43633.4]
  assign regs_124_io_in = 64'h0; // @[RegFile.scala 75:16:@43632.4]
  assign regs_124_io_reset = reset; // @[RegFile.scala 78:19:@43636.4]
  assign regs_124_io_enable = 1'h1; // @[RegFile.scala 74:20:@43630.4]
  assign regs_125_clock = clock; // @[:@43639.4]
  assign regs_125_reset = io_reset; // @[:@43640.4 RegFile.scala 76:16:@43647.4]
  assign regs_125_io_in = 64'h0; // @[RegFile.scala 75:16:@43646.4]
  assign regs_125_io_reset = reset; // @[RegFile.scala 78:19:@43650.4]
  assign regs_125_io_enable = 1'h1; // @[RegFile.scala 74:20:@43644.4]
  assign regs_126_clock = clock; // @[:@43653.4]
  assign regs_126_reset = io_reset; // @[:@43654.4 RegFile.scala 76:16:@43661.4]
  assign regs_126_io_in = 64'h0; // @[RegFile.scala 75:16:@43660.4]
  assign regs_126_io_reset = reset; // @[RegFile.scala 78:19:@43664.4]
  assign regs_126_io_enable = 1'h1; // @[RegFile.scala 74:20:@43658.4]
  assign regs_127_clock = clock; // @[:@43667.4]
  assign regs_127_reset = io_reset; // @[:@43668.4 RegFile.scala 76:16:@43675.4]
  assign regs_127_io_in = 64'h0; // @[RegFile.scala 75:16:@43674.4]
  assign regs_127_io_reset = reset; // @[RegFile.scala 78:19:@43678.4]
  assign regs_127_io_enable = 1'h1; // @[RegFile.scala 74:20:@43672.4]
  assign regs_128_clock = clock; // @[:@43681.4]
  assign regs_128_reset = io_reset; // @[:@43682.4 RegFile.scala 76:16:@43689.4]
  assign regs_128_io_in = 64'h0; // @[RegFile.scala 75:16:@43688.4]
  assign regs_128_io_reset = reset; // @[RegFile.scala 78:19:@43692.4]
  assign regs_128_io_enable = 1'h1; // @[RegFile.scala 74:20:@43686.4]
  assign regs_129_clock = clock; // @[:@43695.4]
  assign regs_129_reset = io_reset; // @[:@43696.4 RegFile.scala 76:16:@43703.4]
  assign regs_129_io_in = 64'h0; // @[RegFile.scala 75:16:@43702.4]
  assign regs_129_io_reset = reset; // @[RegFile.scala 78:19:@43706.4]
  assign regs_129_io_enable = 1'h1; // @[RegFile.scala 74:20:@43700.4]
  assign regs_130_clock = clock; // @[:@43709.4]
  assign regs_130_reset = io_reset; // @[:@43710.4 RegFile.scala 76:16:@43717.4]
  assign regs_130_io_in = 64'h0; // @[RegFile.scala 75:16:@43716.4]
  assign regs_130_io_reset = reset; // @[RegFile.scala 78:19:@43720.4]
  assign regs_130_io_enable = 1'h1; // @[RegFile.scala 74:20:@43714.4]
  assign regs_131_clock = clock; // @[:@43723.4]
  assign regs_131_reset = io_reset; // @[:@43724.4 RegFile.scala 76:16:@43731.4]
  assign regs_131_io_in = 64'h0; // @[RegFile.scala 75:16:@43730.4]
  assign regs_131_io_reset = reset; // @[RegFile.scala 78:19:@43734.4]
  assign regs_131_io_enable = 1'h1; // @[RegFile.scala 74:20:@43728.4]
  assign regs_132_clock = clock; // @[:@43737.4]
  assign regs_132_reset = io_reset; // @[:@43738.4 RegFile.scala 76:16:@43745.4]
  assign regs_132_io_in = 64'h0; // @[RegFile.scala 75:16:@43744.4]
  assign regs_132_io_reset = reset; // @[RegFile.scala 78:19:@43748.4]
  assign regs_132_io_enable = 1'h1; // @[RegFile.scala 74:20:@43742.4]
  assign regs_133_clock = clock; // @[:@43751.4]
  assign regs_133_reset = io_reset; // @[:@43752.4 RegFile.scala 76:16:@43759.4]
  assign regs_133_io_in = 64'h0; // @[RegFile.scala 75:16:@43758.4]
  assign regs_133_io_reset = reset; // @[RegFile.scala 78:19:@43762.4]
  assign regs_133_io_enable = 1'h1; // @[RegFile.scala 74:20:@43756.4]
  assign regs_134_clock = clock; // @[:@43765.4]
  assign regs_134_reset = io_reset; // @[:@43766.4 RegFile.scala 76:16:@43773.4]
  assign regs_134_io_in = 64'h0; // @[RegFile.scala 75:16:@43772.4]
  assign regs_134_io_reset = reset; // @[RegFile.scala 78:19:@43776.4]
  assign regs_134_io_enable = 1'h1; // @[RegFile.scala 74:20:@43770.4]
  assign regs_135_clock = clock; // @[:@43779.4]
  assign regs_135_reset = io_reset; // @[:@43780.4 RegFile.scala 76:16:@43787.4]
  assign regs_135_io_in = 64'h0; // @[RegFile.scala 75:16:@43786.4]
  assign regs_135_io_reset = reset; // @[RegFile.scala 78:19:@43790.4]
  assign regs_135_io_enable = 1'h1; // @[RegFile.scala 74:20:@43784.4]
  assign regs_136_clock = clock; // @[:@43793.4]
  assign regs_136_reset = io_reset; // @[:@43794.4 RegFile.scala 76:16:@43801.4]
  assign regs_136_io_in = 64'h0; // @[RegFile.scala 75:16:@43800.4]
  assign regs_136_io_reset = reset; // @[RegFile.scala 78:19:@43804.4]
  assign regs_136_io_enable = 1'h1; // @[RegFile.scala 74:20:@43798.4]
  assign regs_137_clock = clock; // @[:@43807.4]
  assign regs_137_reset = io_reset; // @[:@43808.4 RegFile.scala 76:16:@43815.4]
  assign regs_137_io_in = 64'h0; // @[RegFile.scala 75:16:@43814.4]
  assign regs_137_io_reset = reset; // @[RegFile.scala 78:19:@43818.4]
  assign regs_137_io_enable = 1'h1; // @[RegFile.scala 74:20:@43812.4]
  assign regs_138_clock = clock; // @[:@43821.4]
  assign regs_138_reset = io_reset; // @[:@43822.4 RegFile.scala 76:16:@43829.4]
  assign regs_138_io_in = 64'h0; // @[RegFile.scala 75:16:@43828.4]
  assign regs_138_io_reset = reset; // @[RegFile.scala 78:19:@43832.4]
  assign regs_138_io_enable = 1'h1; // @[RegFile.scala 74:20:@43826.4]
  assign regs_139_clock = clock; // @[:@43835.4]
  assign regs_139_reset = io_reset; // @[:@43836.4 RegFile.scala 76:16:@43843.4]
  assign regs_139_io_in = 64'h0; // @[RegFile.scala 75:16:@43842.4]
  assign regs_139_io_reset = reset; // @[RegFile.scala 78:19:@43846.4]
  assign regs_139_io_enable = 1'h1; // @[RegFile.scala 74:20:@43840.4]
  assign regs_140_clock = clock; // @[:@43849.4]
  assign regs_140_reset = io_reset; // @[:@43850.4 RegFile.scala 76:16:@43857.4]
  assign regs_140_io_in = 64'h0; // @[RegFile.scala 75:16:@43856.4]
  assign regs_140_io_reset = reset; // @[RegFile.scala 78:19:@43860.4]
  assign regs_140_io_enable = 1'h1; // @[RegFile.scala 74:20:@43854.4]
  assign regs_141_clock = clock; // @[:@43863.4]
  assign regs_141_reset = io_reset; // @[:@43864.4 RegFile.scala 76:16:@43871.4]
  assign regs_141_io_in = 64'h0; // @[RegFile.scala 75:16:@43870.4]
  assign regs_141_io_reset = reset; // @[RegFile.scala 78:19:@43874.4]
  assign regs_141_io_enable = 1'h1; // @[RegFile.scala 74:20:@43868.4]
  assign regs_142_clock = clock; // @[:@43877.4]
  assign regs_142_reset = io_reset; // @[:@43878.4 RegFile.scala 76:16:@43885.4]
  assign regs_142_io_in = 64'h0; // @[RegFile.scala 75:16:@43884.4]
  assign regs_142_io_reset = reset; // @[RegFile.scala 78:19:@43888.4]
  assign regs_142_io_enable = 1'h1; // @[RegFile.scala 74:20:@43882.4]
  assign regs_143_clock = clock; // @[:@43891.4]
  assign regs_143_reset = io_reset; // @[:@43892.4 RegFile.scala 76:16:@43899.4]
  assign regs_143_io_in = 64'h0; // @[RegFile.scala 75:16:@43898.4]
  assign regs_143_io_reset = reset; // @[RegFile.scala 78:19:@43902.4]
  assign regs_143_io_enable = 1'h1; // @[RegFile.scala 74:20:@43896.4]
  assign regs_144_clock = clock; // @[:@43905.4]
  assign regs_144_reset = io_reset; // @[:@43906.4 RegFile.scala 76:16:@43913.4]
  assign regs_144_io_in = 64'h0; // @[RegFile.scala 75:16:@43912.4]
  assign regs_144_io_reset = reset; // @[RegFile.scala 78:19:@43916.4]
  assign regs_144_io_enable = 1'h1; // @[RegFile.scala 74:20:@43910.4]
  assign regs_145_clock = clock; // @[:@43919.4]
  assign regs_145_reset = io_reset; // @[:@43920.4 RegFile.scala 76:16:@43927.4]
  assign regs_145_io_in = 64'h0; // @[RegFile.scala 75:16:@43926.4]
  assign regs_145_io_reset = reset; // @[RegFile.scala 78:19:@43930.4]
  assign regs_145_io_enable = 1'h1; // @[RegFile.scala 74:20:@43924.4]
  assign regs_146_clock = clock; // @[:@43933.4]
  assign regs_146_reset = io_reset; // @[:@43934.4 RegFile.scala 76:16:@43941.4]
  assign regs_146_io_in = 64'h0; // @[RegFile.scala 75:16:@43940.4]
  assign regs_146_io_reset = reset; // @[RegFile.scala 78:19:@43944.4]
  assign regs_146_io_enable = 1'h1; // @[RegFile.scala 74:20:@43938.4]
  assign regs_147_clock = clock; // @[:@43947.4]
  assign regs_147_reset = io_reset; // @[:@43948.4 RegFile.scala 76:16:@43955.4]
  assign regs_147_io_in = 64'h0; // @[RegFile.scala 75:16:@43954.4]
  assign regs_147_io_reset = reset; // @[RegFile.scala 78:19:@43958.4]
  assign regs_147_io_enable = 1'h1; // @[RegFile.scala 74:20:@43952.4]
  assign regs_148_clock = clock; // @[:@43961.4]
  assign regs_148_reset = io_reset; // @[:@43962.4 RegFile.scala 76:16:@43969.4]
  assign regs_148_io_in = 64'h0; // @[RegFile.scala 75:16:@43968.4]
  assign regs_148_io_reset = reset; // @[RegFile.scala 78:19:@43972.4]
  assign regs_148_io_enable = 1'h1; // @[RegFile.scala 74:20:@43966.4]
  assign regs_149_clock = clock; // @[:@43975.4]
  assign regs_149_reset = io_reset; // @[:@43976.4 RegFile.scala 76:16:@43983.4]
  assign regs_149_io_in = 64'h0; // @[RegFile.scala 75:16:@43982.4]
  assign regs_149_io_reset = reset; // @[RegFile.scala 78:19:@43986.4]
  assign regs_149_io_enable = 1'h1; // @[RegFile.scala 74:20:@43980.4]
  assign regs_150_clock = clock; // @[:@43989.4]
  assign regs_150_reset = io_reset; // @[:@43990.4 RegFile.scala 76:16:@43997.4]
  assign regs_150_io_in = 64'h0; // @[RegFile.scala 75:16:@43996.4]
  assign regs_150_io_reset = reset; // @[RegFile.scala 78:19:@44000.4]
  assign regs_150_io_enable = 1'h1; // @[RegFile.scala 74:20:@43994.4]
  assign regs_151_clock = clock; // @[:@44003.4]
  assign regs_151_reset = io_reset; // @[:@44004.4 RegFile.scala 76:16:@44011.4]
  assign regs_151_io_in = 64'h0; // @[RegFile.scala 75:16:@44010.4]
  assign regs_151_io_reset = reset; // @[RegFile.scala 78:19:@44014.4]
  assign regs_151_io_enable = 1'h1; // @[RegFile.scala 74:20:@44008.4]
  assign regs_152_clock = clock; // @[:@44017.4]
  assign regs_152_reset = io_reset; // @[:@44018.4 RegFile.scala 76:16:@44025.4]
  assign regs_152_io_in = 64'h0; // @[RegFile.scala 75:16:@44024.4]
  assign regs_152_io_reset = reset; // @[RegFile.scala 78:19:@44028.4]
  assign regs_152_io_enable = 1'h1; // @[RegFile.scala 74:20:@44022.4]
  assign regs_153_clock = clock; // @[:@44031.4]
  assign regs_153_reset = io_reset; // @[:@44032.4 RegFile.scala 76:16:@44039.4]
  assign regs_153_io_in = 64'h0; // @[RegFile.scala 75:16:@44038.4]
  assign regs_153_io_reset = reset; // @[RegFile.scala 78:19:@44042.4]
  assign regs_153_io_enable = 1'h1; // @[RegFile.scala 74:20:@44036.4]
  assign regs_154_clock = clock; // @[:@44045.4]
  assign regs_154_reset = io_reset; // @[:@44046.4 RegFile.scala 76:16:@44053.4]
  assign regs_154_io_in = 64'h0; // @[RegFile.scala 75:16:@44052.4]
  assign regs_154_io_reset = reset; // @[RegFile.scala 78:19:@44056.4]
  assign regs_154_io_enable = 1'h1; // @[RegFile.scala 74:20:@44050.4]
  assign regs_155_clock = clock; // @[:@44059.4]
  assign regs_155_reset = io_reset; // @[:@44060.4 RegFile.scala 76:16:@44067.4]
  assign regs_155_io_in = 64'h0; // @[RegFile.scala 75:16:@44066.4]
  assign regs_155_io_reset = reset; // @[RegFile.scala 78:19:@44070.4]
  assign regs_155_io_enable = 1'h1; // @[RegFile.scala 74:20:@44064.4]
  assign regs_156_clock = clock; // @[:@44073.4]
  assign regs_156_reset = io_reset; // @[:@44074.4 RegFile.scala 76:16:@44081.4]
  assign regs_156_io_in = 64'h0; // @[RegFile.scala 75:16:@44080.4]
  assign regs_156_io_reset = reset; // @[RegFile.scala 78:19:@44084.4]
  assign regs_156_io_enable = 1'h1; // @[RegFile.scala 74:20:@44078.4]
  assign regs_157_clock = clock; // @[:@44087.4]
  assign regs_157_reset = io_reset; // @[:@44088.4 RegFile.scala 76:16:@44095.4]
  assign regs_157_io_in = 64'h0; // @[RegFile.scala 75:16:@44094.4]
  assign regs_157_io_reset = reset; // @[RegFile.scala 78:19:@44098.4]
  assign regs_157_io_enable = 1'h1; // @[RegFile.scala 74:20:@44092.4]
  assign regs_158_clock = clock; // @[:@44101.4]
  assign regs_158_reset = io_reset; // @[:@44102.4 RegFile.scala 76:16:@44109.4]
  assign regs_158_io_in = 64'h0; // @[RegFile.scala 75:16:@44108.4]
  assign regs_158_io_reset = reset; // @[RegFile.scala 78:19:@44112.4]
  assign regs_158_io_enable = 1'h1; // @[RegFile.scala 74:20:@44106.4]
  assign regs_159_clock = clock; // @[:@44115.4]
  assign regs_159_reset = io_reset; // @[:@44116.4 RegFile.scala 76:16:@44123.4]
  assign regs_159_io_in = 64'h0; // @[RegFile.scala 75:16:@44122.4]
  assign regs_159_io_reset = reset; // @[RegFile.scala 78:19:@44126.4]
  assign regs_159_io_enable = 1'h1; // @[RegFile.scala 74:20:@44120.4]
  assign regs_160_clock = clock; // @[:@44129.4]
  assign regs_160_reset = io_reset; // @[:@44130.4 RegFile.scala 76:16:@44137.4]
  assign regs_160_io_in = 64'h0; // @[RegFile.scala 75:16:@44136.4]
  assign regs_160_io_reset = reset; // @[RegFile.scala 78:19:@44140.4]
  assign regs_160_io_enable = 1'h1; // @[RegFile.scala 74:20:@44134.4]
  assign regs_161_clock = clock; // @[:@44143.4]
  assign regs_161_reset = io_reset; // @[:@44144.4 RegFile.scala 76:16:@44151.4]
  assign regs_161_io_in = 64'h0; // @[RegFile.scala 75:16:@44150.4]
  assign regs_161_io_reset = reset; // @[RegFile.scala 78:19:@44154.4]
  assign regs_161_io_enable = 1'h1; // @[RegFile.scala 74:20:@44148.4]
  assign regs_162_clock = clock; // @[:@44157.4]
  assign regs_162_reset = io_reset; // @[:@44158.4 RegFile.scala 76:16:@44165.4]
  assign regs_162_io_in = 64'h0; // @[RegFile.scala 75:16:@44164.4]
  assign regs_162_io_reset = reset; // @[RegFile.scala 78:19:@44168.4]
  assign regs_162_io_enable = 1'h1; // @[RegFile.scala 74:20:@44162.4]
  assign regs_163_clock = clock; // @[:@44171.4]
  assign regs_163_reset = io_reset; // @[:@44172.4 RegFile.scala 76:16:@44179.4]
  assign regs_163_io_in = 64'h0; // @[RegFile.scala 75:16:@44178.4]
  assign regs_163_io_reset = reset; // @[RegFile.scala 78:19:@44182.4]
  assign regs_163_io_enable = 1'h1; // @[RegFile.scala 74:20:@44176.4]
  assign regs_164_clock = clock; // @[:@44185.4]
  assign regs_164_reset = io_reset; // @[:@44186.4 RegFile.scala 76:16:@44193.4]
  assign regs_164_io_in = 64'h0; // @[RegFile.scala 75:16:@44192.4]
  assign regs_164_io_reset = reset; // @[RegFile.scala 78:19:@44196.4]
  assign regs_164_io_enable = 1'h1; // @[RegFile.scala 74:20:@44190.4]
  assign regs_165_clock = clock; // @[:@44199.4]
  assign regs_165_reset = io_reset; // @[:@44200.4 RegFile.scala 76:16:@44207.4]
  assign regs_165_io_in = 64'h0; // @[RegFile.scala 75:16:@44206.4]
  assign regs_165_io_reset = reset; // @[RegFile.scala 78:19:@44210.4]
  assign regs_165_io_enable = 1'h1; // @[RegFile.scala 74:20:@44204.4]
  assign regs_166_clock = clock; // @[:@44213.4]
  assign regs_166_reset = io_reset; // @[:@44214.4 RegFile.scala 76:16:@44221.4]
  assign regs_166_io_in = 64'h0; // @[RegFile.scala 75:16:@44220.4]
  assign regs_166_io_reset = reset; // @[RegFile.scala 78:19:@44224.4]
  assign regs_166_io_enable = 1'h1; // @[RegFile.scala 74:20:@44218.4]
  assign regs_167_clock = clock; // @[:@44227.4]
  assign regs_167_reset = io_reset; // @[:@44228.4 RegFile.scala 76:16:@44235.4]
  assign regs_167_io_in = 64'h0; // @[RegFile.scala 75:16:@44234.4]
  assign regs_167_io_reset = reset; // @[RegFile.scala 78:19:@44238.4]
  assign regs_167_io_enable = 1'h1; // @[RegFile.scala 74:20:@44232.4]
  assign regs_168_clock = clock; // @[:@44241.4]
  assign regs_168_reset = io_reset; // @[:@44242.4 RegFile.scala 76:16:@44249.4]
  assign regs_168_io_in = 64'h0; // @[RegFile.scala 75:16:@44248.4]
  assign regs_168_io_reset = reset; // @[RegFile.scala 78:19:@44252.4]
  assign regs_168_io_enable = 1'h1; // @[RegFile.scala 74:20:@44246.4]
  assign regs_169_clock = clock; // @[:@44255.4]
  assign regs_169_reset = io_reset; // @[:@44256.4 RegFile.scala 76:16:@44263.4]
  assign regs_169_io_in = 64'h0; // @[RegFile.scala 75:16:@44262.4]
  assign regs_169_io_reset = reset; // @[RegFile.scala 78:19:@44266.4]
  assign regs_169_io_enable = 1'h1; // @[RegFile.scala 74:20:@44260.4]
  assign regs_170_clock = clock; // @[:@44269.4]
  assign regs_170_reset = io_reset; // @[:@44270.4 RegFile.scala 76:16:@44277.4]
  assign regs_170_io_in = 64'h0; // @[RegFile.scala 75:16:@44276.4]
  assign regs_170_io_reset = reset; // @[RegFile.scala 78:19:@44280.4]
  assign regs_170_io_enable = 1'h1; // @[RegFile.scala 74:20:@44274.4]
  assign regs_171_clock = clock; // @[:@44283.4]
  assign regs_171_reset = io_reset; // @[:@44284.4 RegFile.scala 76:16:@44291.4]
  assign regs_171_io_in = 64'h0; // @[RegFile.scala 75:16:@44290.4]
  assign regs_171_io_reset = reset; // @[RegFile.scala 78:19:@44294.4]
  assign regs_171_io_enable = 1'h1; // @[RegFile.scala 74:20:@44288.4]
  assign regs_172_clock = clock; // @[:@44297.4]
  assign regs_172_reset = io_reset; // @[:@44298.4 RegFile.scala 76:16:@44305.4]
  assign regs_172_io_in = 64'h0; // @[RegFile.scala 75:16:@44304.4]
  assign regs_172_io_reset = reset; // @[RegFile.scala 78:19:@44308.4]
  assign regs_172_io_enable = 1'h1; // @[RegFile.scala 74:20:@44302.4]
  assign regs_173_clock = clock; // @[:@44311.4]
  assign regs_173_reset = io_reset; // @[:@44312.4 RegFile.scala 76:16:@44319.4]
  assign regs_173_io_in = 64'h0; // @[RegFile.scala 75:16:@44318.4]
  assign regs_173_io_reset = reset; // @[RegFile.scala 78:19:@44322.4]
  assign regs_173_io_enable = 1'h1; // @[RegFile.scala 74:20:@44316.4]
  assign regs_174_clock = clock; // @[:@44325.4]
  assign regs_174_reset = io_reset; // @[:@44326.4 RegFile.scala 76:16:@44333.4]
  assign regs_174_io_in = 64'h0; // @[RegFile.scala 75:16:@44332.4]
  assign regs_174_io_reset = reset; // @[RegFile.scala 78:19:@44336.4]
  assign regs_174_io_enable = 1'h1; // @[RegFile.scala 74:20:@44330.4]
  assign regs_175_clock = clock; // @[:@44339.4]
  assign regs_175_reset = io_reset; // @[:@44340.4 RegFile.scala 76:16:@44347.4]
  assign regs_175_io_in = 64'h0; // @[RegFile.scala 75:16:@44346.4]
  assign regs_175_io_reset = reset; // @[RegFile.scala 78:19:@44350.4]
  assign regs_175_io_enable = 1'h1; // @[RegFile.scala 74:20:@44344.4]
  assign regs_176_clock = clock; // @[:@44353.4]
  assign regs_176_reset = io_reset; // @[:@44354.4 RegFile.scala 76:16:@44361.4]
  assign regs_176_io_in = 64'h0; // @[RegFile.scala 75:16:@44360.4]
  assign regs_176_io_reset = reset; // @[RegFile.scala 78:19:@44364.4]
  assign regs_176_io_enable = 1'h1; // @[RegFile.scala 74:20:@44358.4]
  assign regs_177_clock = clock; // @[:@44367.4]
  assign regs_177_reset = io_reset; // @[:@44368.4 RegFile.scala 76:16:@44375.4]
  assign regs_177_io_in = 64'h0; // @[RegFile.scala 75:16:@44374.4]
  assign regs_177_io_reset = reset; // @[RegFile.scala 78:19:@44378.4]
  assign regs_177_io_enable = 1'h1; // @[RegFile.scala 74:20:@44372.4]
  assign regs_178_clock = clock; // @[:@44381.4]
  assign regs_178_reset = io_reset; // @[:@44382.4 RegFile.scala 76:16:@44389.4]
  assign regs_178_io_in = 64'h0; // @[RegFile.scala 75:16:@44388.4]
  assign regs_178_io_reset = reset; // @[RegFile.scala 78:19:@44392.4]
  assign regs_178_io_enable = 1'h1; // @[RegFile.scala 74:20:@44386.4]
  assign regs_179_clock = clock; // @[:@44395.4]
  assign regs_179_reset = io_reset; // @[:@44396.4 RegFile.scala 76:16:@44403.4]
  assign regs_179_io_in = 64'h0; // @[RegFile.scala 75:16:@44402.4]
  assign regs_179_io_reset = reset; // @[RegFile.scala 78:19:@44406.4]
  assign regs_179_io_enable = 1'h1; // @[RegFile.scala 74:20:@44400.4]
  assign regs_180_clock = clock; // @[:@44409.4]
  assign regs_180_reset = io_reset; // @[:@44410.4 RegFile.scala 76:16:@44417.4]
  assign regs_180_io_in = 64'h0; // @[RegFile.scala 75:16:@44416.4]
  assign regs_180_io_reset = reset; // @[RegFile.scala 78:19:@44420.4]
  assign regs_180_io_enable = 1'h1; // @[RegFile.scala 74:20:@44414.4]
  assign regs_181_clock = clock; // @[:@44423.4]
  assign regs_181_reset = io_reset; // @[:@44424.4 RegFile.scala 76:16:@44431.4]
  assign regs_181_io_in = 64'h0; // @[RegFile.scala 75:16:@44430.4]
  assign regs_181_io_reset = reset; // @[RegFile.scala 78:19:@44434.4]
  assign regs_181_io_enable = 1'h1; // @[RegFile.scala 74:20:@44428.4]
  assign regs_182_clock = clock; // @[:@44437.4]
  assign regs_182_reset = io_reset; // @[:@44438.4 RegFile.scala 76:16:@44445.4]
  assign regs_182_io_in = 64'h0; // @[RegFile.scala 75:16:@44444.4]
  assign regs_182_io_reset = reset; // @[RegFile.scala 78:19:@44448.4]
  assign regs_182_io_enable = 1'h1; // @[RegFile.scala 74:20:@44442.4]
  assign regs_183_clock = clock; // @[:@44451.4]
  assign regs_183_reset = io_reset; // @[:@44452.4 RegFile.scala 76:16:@44459.4]
  assign regs_183_io_in = 64'h0; // @[RegFile.scala 75:16:@44458.4]
  assign regs_183_io_reset = reset; // @[RegFile.scala 78:19:@44462.4]
  assign regs_183_io_enable = 1'h1; // @[RegFile.scala 74:20:@44456.4]
  assign regs_184_clock = clock; // @[:@44465.4]
  assign regs_184_reset = io_reset; // @[:@44466.4 RegFile.scala 76:16:@44473.4]
  assign regs_184_io_in = 64'h0; // @[RegFile.scala 75:16:@44472.4]
  assign regs_184_io_reset = reset; // @[RegFile.scala 78:19:@44476.4]
  assign regs_184_io_enable = 1'h1; // @[RegFile.scala 74:20:@44470.4]
  assign regs_185_clock = clock; // @[:@44479.4]
  assign regs_185_reset = io_reset; // @[:@44480.4 RegFile.scala 76:16:@44487.4]
  assign regs_185_io_in = 64'h0; // @[RegFile.scala 75:16:@44486.4]
  assign regs_185_io_reset = reset; // @[RegFile.scala 78:19:@44490.4]
  assign regs_185_io_enable = 1'h1; // @[RegFile.scala 74:20:@44484.4]
  assign regs_186_clock = clock; // @[:@44493.4]
  assign regs_186_reset = io_reset; // @[:@44494.4 RegFile.scala 76:16:@44501.4]
  assign regs_186_io_in = 64'h0; // @[RegFile.scala 75:16:@44500.4]
  assign regs_186_io_reset = reset; // @[RegFile.scala 78:19:@44504.4]
  assign regs_186_io_enable = 1'h1; // @[RegFile.scala 74:20:@44498.4]
  assign regs_187_clock = clock; // @[:@44507.4]
  assign regs_187_reset = io_reset; // @[:@44508.4 RegFile.scala 76:16:@44515.4]
  assign regs_187_io_in = 64'h0; // @[RegFile.scala 75:16:@44514.4]
  assign regs_187_io_reset = reset; // @[RegFile.scala 78:19:@44518.4]
  assign regs_187_io_enable = 1'h1; // @[RegFile.scala 74:20:@44512.4]
  assign regs_188_clock = clock; // @[:@44521.4]
  assign regs_188_reset = io_reset; // @[:@44522.4 RegFile.scala 76:16:@44529.4]
  assign regs_188_io_in = 64'h0; // @[RegFile.scala 75:16:@44528.4]
  assign regs_188_io_reset = reset; // @[RegFile.scala 78:19:@44532.4]
  assign regs_188_io_enable = 1'h1; // @[RegFile.scala 74:20:@44526.4]
  assign regs_189_clock = clock; // @[:@44535.4]
  assign regs_189_reset = io_reset; // @[:@44536.4 RegFile.scala 76:16:@44543.4]
  assign regs_189_io_in = 64'h0; // @[RegFile.scala 75:16:@44542.4]
  assign regs_189_io_reset = reset; // @[RegFile.scala 78:19:@44546.4]
  assign regs_189_io_enable = 1'h1; // @[RegFile.scala 74:20:@44540.4]
  assign regs_190_clock = clock; // @[:@44549.4]
  assign regs_190_reset = io_reset; // @[:@44550.4 RegFile.scala 76:16:@44557.4]
  assign regs_190_io_in = 64'h0; // @[RegFile.scala 75:16:@44556.4]
  assign regs_190_io_reset = reset; // @[RegFile.scala 78:19:@44560.4]
  assign regs_190_io_enable = 1'h1; // @[RegFile.scala 74:20:@44554.4]
  assign regs_191_clock = clock; // @[:@44563.4]
  assign regs_191_reset = io_reset; // @[:@44564.4 RegFile.scala 76:16:@44571.4]
  assign regs_191_io_in = 64'h0; // @[RegFile.scala 75:16:@44570.4]
  assign regs_191_io_reset = reset; // @[RegFile.scala 78:19:@44574.4]
  assign regs_191_io_enable = 1'h1; // @[RegFile.scala 74:20:@44568.4]
  assign regs_192_clock = clock; // @[:@44577.4]
  assign regs_192_reset = io_reset; // @[:@44578.4 RegFile.scala 76:16:@44585.4]
  assign regs_192_io_in = 64'h0; // @[RegFile.scala 75:16:@44584.4]
  assign regs_192_io_reset = reset; // @[RegFile.scala 78:19:@44588.4]
  assign regs_192_io_enable = 1'h1; // @[RegFile.scala 74:20:@44582.4]
  assign regs_193_clock = clock; // @[:@44591.4]
  assign regs_193_reset = io_reset; // @[:@44592.4 RegFile.scala 76:16:@44599.4]
  assign regs_193_io_in = 64'h0; // @[RegFile.scala 75:16:@44598.4]
  assign regs_193_io_reset = reset; // @[RegFile.scala 78:19:@44602.4]
  assign regs_193_io_enable = 1'h1; // @[RegFile.scala 74:20:@44596.4]
  assign regs_194_clock = clock; // @[:@44605.4]
  assign regs_194_reset = io_reset; // @[:@44606.4 RegFile.scala 76:16:@44613.4]
  assign regs_194_io_in = 64'h0; // @[RegFile.scala 75:16:@44612.4]
  assign regs_194_io_reset = reset; // @[RegFile.scala 78:19:@44616.4]
  assign regs_194_io_enable = 1'h1; // @[RegFile.scala 74:20:@44610.4]
  assign regs_195_clock = clock; // @[:@44619.4]
  assign regs_195_reset = io_reset; // @[:@44620.4 RegFile.scala 76:16:@44627.4]
  assign regs_195_io_in = 64'h0; // @[RegFile.scala 75:16:@44626.4]
  assign regs_195_io_reset = reset; // @[RegFile.scala 78:19:@44630.4]
  assign regs_195_io_enable = 1'h1; // @[RegFile.scala 74:20:@44624.4]
  assign regs_196_clock = clock; // @[:@44633.4]
  assign regs_196_reset = io_reset; // @[:@44634.4 RegFile.scala 76:16:@44641.4]
  assign regs_196_io_in = 64'h0; // @[RegFile.scala 75:16:@44640.4]
  assign regs_196_io_reset = reset; // @[RegFile.scala 78:19:@44644.4]
  assign regs_196_io_enable = 1'h1; // @[RegFile.scala 74:20:@44638.4]
  assign regs_197_clock = clock; // @[:@44647.4]
  assign regs_197_reset = io_reset; // @[:@44648.4 RegFile.scala 76:16:@44655.4]
  assign regs_197_io_in = 64'h0; // @[RegFile.scala 75:16:@44654.4]
  assign regs_197_io_reset = reset; // @[RegFile.scala 78:19:@44658.4]
  assign regs_197_io_enable = 1'h1; // @[RegFile.scala 74:20:@44652.4]
  assign regs_198_clock = clock; // @[:@44661.4]
  assign regs_198_reset = io_reset; // @[:@44662.4 RegFile.scala 76:16:@44669.4]
  assign regs_198_io_in = 64'h0; // @[RegFile.scala 75:16:@44668.4]
  assign regs_198_io_reset = reset; // @[RegFile.scala 78:19:@44672.4]
  assign regs_198_io_enable = 1'h1; // @[RegFile.scala 74:20:@44666.4]
  assign regs_199_clock = clock; // @[:@44675.4]
  assign regs_199_reset = io_reset; // @[:@44676.4 RegFile.scala 76:16:@44683.4]
  assign regs_199_io_in = 64'h0; // @[RegFile.scala 75:16:@44682.4]
  assign regs_199_io_reset = reset; // @[RegFile.scala 78:19:@44686.4]
  assign regs_199_io_enable = 1'h1; // @[RegFile.scala 74:20:@44680.4]
  assign regs_200_clock = clock; // @[:@44689.4]
  assign regs_200_reset = io_reset; // @[:@44690.4 RegFile.scala 76:16:@44697.4]
  assign regs_200_io_in = 64'h0; // @[RegFile.scala 75:16:@44696.4]
  assign regs_200_io_reset = reset; // @[RegFile.scala 78:19:@44700.4]
  assign regs_200_io_enable = 1'h1; // @[RegFile.scala 74:20:@44694.4]
  assign regs_201_clock = clock; // @[:@44703.4]
  assign regs_201_reset = io_reset; // @[:@44704.4 RegFile.scala 76:16:@44711.4]
  assign regs_201_io_in = 64'h0; // @[RegFile.scala 75:16:@44710.4]
  assign regs_201_io_reset = reset; // @[RegFile.scala 78:19:@44714.4]
  assign regs_201_io_enable = 1'h1; // @[RegFile.scala 74:20:@44708.4]
  assign regs_202_clock = clock; // @[:@44717.4]
  assign regs_202_reset = io_reset; // @[:@44718.4 RegFile.scala 76:16:@44725.4]
  assign regs_202_io_in = 64'h0; // @[RegFile.scala 75:16:@44724.4]
  assign regs_202_io_reset = reset; // @[RegFile.scala 78:19:@44728.4]
  assign regs_202_io_enable = 1'h1; // @[RegFile.scala 74:20:@44722.4]
  assign regs_203_clock = clock; // @[:@44731.4]
  assign regs_203_reset = io_reset; // @[:@44732.4 RegFile.scala 76:16:@44739.4]
  assign regs_203_io_in = 64'h0; // @[RegFile.scala 75:16:@44738.4]
  assign regs_203_io_reset = reset; // @[RegFile.scala 78:19:@44742.4]
  assign regs_203_io_enable = 1'h1; // @[RegFile.scala 74:20:@44736.4]
  assign regs_204_clock = clock; // @[:@44745.4]
  assign regs_204_reset = io_reset; // @[:@44746.4 RegFile.scala 76:16:@44753.4]
  assign regs_204_io_in = 64'h0; // @[RegFile.scala 75:16:@44752.4]
  assign regs_204_io_reset = reset; // @[RegFile.scala 78:19:@44756.4]
  assign regs_204_io_enable = 1'h1; // @[RegFile.scala 74:20:@44750.4]
  assign regs_205_clock = clock; // @[:@44759.4]
  assign regs_205_reset = io_reset; // @[:@44760.4 RegFile.scala 76:16:@44767.4]
  assign regs_205_io_in = 64'h0; // @[RegFile.scala 75:16:@44766.4]
  assign regs_205_io_reset = reset; // @[RegFile.scala 78:19:@44770.4]
  assign regs_205_io_enable = 1'h1; // @[RegFile.scala 74:20:@44764.4]
  assign regs_206_clock = clock; // @[:@44773.4]
  assign regs_206_reset = io_reset; // @[:@44774.4 RegFile.scala 76:16:@44781.4]
  assign regs_206_io_in = 64'h0; // @[RegFile.scala 75:16:@44780.4]
  assign regs_206_io_reset = reset; // @[RegFile.scala 78:19:@44784.4]
  assign regs_206_io_enable = 1'h1; // @[RegFile.scala 74:20:@44778.4]
  assign regs_207_clock = clock; // @[:@44787.4]
  assign regs_207_reset = io_reset; // @[:@44788.4 RegFile.scala 76:16:@44795.4]
  assign regs_207_io_in = 64'h0; // @[RegFile.scala 75:16:@44794.4]
  assign regs_207_io_reset = reset; // @[RegFile.scala 78:19:@44798.4]
  assign regs_207_io_enable = 1'h1; // @[RegFile.scala 74:20:@44792.4]
  assign regs_208_clock = clock; // @[:@44801.4]
  assign regs_208_reset = io_reset; // @[:@44802.4 RegFile.scala 76:16:@44809.4]
  assign regs_208_io_in = 64'h0; // @[RegFile.scala 75:16:@44808.4]
  assign regs_208_io_reset = reset; // @[RegFile.scala 78:19:@44812.4]
  assign regs_208_io_enable = 1'h1; // @[RegFile.scala 74:20:@44806.4]
  assign regs_209_clock = clock; // @[:@44815.4]
  assign regs_209_reset = io_reset; // @[:@44816.4 RegFile.scala 76:16:@44823.4]
  assign regs_209_io_in = 64'h0; // @[RegFile.scala 75:16:@44822.4]
  assign regs_209_io_reset = reset; // @[RegFile.scala 78:19:@44826.4]
  assign regs_209_io_enable = 1'h1; // @[RegFile.scala 74:20:@44820.4]
  assign regs_210_clock = clock; // @[:@44829.4]
  assign regs_210_reset = io_reset; // @[:@44830.4 RegFile.scala 76:16:@44837.4]
  assign regs_210_io_in = 64'h0; // @[RegFile.scala 75:16:@44836.4]
  assign regs_210_io_reset = reset; // @[RegFile.scala 78:19:@44840.4]
  assign regs_210_io_enable = 1'h1; // @[RegFile.scala 74:20:@44834.4]
  assign regs_211_clock = clock; // @[:@44843.4]
  assign regs_211_reset = io_reset; // @[:@44844.4 RegFile.scala 76:16:@44851.4]
  assign regs_211_io_in = 64'h0; // @[RegFile.scala 75:16:@44850.4]
  assign regs_211_io_reset = reset; // @[RegFile.scala 78:19:@44854.4]
  assign regs_211_io_enable = 1'h1; // @[RegFile.scala 74:20:@44848.4]
  assign regs_212_clock = clock; // @[:@44857.4]
  assign regs_212_reset = io_reset; // @[:@44858.4 RegFile.scala 76:16:@44865.4]
  assign regs_212_io_in = 64'h0; // @[RegFile.scala 75:16:@44864.4]
  assign regs_212_io_reset = reset; // @[RegFile.scala 78:19:@44868.4]
  assign regs_212_io_enable = 1'h1; // @[RegFile.scala 74:20:@44862.4]
  assign regs_213_clock = clock; // @[:@44871.4]
  assign regs_213_reset = io_reset; // @[:@44872.4 RegFile.scala 76:16:@44879.4]
  assign regs_213_io_in = 64'h0; // @[RegFile.scala 75:16:@44878.4]
  assign regs_213_io_reset = reset; // @[RegFile.scala 78:19:@44882.4]
  assign regs_213_io_enable = 1'h1; // @[RegFile.scala 74:20:@44876.4]
  assign regs_214_clock = clock; // @[:@44885.4]
  assign regs_214_reset = io_reset; // @[:@44886.4 RegFile.scala 76:16:@44893.4]
  assign regs_214_io_in = 64'h0; // @[RegFile.scala 75:16:@44892.4]
  assign regs_214_io_reset = reset; // @[RegFile.scala 78:19:@44896.4]
  assign regs_214_io_enable = 1'h1; // @[RegFile.scala 74:20:@44890.4]
  assign regs_215_clock = clock; // @[:@44899.4]
  assign regs_215_reset = io_reset; // @[:@44900.4 RegFile.scala 76:16:@44907.4]
  assign regs_215_io_in = 64'h0; // @[RegFile.scala 75:16:@44906.4]
  assign regs_215_io_reset = reset; // @[RegFile.scala 78:19:@44910.4]
  assign regs_215_io_enable = 1'h1; // @[RegFile.scala 74:20:@44904.4]
  assign regs_216_clock = clock; // @[:@44913.4]
  assign regs_216_reset = io_reset; // @[:@44914.4 RegFile.scala 76:16:@44921.4]
  assign regs_216_io_in = 64'h0; // @[RegFile.scala 75:16:@44920.4]
  assign regs_216_io_reset = reset; // @[RegFile.scala 78:19:@44924.4]
  assign regs_216_io_enable = 1'h1; // @[RegFile.scala 74:20:@44918.4]
  assign regs_217_clock = clock; // @[:@44927.4]
  assign regs_217_reset = io_reset; // @[:@44928.4 RegFile.scala 76:16:@44935.4]
  assign regs_217_io_in = 64'h0; // @[RegFile.scala 75:16:@44934.4]
  assign regs_217_io_reset = reset; // @[RegFile.scala 78:19:@44938.4]
  assign regs_217_io_enable = 1'h1; // @[RegFile.scala 74:20:@44932.4]
  assign regs_218_clock = clock; // @[:@44941.4]
  assign regs_218_reset = io_reset; // @[:@44942.4 RegFile.scala 76:16:@44949.4]
  assign regs_218_io_in = 64'h0; // @[RegFile.scala 75:16:@44948.4]
  assign regs_218_io_reset = reset; // @[RegFile.scala 78:19:@44952.4]
  assign regs_218_io_enable = 1'h1; // @[RegFile.scala 74:20:@44946.4]
  assign regs_219_clock = clock; // @[:@44955.4]
  assign regs_219_reset = io_reset; // @[:@44956.4 RegFile.scala 76:16:@44963.4]
  assign regs_219_io_in = 64'h0; // @[RegFile.scala 75:16:@44962.4]
  assign regs_219_io_reset = reset; // @[RegFile.scala 78:19:@44966.4]
  assign regs_219_io_enable = 1'h1; // @[RegFile.scala 74:20:@44960.4]
  assign regs_220_clock = clock; // @[:@44969.4]
  assign regs_220_reset = io_reset; // @[:@44970.4 RegFile.scala 76:16:@44977.4]
  assign regs_220_io_in = 64'h0; // @[RegFile.scala 75:16:@44976.4]
  assign regs_220_io_reset = reset; // @[RegFile.scala 78:19:@44980.4]
  assign regs_220_io_enable = 1'h1; // @[RegFile.scala 74:20:@44974.4]
  assign regs_221_clock = clock; // @[:@44983.4]
  assign regs_221_reset = io_reset; // @[:@44984.4 RegFile.scala 76:16:@44991.4]
  assign regs_221_io_in = 64'h0; // @[RegFile.scala 75:16:@44990.4]
  assign regs_221_io_reset = reset; // @[RegFile.scala 78:19:@44994.4]
  assign regs_221_io_enable = 1'h1; // @[RegFile.scala 74:20:@44988.4]
  assign regs_222_clock = clock; // @[:@44997.4]
  assign regs_222_reset = io_reset; // @[:@44998.4 RegFile.scala 76:16:@45005.4]
  assign regs_222_io_in = 64'h0; // @[RegFile.scala 75:16:@45004.4]
  assign regs_222_io_reset = reset; // @[RegFile.scala 78:19:@45008.4]
  assign regs_222_io_enable = 1'h1; // @[RegFile.scala 74:20:@45002.4]
  assign regs_223_clock = clock; // @[:@45011.4]
  assign regs_223_reset = io_reset; // @[:@45012.4 RegFile.scala 76:16:@45019.4]
  assign regs_223_io_in = 64'h0; // @[RegFile.scala 75:16:@45018.4]
  assign regs_223_io_reset = reset; // @[RegFile.scala 78:19:@45022.4]
  assign regs_223_io_enable = 1'h1; // @[RegFile.scala 74:20:@45016.4]
  assign regs_224_clock = clock; // @[:@45025.4]
  assign regs_224_reset = io_reset; // @[:@45026.4 RegFile.scala 76:16:@45033.4]
  assign regs_224_io_in = 64'h0; // @[RegFile.scala 75:16:@45032.4]
  assign regs_224_io_reset = reset; // @[RegFile.scala 78:19:@45036.4]
  assign regs_224_io_enable = 1'h1; // @[RegFile.scala 74:20:@45030.4]
  assign regs_225_clock = clock; // @[:@45039.4]
  assign regs_225_reset = io_reset; // @[:@45040.4 RegFile.scala 76:16:@45047.4]
  assign regs_225_io_in = 64'h0; // @[RegFile.scala 75:16:@45046.4]
  assign regs_225_io_reset = reset; // @[RegFile.scala 78:19:@45050.4]
  assign regs_225_io_enable = 1'h1; // @[RegFile.scala 74:20:@45044.4]
  assign regs_226_clock = clock; // @[:@45053.4]
  assign regs_226_reset = io_reset; // @[:@45054.4 RegFile.scala 76:16:@45061.4]
  assign regs_226_io_in = 64'h0; // @[RegFile.scala 75:16:@45060.4]
  assign regs_226_io_reset = reset; // @[RegFile.scala 78:19:@45064.4]
  assign regs_226_io_enable = 1'h1; // @[RegFile.scala 74:20:@45058.4]
  assign regs_227_clock = clock; // @[:@45067.4]
  assign regs_227_reset = io_reset; // @[:@45068.4 RegFile.scala 76:16:@45075.4]
  assign regs_227_io_in = 64'h0; // @[RegFile.scala 75:16:@45074.4]
  assign regs_227_io_reset = reset; // @[RegFile.scala 78:19:@45078.4]
  assign regs_227_io_enable = 1'h1; // @[RegFile.scala 74:20:@45072.4]
  assign regs_228_clock = clock; // @[:@45081.4]
  assign regs_228_reset = io_reset; // @[:@45082.4 RegFile.scala 76:16:@45089.4]
  assign regs_228_io_in = 64'h0; // @[RegFile.scala 75:16:@45088.4]
  assign regs_228_io_reset = reset; // @[RegFile.scala 78:19:@45092.4]
  assign regs_228_io_enable = 1'h1; // @[RegFile.scala 74:20:@45086.4]
  assign regs_229_clock = clock; // @[:@45095.4]
  assign regs_229_reset = io_reset; // @[:@45096.4 RegFile.scala 76:16:@45103.4]
  assign regs_229_io_in = 64'h0; // @[RegFile.scala 75:16:@45102.4]
  assign regs_229_io_reset = reset; // @[RegFile.scala 78:19:@45106.4]
  assign regs_229_io_enable = 1'h1; // @[RegFile.scala 74:20:@45100.4]
  assign regs_230_clock = clock; // @[:@45109.4]
  assign regs_230_reset = io_reset; // @[:@45110.4 RegFile.scala 76:16:@45117.4]
  assign regs_230_io_in = 64'h0; // @[RegFile.scala 75:16:@45116.4]
  assign regs_230_io_reset = reset; // @[RegFile.scala 78:19:@45120.4]
  assign regs_230_io_enable = 1'h1; // @[RegFile.scala 74:20:@45114.4]
  assign regs_231_clock = clock; // @[:@45123.4]
  assign regs_231_reset = io_reset; // @[:@45124.4 RegFile.scala 76:16:@45131.4]
  assign regs_231_io_in = 64'h0; // @[RegFile.scala 75:16:@45130.4]
  assign regs_231_io_reset = reset; // @[RegFile.scala 78:19:@45134.4]
  assign regs_231_io_enable = 1'h1; // @[RegFile.scala 74:20:@45128.4]
  assign regs_232_clock = clock; // @[:@45137.4]
  assign regs_232_reset = io_reset; // @[:@45138.4 RegFile.scala 76:16:@45145.4]
  assign regs_232_io_in = 64'h0; // @[RegFile.scala 75:16:@45144.4]
  assign regs_232_io_reset = reset; // @[RegFile.scala 78:19:@45148.4]
  assign regs_232_io_enable = 1'h1; // @[RegFile.scala 74:20:@45142.4]
  assign regs_233_clock = clock; // @[:@45151.4]
  assign regs_233_reset = io_reset; // @[:@45152.4 RegFile.scala 76:16:@45159.4]
  assign regs_233_io_in = 64'h0; // @[RegFile.scala 75:16:@45158.4]
  assign regs_233_io_reset = reset; // @[RegFile.scala 78:19:@45162.4]
  assign regs_233_io_enable = 1'h1; // @[RegFile.scala 74:20:@45156.4]
  assign regs_234_clock = clock; // @[:@45165.4]
  assign regs_234_reset = io_reset; // @[:@45166.4 RegFile.scala 76:16:@45173.4]
  assign regs_234_io_in = 64'h0; // @[RegFile.scala 75:16:@45172.4]
  assign regs_234_io_reset = reset; // @[RegFile.scala 78:19:@45176.4]
  assign regs_234_io_enable = 1'h1; // @[RegFile.scala 74:20:@45170.4]
  assign regs_235_clock = clock; // @[:@45179.4]
  assign regs_235_reset = io_reset; // @[:@45180.4 RegFile.scala 76:16:@45187.4]
  assign regs_235_io_in = 64'h0; // @[RegFile.scala 75:16:@45186.4]
  assign regs_235_io_reset = reset; // @[RegFile.scala 78:19:@45190.4]
  assign regs_235_io_enable = 1'h1; // @[RegFile.scala 74:20:@45184.4]
  assign regs_236_clock = clock; // @[:@45193.4]
  assign regs_236_reset = io_reset; // @[:@45194.4 RegFile.scala 76:16:@45201.4]
  assign regs_236_io_in = 64'h0; // @[RegFile.scala 75:16:@45200.4]
  assign regs_236_io_reset = reset; // @[RegFile.scala 78:19:@45204.4]
  assign regs_236_io_enable = 1'h1; // @[RegFile.scala 74:20:@45198.4]
  assign regs_237_clock = clock; // @[:@45207.4]
  assign regs_237_reset = io_reset; // @[:@45208.4 RegFile.scala 76:16:@45215.4]
  assign regs_237_io_in = 64'h0; // @[RegFile.scala 75:16:@45214.4]
  assign regs_237_io_reset = reset; // @[RegFile.scala 78:19:@45218.4]
  assign regs_237_io_enable = 1'h1; // @[RegFile.scala 74:20:@45212.4]
  assign regs_238_clock = clock; // @[:@45221.4]
  assign regs_238_reset = io_reset; // @[:@45222.4 RegFile.scala 76:16:@45229.4]
  assign regs_238_io_in = 64'h0; // @[RegFile.scala 75:16:@45228.4]
  assign regs_238_io_reset = reset; // @[RegFile.scala 78:19:@45232.4]
  assign regs_238_io_enable = 1'h1; // @[RegFile.scala 74:20:@45226.4]
  assign regs_239_clock = clock; // @[:@45235.4]
  assign regs_239_reset = io_reset; // @[:@45236.4 RegFile.scala 76:16:@45243.4]
  assign regs_239_io_in = 64'h0; // @[RegFile.scala 75:16:@45242.4]
  assign regs_239_io_reset = reset; // @[RegFile.scala 78:19:@45246.4]
  assign regs_239_io_enable = 1'h1; // @[RegFile.scala 74:20:@45240.4]
  assign regs_240_clock = clock; // @[:@45249.4]
  assign regs_240_reset = io_reset; // @[:@45250.4 RegFile.scala 76:16:@45257.4]
  assign regs_240_io_in = 64'h0; // @[RegFile.scala 75:16:@45256.4]
  assign regs_240_io_reset = reset; // @[RegFile.scala 78:19:@45260.4]
  assign regs_240_io_enable = 1'h1; // @[RegFile.scala 74:20:@45254.4]
  assign regs_241_clock = clock; // @[:@45263.4]
  assign regs_241_reset = io_reset; // @[:@45264.4 RegFile.scala 76:16:@45271.4]
  assign regs_241_io_in = 64'h0; // @[RegFile.scala 75:16:@45270.4]
  assign regs_241_io_reset = reset; // @[RegFile.scala 78:19:@45274.4]
  assign regs_241_io_enable = 1'h1; // @[RegFile.scala 74:20:@45268.4]
  assign regs_242_clock = clock; // @[:@45277.4]
  assign regs_242_reset = io_reset; // @[:@45278.4 RegFile.scala 76:16:@45285.4]
  assign regs_242_io_in = 64'h0; // @[RegFile.scala 75:16:@45284.4]
  assign regs_242_io_reset = reset; // @[RegFile.scala 78:19:@45288.4]
  assign regs_242_io_enable = 1'h1; // @[RegFile.scala 74:20:@45282.4]
  assign regs_243_clock = clock; // @[:@45291.4]
  assign regs_243_reset = io_reset; // @[:@45292.4 RegFile.scala 76:16:@45299.4]
  assign regs_243_io_in = 64'h0; // @[RegFile.scala 75:16:@45298.4]
  assign regs_243_io_reset = reset; // @[RegFile.scala 78:19:@45302.4]
  assign regs_243_io_enable = 1'h1; // @[RegFile.scala 74:20:@45296.4]
  assign regs_244_clock = clock; // @[:@45305.4]
  assign regs_244_reset = io_reset; // @[:@45306.4 RegFile.scala 76:16:@45313.4]
  assign regs_244_io_in = 64'h0; // @[RegFile.scala 75:16:@45312.4]
  assign regs_244_io_reset = reset; // @[RegFile.scala 78:19:@45316.4]
  assign regs_244_io_enable = 1'h1; // @[RegFile.scala 74:20:@45310.4]
  assign regs_245_clock = clock; // @[:@45319.4]
  assign regs_245_reset = io_reset; // @[:@45320.4 RegFile.scala 76:16:@45327.4]
  assign regs_245_io_in = 64'h0; // @[RegFile.scala 75:16:@45326.4]
  assign regs_245_io_reset = reset; // @[RegFile.scala 78:19:@45330.4]
  assign regs_245_io_enable = 1'h1; // @[RegFile.scala 74:20:@45324.4]
  assign regs_246_clock = clock; // @[:@45333.4]
  assign regs_246_reset = io_reset; // @[:@45334.4 RegFile.scala 76:16:@45341.4]
  assign regs_246_io_in = 64'h0; // @[RegFile.scala 75:16:@45340.4]
  assign regs_246_io_reset = reset; // @[RegFile.scala 78:19:@45344.4]
  assign regs_246_io_enable = 1'h1; // @[RegFile.scala 74:20:@45338.4]
  assign regs_247_clock = clock; // @[:@45347.4]
  assign regs_247_reset = io_reset; // @[:@45348.4 RegFile.scala 76:16:@45355.4]
  assign regs_247_io_in = 64'h0; // @[RegFile.scala 75:16:@45354.4]
  assign regs_247_io_reset = reset; // @[RegFile.scala 78:19:@45358.4]
  assign regs_247_io_enable = 1'h1; // @[RegFile.scala 74:20:@45352.4]
  assign regs_248_clock = clock; // @[:@45361.4]
  assign regs_248_reset = io_reset; // @[:@45362.4 RegFile.scala 76:16:@45369.4]
  assign regs_248_io_in = 64'h0; // @[RegFile.scala 75:16:@45368.4]
  assign regs_248_io_reset = reset; // @[RegFile.scala 78:19:@45372.4]
  assign regs_248_io_enable = 1'h1; // @[RegFile.scala 74:20:@45366.4]
  assign regs_249_clock = clock; // @[:@45375.4]
  assign regs_249_reset = io_reset; // @[:@45376.4 RegFile.scala 76:16:@45383.4]
  assign regs_249_io_in = 64'h0; // @[RegFile.scala 75:16:@45382.4]
  assign regs_249_io_reset = reset; // @[RegFile.scala 78:19:@45386.4]
  assign regs_249_io_enable = 1'h1; // @[RegFile.scala 74:20:@45380.4]
  assign regs_250_clock = clock; // @[:@45389.4]
  assign regs_250_reset = io_reset; // @[:@45390.4 RegFile.scala 76:16:@45397.4]
  assign regs_250_io_in = 64'h0; // @[RegFile.scala 75:16:@45396.4]
  assign regs_250_io_reset = reset; // @[RegFile.scala 78:19:@45400.4]
  assign regs_250_io_enable = 1'h1; // @[RegFile.scala 74:20:@45394.4]
  assign regs_251_clock = clock; // @[:@45403.4]
  assign regs_251_reset = io_reset; // @[:@45404.4 RegFile.scala 76:16:@45411.4]
  assign regs_251_io_in = 64'h0; // @[RegFile.scala 75:16:@45410.4]
  assign regs_251_io_reset = reset; // @[RegFile.scala 78:19:@45414.4]
  assign regs_251_io_enable = 1'h1; // @[RegFile.scala 74:20:@45408.4]
  assign regs_252_clock = clock; // @[:@45417.4]
  assign regs_252_reset = io_reset; // @[:@45418.4 RegFile.scala 76:16:@45425.4]
  assign regs_252_io_in = 64'h0; // @[RegFile.scala 75:16:@45424.4]
  assign regs_252_io_reset = reset; // @[RegFile.scala 78:19:@45428.4]
  assign regs_252_io_enable = 1'h1; // @[RegFile.scala 74:20:@45422.4]
  assign regs_253_clock = clock; // @[:@45431.4]
  assign regs_253_reset = io_reset; // @[:@45432.4 RegFile.scala 76:16:@45439.4]
  assign regs_253_io_in = 64'h0; // @[RegFile.scala 75:16:@45438.4]
  assign regs_253_io_reset = reset; // @[RegFile.scala 78:19:@45442.4]
  assign regs_253_io_enable = 1'h1; // @[RegFile.scala 74:20:@45436.4]
  assign regs_254_clock = clock; // @[:@45445.4]
  assign regs_254_reset = io_reset; // @[:@45446.4 RegFile.scala 76:16:@45453.4]
  assign regs_254_io_in = 64'h0; // @[RegFile.scala 75:16:@45452.4]
  assign regs_254_io_reset = reset; // @[RegFile.scala 78:19:@45456.4]
  assign regs_254_io_enable = 1'h1; // @[RegFile.scala 74:20:@45450.4]
  assign regs_255_clock = clock; // @[:@45459.4]
  assign regs_255_reset = io_reset; // @[:@45460.4 RegFile.scala 76:16:@45467.4]
  assign regs_255_io_in = 64'h0; // @[RegFile.scala 75:16:@45466.4]
  assign regs_255_io_reset = reset; // @[RegFile.scala 78:19:@45470.4]
  assign regs_255_io_enable = 1'h1; // @[RegFile.scala 74:20:@45464.4]
  assign regs_256_clock = clock; // @[:@45473.4]
  assign regs_256_reset = io_reset; // @[:@45474.4 RegFile.scala 76:16:@45481.4]
  assign regs_256_io_in = 64'h0; // @[RegFile.scala 75:16:@45480.4]
  assign regs_256_io_reset = reset; // @[RegFile.scala 78:19:@45484.4]
  assign regs_256_io_enable = 1'h1; // @[RegFile.scala 74:20:@45478.4]
  assign regs_257_clock = clock; // @[:@45487.4]
  assign regs_257_reset = io_reset; // @[:@45488.4 RegFile.scala 76:16:@45495.4]
  assign regs_257_io_in = 64'h0; // @[RegFile.scala 75:16:@45494.4]
  assign regs_257_io_reset = reset; // @[RegFile.scala 78:19:@45498.4]
  assign regs_257_io_enable = 1'h1; // @[RegFile.scala 74:20:@45492.4]
  assign regs_258_clock = clock; // @[:@45501.4]
  assign regs_258_reset = io_reset; // @[:@45502.4 RegFile.scala 76:16:@45509.4]
  assign regs_258_io_in = 64'h0; // @[RegFile.scala 75:16:@45508.4]
  assign regs_258_io_reset = reset; // @[RegFile.scala 78:19:@45512.4]
  assign regs_258_io_enable = 1'h1; // @[RegFile.scala 74:20:@45506.4]
  assign regs_259_clock = clock; // @[:@45515.4]
  assign regs_259_reset = io_reset; // @[:@45516.4 RegFile.scala 76:16:@45523.4]
  assign regs_259_io_in = 64'h0; // @[RegFile.scala 75:16:@45522.4]
  assign regs_259_io_reset = reset; // @[RegFile.scala 78:19:@45526.4]
  assign regs_259_io_enable = 1'h1; // @[RegFile.scala 74:20:@45520.4]
  assign regs_260_clock = clock; // @[:@45529.4]
  assign regs_260_reset = io_reset; // @[:@45530.4 RegFile.scala 76:16:@45537.4]
  assign regs_260_io_in = 64'h0; // @[RegFile.scala 75:16:@45536.4]
  assign regs_260_io_reset = reset; // @[RegFile.scala 78:19:@45540.4]
  assign regs_260_io_enable = 1'h1; // @[RegFile.scala 74:20:@45534.4]
  assign regs_261_clock = clock; // @[:@45543.4]
  assign regs_261_reset = io_reset; // @[:@45544.4 RegFile.scala 76:16:@45551.4]
  assign regs_261_io_in = 64'h0; // @[RegFile.scala 75:16:@45550.4]
  assign regs_261_io_reset = reset; // @[RegFile.scala 78:19:@45554.4]
  assign regs_261_io_enable = 1'h1; // @[RegFile.scala 74:20:@45548.4]
  assign regs_262_clock = clock; // @[:@45557.4]
  assign regs_262_reset = io_reset; // @[:@45558.4 RegFile.scala 76:16:@45565.4]
  assign regs_262_io_in = 64'h0; // @[RegFile.scala 75:16:@45564.4]
  assign regs_262_io_reset = reset; // @[RegFile.scala 78:19:@45568.4]
  assign regs_262_io_enable = 1'h1; // @[RegFile.scala 74:20:@45562.4]
  assign regs_263_clock = clock; // @[:@45571.4]
  assign regs_263_reset = io_reset; // @[:@45572.4 RegFile.scala 76:16:@45579.4]
  assign regs_263_io_in = 64'h0; // @[RegFile.scala 75:16:@45578.4]
  assign regs_263_io_reset = reset; // @[RegFile.scala 78:19:@45582.4]
  assign regs_263_io_enable = 1'h1; // @[RegFile.scala 74:20:@45576.4]
  assign regs_264_clock = clock; // @[:@45585.4]
  assign regs_264_reset = io_reset; // @[:@45586.4 RegFile.scala 76:16:@45593.4]
  assign regs_264_io_in = 64'h0; // @[RegFile.scala 75:16:@45592.4]
  assign regs_264_io_reset = reset; // @[RegFile.scala 78:19:@45596.4]
  assign regs_264_io_enable = 1'h1; // @[RegFile.scala 74:20:@45590.4]
  assign regs_265_clock = clock; // @[:@45599.4]
  assign regs_265_reset = io_reset; // @[:@45600.4 RegFile.scala 76:16:@45607.4]
  assign regs_265_io_in = 64'h0; // @[RegFile.scala 75:16:@45606.4]
  assign regs_265_io_reset = reset; // @[RegFile.scala 78:19:@45610.4]
  assign regs_265_io_enable = 1'h1; // @[RegFile.scala 74:20:@45604.4]
  assign regs_266_clock = clock; // @[:@45613.4]
  assign regs_266_reset = io_reset; // @[:@45614.4 RegFile.scala 76:16:@45621.4]
  assign regs_266_io_in = 64'h0; // @[RegFile.scala 75:16:@45620.4]
  assign regs_266_io_reset = reset; // @[RegFile.scala 78:19:@45624.4]
  assign regs_266_io_enable = 1'h1; // @[RegFile.scala 74:20:@45618.4]
  assign regs_267_clock = clock; // @[:@45627.4]
  assign regs_267_reset = io_reset; // @[:@45628.4 RegFile.scala 76:16:@45635.4]
  assign regs_267_io_in = 64'h0; // @[RegFile.scala 75:16:@45634.4]
  assign regs_267_io_reset = reset; // @[RegFile.scala 78:19:@45638.4]
  assign regs_267_io_enable = 1'h1; // @[RegFile.scala 74:20:@45632.4]
  assign regs_268_clock = clock; // @[:@45641.4]
  assign regs_268_reset = io_reset; // @[:@45642.4 RegFile.scala 76:16:@45649.4]
  assign regs_268_io_in = 64'h0; // @[RegFile.scala 75:16:@45648.4]
  assign regs_268_io_reset = reset; // @[RegFile.scala 78:19:@45652.4]
  assign regs_268_io_enable = 1'h1; // @[RegFile.scala 74:20:@45646.4]
  assign regs_269_clock = clock; // @[:@45655.4]
  assign regs_269_reset = io_reset; // @[:@45656.4 RegFile.scala 76:16:@45663.4]
  assign regs_269_io_in = 64'h0; // @[RegFile.scala 75:16:@45662.4]
  assign regs_269_io_reset = reset; // @[RegFile.scala 78:19:@45666.4]
  assign regs_269_io_enable = 1'h1; // @[RegFile.scala 74:20:@45660.4]
  assign regs_270_clock = clock; // @[:@45669.4]
  assign regs_270_reset = io_reset; // @[:@45670.4 RegFile.scala 76:16:@45677.4]
  assign regs_270_io_in = 64'h0; // @[RegFile.scala 75:16:@45676.4]
  assign regs_270_io_reset = reset; // @[RegFile.scala 78:19:@45680.4]
  assign regs_270_io_enable = 1'h1; // @[RegFile.scala 74:20:@45674.4]
  assign regs_271_clock = clock; // @[:@45683.4]
  assign regs_271_reset = io_reset; // @[:@45684.4 RegFile.scala 76:16:@45691.4]
  assign regs_271_io_in = 64'h0; // @[RegFile.scala 75:16:@45690.4]
  assign regs_271_io_reset = reset; // @[RegFile.scala 78:19:@45694.4]
  assign regs_271_io_enable = 1'h1; // @[RegFile.scala 74:20:@45688.4]
  assign regs_272_clock = clock; // @[:@45697.4]
  assign regs_272_reset = io_reset; // @[:@45698.4 RegFile.scala 76:16:@45705.4]
  assign regs_272_io_in = 64'h0; // @[RegFile.scala 75:16:@45704.4]
  assign regs_272_io_reset = reset; // @[RegFile.scala 78:19:@45708.4]
  assign regs_272_io_enable = 1'h1; // @[RegFile.scala 74:20:@45702.4]
  assign regs_273_clock = clock; // @[:@45711.4]
  assign regs_273_reset = io_reset; // @[:@45712.4 RegFile.scala 76:16:@45719.4]
  assign regs_273_io_in = 64'h0; // @[RegFile.scala 75:16:@45718.4]
  assign regs_273_io_reset = reset; // @[RegFile.scala 78:19:@45722.4]
  assign regs_273_io_enable = 1'h1; // @[RegFile.scala 74:20:@45716.4]
  assign regs_274_clock = clock; // @[:@45725.4]
  assign regs_274_reset = io_reset; // @[:@45726.4 RegFile.scala 76:16:@45733.4]
  assign regs_274_io_in = 64'h0; // @[RegFile.scala 75:16:@45732.4]
  assign regs_274_io_reset = reset; // @[RegFile.scala 78:19:@45736.4]
  assign regs_274_io_enable = 1'h1; // @[RegFile.scala 74:20:@45730.4]
  assign regs_275_clock = clock; // @[:@45739.4]
  assign regs_275_reset = io_reset; // @[:@45740.4 RegFile.scala 76:16:@45747.4]
  assign regs_275_io_in = 64'h0; // @[RegFile.scala 75:16:@45746.4]
  assign regs_275_io_reset = reset; // @[RegFile.scala 78:19:@45750.4]
  assign regs_275_io_enable = 1'h1; // @[RegFile.scala 74:20:@45744.4]
  assign regs_276_clock = clock; // @[:@45753.4]
  assign regs_276_reset = io_reset; // @[:@45754.4 RegFile.scala 76:16:@45761.4]
  assign regs_276_io_in = 64'h0; // @[RegFile.scala 75:16:@45760.4]
  assign regs_276_io_reset = reset; // @[RegFile.scala 78:19:@45764.4]
  assign regs_276_io_enable = 1'h1; // @[RegFile.scala 74:20:@45758.4]
  assign regs_277_clock = clock; // @[:@45767.4]
  assign regs_277_reset = io_reset; // @[:@45768.4 RegFile.scala 76:16:@45775.4]
  assign regs_277_io_in = 64'h0; // @[RegFile.scala 75:16:@45774.4]
  assign regs_277_io_reset = reset; // @[RegFile.scala 78:19:@45778.4]
  assign regs_277_io_enable = 1'h1; // @[RegFile.scala 74:20:@45772.4]
  assign regs_278_clock = clock; // @[:@45781.4]
  assign regs_278_reset = io_reset; // @[:@45782.4 RegFile.scala 76:16:@45789.4]
  assign regs_278_io_in = 64'h0; // @[RegFile.scala 75:16:@45788.4]
  assign regs_278_io_reset = reset; // @[RegFile.scala 78:19:@45792.4]
  assign regs_278_io_enable = 1'h1; // @[RegFile.scala 74:20:@45786.4]
  assign regs_279_clock = clock; // @[:@45795.4]
  assign regs_279_reset = io_reset; // @[:@45796.4 RegFile.scala 76:16:@45803.4]
  assign regs_279_io_in = 64'h0; // @[RegFile.scala 75:16:@45802.4]
  assign regs_279_io_reset = reset; // @[RegFile.scala 78:19:@45806.4]
  assign regs_279_io_enable = 1'h1; // @[RegFile.scala 74:20:@45800.4]
  assign regs_280_clock = clock; // @[:@45809.4]
  assign regs_280_reset = io_reset; // @[:@45810.4 RegFile.scala 76:16:@45817.4]
  assign regs_280_io_in = 64'h0; // @[RegFile.scala 75:16:@45816.4]
  assign regs_280_io_reset = reset; // @[RegFile.scala 78:19:@45820.4]
  assign regs_280_io_enable = 1'h1; // @[RegFile.scala 74:20:@45814.4]
  assign regs_281_clock = clock; // @[:@45823.4]
  assign regs_281_reset = io_reset; // @[:@45824.4 RegFile.scala 76:16:@45831.4]
  assign regs_281_io_in = 64'h0; // @[RegFile.scala 75:16:@45830.4]
  assign regs_281_io_reset = reset; // @[RegFile.scala 78:19:@45834.4]
  assign regs_281_io_enable = 1'h1; // @[RegFile.scala 74:20:@45828.4]
  assign regs_282_clock = clock; // @[:@45837.4]
  assign regs_282_reset = io_reset; // @[:@45838.4 RegFile.scala 76:16:@45845.4]
  assign regs_282_io_in = 64'h0; // @[RegFile.scala 75:16:@45844.4]
  assign regs_282_io_reset = reset; // @[RegFile.scala 78:19:@45848.4]
  assign regs_282_io_enable = 1'h1; // @[RegFile.scala 74:20:@45842.4]
  assign regs_283_clock = clock; // @[:@45851.4]
  assign regs_283_reset = io_reset; // @[:@45852.4 RegFile.scala 76:16:@45859.4]
  assign regs_283_io_in = 64'h0; // @[RegFile.scala 75:16:@45858.4]
  assign regs_283_io_reset = reset; // @[RegFile.scala 78:19:@45862.4]
  assign regs_283_io_enable = 1'h1; // @[RegFile.scala 74:20:@45856.4]
  assign regs_284_clock = clock; // @[:@45865.4]
  assign regs_284_reset = io_reset; // @[:@45866.4 RegFile.scala 76:16:@45873.4]
  assign regs_284_io_in = 64'h0; // @[RegFile.scala 75:16:@45872.4]
  assign regs_284_io_reset = reset; // @[RegFile.scala 78:19:@45876.4]
  assign regs_284_io_enable = 1'h1; // @[RegFile.scala 74:20:@45870.4]
  assign regs_285_clock = clock; // @[:@45879.4]
  assign regs_285_reset = io_reset; // @[:@45880.4 RegFile.scala 76:16:@45887.4]
  assign regs_285_io_in = 64'h0; // @[RegFile.scala 75:16:@45886.4]
  assign regs_285_io_reset = reset; // @[RegFile.scala 78:19:@45890.4]
  assign regs_285_io_enable = 1'h1; // @[RegFile.scala 74:20:@45884.4]
  assign regs_286_clock = clock; // @[:@45893.4]
  assign regs_286_reset = io_reset; // @[:@45894.4 RegFile.scala 76:16:@45901.4]
  assign regs_286_io_in = 64'h0; // @[RegFile.scala 75:16:@45900.4]
  assign regs_286_io_reset = reset; // @[RegFile.scala 78:19:@45904.4]
  assign regs_286_io_enable = 1'h1; // @[RegFile.scala 74:20:@45898.4]
  assign regs_287_clock = clock; // @[:@45907.4]
  assign regs_287_reset = io_reset; // @[:@45908.4 RegFile.scala 76:16:@45915.4]
  assign regs_287_io_in = 64'h0; // @[RegFile.scala 75:16:@45914.4]
  assign regs_287_io_reset = reset; // @[RegFile.scala 78:19:@45918.4]
  assign regs_287_io_enable = 1'h1; // @[RegFile.scala 74:20:@45912.4]
  assign regs_288_clock = clock; // @[:@45921.4]
  assign regs_288_reset = io_reset; // @[:@45922.4 RegFile.scala 76:16:@45929.4]
  assign regs_288_io_in = 64'h0; // @[RegFile.scala 75:16:@45928.4]
  assign regs_288_io_reset = reset; // @[RegFile.scala 78:19:@45932.4]
  assign regs_288_io_enable = 1'h1; // @[RegFile.scala 74:20:@45926.4]
  assign regs_289_clock = clock; // @[:@45935.4]
  assign regs_289_reset = io_reset; // @[:@45936.4 RegFile.scala 76:16:@45943.4]
  assign regs_289_io_in = 64'h0; // @[RegFile.scala 75:16:@45942.4]
  assign regs_289_io_reset = reset; // @[RegFile.scala 78:19:@45946.4]
  assign regs_289_io_enable = 1'h1; // @[RegFile.scala 74:20:@45940.4]
  assign regs_290_clock = clock; // @[:@45949.4]
  assign regs_290_reset = io_reset; // @[:@45950.4 RegFile.scala 76:16:@45957.4]
  assign regs_290_io_in = 64'h0; // @[RegFile.scala 75:16:@45956.4]
  assign regs_290_io_reset = reset; // @[RegFile.scala 78:19:@45960.4]
  assign regs_290_io_enable = 1'h1; // @[RegFile.scala 74:20:@45954.4]
  assign regs_291_clock = clock; // @[:@45963.4]
  assign regs_291_reset = io_reset; // @[:@45964.4 RegFile.scala 76:16:@45971.4]
  assign regs_291_io_in = 64'h0; // @[RegFile.scala 75:16:@45970.4]
  assign regs_291_io_reset = reset; // @[RegFile.scala 78:19:@45974.4]
  assign regs_291_io_enable = 1'h1; // @[RegFile.scala 74:20:@45968.4]
  assign regs_292_clock = clock; // @[:@45977.4]
  assign regs_292_reset = io_reset; // @[:@45978.4 RegFile.scala 76:16:@45985.4]
  assign regs_292_io_in = 64'h0; // @[RegFile.scala 75:16:@45984.4]
  assign regs_292_io_reset = reset; // @[RegFile.scala 78:19:@45988.4]
  assign regs_292_io_enable = 1'h1; // @[RegFile.scala 74:20:@45982.4]
  assign regs_293_clock = clock; // @[:@45991.4]
  assign regs_293_reset = io_reset; // @[:@45992.4 RegFile.scala 76:16:@45999.4]
  assign regs_293_io_in = 64'h0; // @[RegFile.scala 75:16:@45998.4]
  assign regs_293_io_reset = reset; // @[RegFile.scala 78:19:@46002.4]
  assign regs_293_io_enable = 1'h1; // @[RegFile.scala 74:20:@45996.4]
  assign regs_294_clock = clock; // @[:@46005.4]
  assign regs_294_reset = io_reset; // @[:@46006.4 RegFile.scala 76:16:@46013.4]
  assign regs_294_io_in = 64'h0; // @[RegFile.scala 75:16:@46012.4]
  assign regs_294_io_reset = reset; // @[RegFile.scala 78:19:@46016.4]
  assign regs_294_io_enable = 1'h1; // @[RegFile.scala 74:20:@46010.4]
  assign regs_295_clock = clock; // @[:@46019.4]
  assign regs_295_reset = io_reset; // @[:@46020.4 RegFile.scala 76:16:@46027.4]
  assign regs_295_io_in = 64'h0; // @[RegFile.scala 75:16:@46026.4]
  assign regs_295_io_reset = reset; // @[RegFile.scala 78:19:@46030.4]
  assign regs_295_io_enable = 1'h1; // @[RegFile.scala 74:20:@46024.4]
  assign regs_296_clock = clock; // @[:@46033.4]
  assign regs_296_reset = io_reset; // @[:@46034.4 RegFile.scala 76:16:@46041.4]
  assign regs_296_io_in = 64'h0; // @[RegFile.scala 75:16:@46040.4]
  assign regs_296_io_reset = reset; // @[RegFile.scala 78:19:@46044.4]
  assign regs_296_io_enable = 1'h1; // @[RegFile.scala 74:20:@46038.4]
  assign regs_297_clock = clock; // @[:@46047.4]
  assign regs_297_reset = io_reset; // @[:@46048.4 RegFile.scala 76:16:@46055.4]
  assign regs_297_io_in = 64'h0; // @[RegFile.scala 75:16:@46054.4]
  assign regs_297_io_reset = reset; // @[RegFile.scala 78:19:@46058.4]
  assign regs_297_io_enable = 1'h1; // @[RegFile.scala 74:20:@46052.4]
  assign regs_298_clock = clock; // @[:@46061.4]
  assign regs_298_reset = io_reset; // @[:@46062.4 RegFile.scala 76:16:@46069.4]
  assign regs_298_io_in = 64'h0; // @[RegFile.scala 75:16:@46068.4]
  assign regs_298_io_reset = reset; // @[RegFile.scala 78:19:@46072.4]
  assign regs_298_io_enable = 1'h1; // @[RegFile.scala 74:20:@46066.4]
  assign regs_299_clock = clock; // @[:@46075.4]
  assign regs_299_reset = io_reset; // @[:@46076.4 RegFile.scala 76:16:@46083.4]
  assign regs_299_io_in = 64'h0; // @[RegFile.scala 75:16:@46082.4]
  assign regs_299_io_reset = reset; // @[RegFile.scala 78:19:@46086.4]
  assign regs_299_io_enable = 1'h1; // @[RegFile.scala 74:20:@46080.4]
  assign regs_300_clock = clock; // @[:@46089.4]
  assign regs_300_reset = io_reset; // @[:@46090.4 RegFile.scala 76:16:@46097.4]
  assign regs_300_io_in = 64'h0; // @[RegFile.scala 75:16:@46096.4]
  assign regs_300_io_reset = reset; // @[RegFile.scala 78:19:@46100.4]
  assign regs_300_io_enable = 1'h1; // @[RegFile.scala 74:20:@46094.4]
  assign regs_301_clock = clock; // @[:@46103.4]
  assign regs_301_reset = io_reset; // @[:@46104.4 RegFile.scala 76:16:@46111.4]
  assign regs_301_io_in = 64'h0; // @[RegFile.scala 75:16:@46110.4]
  assign regs_301_io_reset = reset; // @[RegFile.scala 78:19:@46114.4]
  assign regs_301_io_enable = 1'h1; // @[RegFile.scala 74:20:@46108.4]
  assign regs_302_clock = clock; // @[:@46117.4]
  assign regs_302_reset = io_reset; // @[:@46118.4 RegFile.scala 76:16:@46125.4]
  assign regs_302_io_in = 64'h0; // @[RegFile.scala 75:16:@46124.4]
  assign regs_302_io_reset = reset; // @[RegFile.scala 78:19:@46128.4]
  assign regs_302_io_enable = 1'h1; // @[RegFile.scala 74:20:@46122.4]
  assign regs_303_clock = clock; // @[:@46131.4]
  assign regs_303_reset = io_reset; // @[:@46132.4 RegFile.scala 76:16:@46139.4]
  assign regs_303_io_in = 64'h0; // @[RegFile.scala 75:16:@46138.4]
  assign regs_303_io_reset = reset; // @[RegFile.scala 78:19:@46142.4]
  assign regs_303_io_enable = 1'h1; // @[RegFile.scala 74:20:@46136.4]
  assign regs_304_clock = clock; // @[:@46145.4]
  assign regs_304_reset = io_reset; // @[:@46146.4 RegFile.scala 76:16:@46153.4]
  assign regs_304_io_in = 64'h0; // @[RegFile.scala 75:16:@46152.4]
  assign regs_304_io_reset = reset; // @[RegFile.scala 78:19:@46156.4]
  assign regs_304_io_enable = 1'h1; // @[RegFile.scala 74:20:@46150.4]
  assign regs_305_clock = clock; // @[:@46159.4]
  assign regs_305_reset = io_reset; // @[:@46160.4 RegFile.scala 76:16:@46167.4]
  assign regs_305_io_in = 64'h0; // @[RegFile.scala 75:16:@46166.4]
  assign regs_305_io_reset = reset; // @[RegFile.scala 78:19:@46170.4]
  assign regs_305_io_enable = 1'h1; // @[RegFile.scala 74:20:@46164.4]
  assign regs_306_clock = clock; // @[:@46173.4]
  assign regs_306_reset = io_reset; // @[:@46174.4 RegFile.scala 76:16:@46181.4]
  assign regs_306_io_in = 64'h0; // @[RegFile.scala 75:16:@46180.4]
  assign regs_306_io_reset = reset; // @[RegFile.scala 78:19:@46184.4]
  assign regs_306_io_enable = 1'h1; // @[RegFile.scala 74:20:@46178.4]
  assign regs_307_clock = clock; // @[:@46187.4]
  assign regs_307_reset = io_reset; // @[:@46188.4 RegFile.scala 76:16:@46195.4]
  assign regs_307_io_in = 64'h0; // @[RegFile.scala 75:16:@46194.4]
  assign regs_307_io_reset = reset; // @[RegFile.scala 78:19:@46198.4]
  assign regs_307_io_enable = 1'h1; // @[RegFile.scala 74:20:@46192.4]
  assign regs_308_clock = clock; // @[:@46201.4]
  assign regs_308_reset = io_reset; // @[:@46202.4 RegFile.scala 76:16:@46209.4]
  assign regs_308_io_in = 64'h0; // @[RegFile.scala 75:16:@46208.4]
  assign regs_308_io_reset = reset; // @[RegFile.scala 78:19:@46212.4]
  assign regs_308_io_enable = 1'h1; // @[RegFile.scala 74:20:@46206.4]
  assign regs_309_clock = clock; // @[:@46215.4]
  assign regs_309_reset = io_reset; // @[:@46216.4 RegFile.scala 76:16:@46223.4]
  assign regs_309_io_in = 64'h0; // @[RegFile.scala 75:16:@46222.4]
  assign regs_309_io_reset = reset; // @[RegFile.scala 78:19:@46226.4]
  assign regs_309_io_enable = 1'h1; // @[RegFile.scala 74:20:@46220.4]
  assign regs_310_clock = clock; // @[:@46229.4]
  assign regs_310_reset = io_reset; // @[:@46230.4 RegFile.scala 76:16:@46237.4]
  assign regs_310_io_in = 64'h0; // @[RegFile.scala 75:16:@46236.4]
  assign regs_310_io_reset = reset; // @[RegFile.scala 78:19:@46240.4]
  assign regs_310_io_enable = 1'h1; // @[RegFile.scala 74:20:@46234.4]
  assign regs_311_clock = clock; // @[:@46243.4]
  assign regs_311_reset = io_reset; // @[:@46244.4 RegFile.scala 76:16:@46251.4]
  assign regs_311_io_in = 64'h0; // @[RegFile.scala 75:16:@46250.4]
  assign regs_311_io_reset = reset; // @[RegFile.scala 78:19:@46254.4]
  assign regs_311_io_enable = 1'h1; // @[RegFile.scala 74:20:@46248.4]
  assign regs_312_clock = clock; // @[:@46257.4]
  assign regs_312_reset = io_reset; // @[:@46258.4 RegFile.scala 76:16:@46265.4]
  assign regs_312_io_in = 64'h0; // @[RegFile.scala 75:16:@46264.4]
  assign regs_312_io_reset = reset; // @[RegFile.scala 78:19:@46268.4]
  assign regs_312_io_enable = 1'h1; // @[RegFile.scala 74:20:@46262.4]
  assign regs_313_clock = clock; // @[:@46271.4]
  assign regs_313_reset = io_reset; // @[:@46272.4 RegFile.scala 76:16:@46279.4]
  assign regs_313_io_in = 64'h0; // @[RegFile.scala 75:16:@46278.4]
  assign regs_313_io_reset = reset; // @[RegFile.scala 78:19:@46282.4]
  assign regs_313_io_enable = 1'h1; // @[RegFile.scala 74:20:@46276.4]
  assign regs_314_clock = clock; // @[:@46285.4]
  assign regs_314_reset = io_reset; // @[:@46286.4 RegFile.scala 76:16:@46293.4]
  assign regs_314_io_in = 64'h0; // @[RegFile.scala 75:16:@46292.4]
  assign regs_314_io_reset = reset; // @[RegFile.scala 78:19:@46296.4]
  assign regs_314_io_enable = 1'h1; // @[RegFile.scala 74:20:@46290.4]
  assign regs_315_clock = clock; // @[:@46299.4]
  assign regs_315_reset = io_reset; // @[:@46300.4 RegFile.scala 76:16:@46307.4]
  assign regs_315_io_in = 64'h0; // @[RegFile.scala 75:16:@46306.4]
  assign regs_315_io_reset = reset; // @[RegFile.scala 78:19:@46310.4]
  assign regs_315_io_enable = 1'h1; // @[RegFile.scala 74:20:@46304.4]
  assign regs_316_clock = clock; // @[:@46313.4]
  assign regs_316_reset = io_reset; // @[:@46314.4 RegFile.scala 76:16:@46321.4]
  assign regs_316_io_in = 64'h0; // @[RegFile.scala 75:16:@46320.4]
  assign regs_316_io_reset = reset; // @[RegFile.scala 78:19:@46324.4]
  assign regs_316_io_enable = 1'h1; // @[RegFile.scala 74:20:@46318.4]
  assign regs_317_clock = clock; // @[:@46327.4]
  assign regs_317_reset = io_reset; // @[:@46328.4 RegFile.scala 76:16:@46335.4]
  assign regs_317_io_in = 64'h0; // @[RegFile.scala 75:16:@46334.4]
  assign regs_317_io_reset = reset; // @[RegFile.scala 78:19:@46338.4]
  assign regs_317_io_enable = 1'h1; // @[RegFile.scala 74:20:@46332.4]
  assign regs_318_clock = clock; // @[:@46341.4]
  assign regs_318_reset = io_reset; // @[:@46342.4 RegFile.scala 76:16:@46349.4]
  assign regs_318_io_in = 64'h0; // @[RegFile.scala 75:16:@46348.4]
  assign regs_318_io_reset = reset; // @[RegFile.scala 78:19:@46352.4]
  assign regs_318_io_enable = 1'h1; // @[RegFile.scala 74:20:@46346.4]
  assign regs_319_clock = clock; // @[:@46355.4]
  assign regs_319_reset = io_reset; // @[:@46356.4 RegFile.scala 76:16:@46363.4]
  assign regs_319_io_in = 64'h0; // @[RegFile.scala 75:16:@46362.4]
  assign regs_319_io_reset = reset; // @[RegFile.scala 78:19:@46366.4]
  assign regs_319_io_enable = 1'h1; // @[RegFile.scala 74:20:@46360.4]
  assign regs_320_clock = clock; // @[:@46369.4]
  assign regs_320_reset = io_reset; // @[:@46370.4 RegFile.scala 76:16:@46377.4]
  assign regs_320_io_in = 64'h0; // @[RegFile.scala 75:16:@46376.4]
  assign regs_320_io_reset = reset; // @[RegFile.scala 78:19:@46380.4]
  assign regs_320_io_enable = 1'h1; // @[RegFile.scala 74:20:@46374.4]
  assign regs_321_clock = clock; // @[:@46383.4]
  assign regs_321_reset = io_reset; // @[:@46384.4 RegFile.scala 76:16:@46391.4]
  assign regs_321_io_in = 64'h0; // @[RegFile.scala 75:16:@46390.4]
  assign regs_321_io_reset = reset; // @[RegFile.scala 78:19:@46394.4]
  assign regs_321_io_enable = 1'h1; // @[RegFile.scala 74:20:@46388.4]
  assign regs_322_clock = clock; // @[:@46397.4]
  assign regs_322_reset = io_reset; // @[:@46398.4 RegFile.scala 76:16:@46405.4]
  assign regs_322_io_in = 64'h0; // @[RegFile.scala 75:16:@46404.4]
  assign regs_322_io_reset = reset; // @[RegFile.scala 78:19:@46408.4]
  assign regs_322_io_enable = 1'h1; // @[RegFile.scala 74:20:@46402.4]
  assign regs_323_clock = clock; // @[:@46411.4]
  assign regs_323_reset = io_reset; // @[:@46412.4 RegFile.scala 76:16:@46419.4]
  assign regs_323_io_in = 64'h0; // @[RegFile.scala 75:16:@46418.4]
  assign regs_323_io_reset = reset; // @[RegFile.scala 78:19:@46422.4]
  assign regs_323_io_enable = 1'h1; // @[RegFile.scala 74:20:@46416.4]
  assign regs_324_clock = clock; // @[:@46425.4]
  assign regs_324_reset = io_reset; // @[:@46426.4 RegFile.scala 76:16:@46433.4]
  assign regs_324_io_in = 64'h0; // @[RegFile.scala 75:16:@46432.4]
  assign regs_324_io_reset = reset; // @[RegFile.scala 78:19:@46436.4]
  assign regs_324_io_enable = 1'h1; // @[RegFile.scala 74:20:@46430.4]
  assign regs_325_clock = clock; // @[:@46439.4]
  assign regs_325_reset = io_reset; // @[:@46440.4 RegFile.scala 76:16:@46447.4]
  assign regs_325_io_in = 64'h0; // @[RegFile.scala 75:16:@46446.4]
  assign regs_325_io_reset = reset; // @[RegFile.scala 78:19:@46450.4]
  assign regs_325_io_enable = 1'h1; // @[RegFile.scala 74:20:@46444.4]
  assign regs_326_clock = clock; // @[:@46453.4]
  assign regs_326_reset = io_reset; // @[:@46454.4 RegFile.scala 76:16:@46461.4]
  assign regs_326_io_in = 64'h0; // @[RegFile.scala 75:16:@46460.4]
  assign regs_326_io_reset = reset; // @[RegFile.scala 78:19:@46464.4]
  assign regs_326_io_enable = 1'h1; // @[RegFile.scala 74:20:@46458.4]
  assign regs_327_clock = clock; // @[:@46467.4]
  assign regs_327_reset = io_reset; // @[:@46468.4 RegFile.scala 76:16:@46475.4]
  assign regs_327_io_in = 64'h0; // @[RegFile.scala 75:16:@46474.4]
  assign regs_327_io_reset = reset; // @[RegFile.scala 78:19:@46478.4]
  assign regs_327_io_enable = 1'h1; // @[RegFile.scala 74:20:@46472.4]
  assign regs_328_clock = clock; // @[:@46481.4]
  assign regs_328_reset = io_reset; // @[:@46482.4 RegFile.scala 76:16:@46489.4]
  assign regs_328_io_in = 64'h0; // @[RegFile.scala 75:16:@46488.4]
  assign regs_328_io_reset = reset; // @[RegFile.scala 78:19:@46492.4]
  assign regs_328_io_enable = 1'h1; // @[RegFile.scala 74:20:@46486.4]
  assign regs_329_clock = clock; // @[:@46495.4]
  assign regs_329_reset = io_reset; // @[:@46496.4 RegFile.scala 76:16:@46503.4]
  assign regs_329_io_in = 64'h0; // @[RegFile.scala 75:16:@46502.4]
  assign regs_329_io_reset = reset; // @[RegFile.scala 78:19:@46506.4]
  assign regs_329_io_enable = 1'h1; // @[RegFile.scala 74:20:@46500.4]
  assign regs_330_clock = clock; // @[:@46509.4]
  assign regs_330_reset = io_reset; // @[:@46510.4 RegFile.scala 76:16:@46517.4]
  assign regs_330_io_in = 64'h0; // @[RegFile.scala 75:16:@46516.4]
  assign regs_330_io_reset = reset; // @[RegFile.scala 78:19:@46520.4]
  assign regs_330_io_enable = 1'h1; // @[RegFile.scala 74:20:@46514.4]
  assign regs_331_clock = clock; // @[:@46523.4]
  assign regs_331_reset = io_reset; // @[:@46524.4 RegFile.scala 76:16:@46531.4]
  assign regs_331_io_in = 64'h0; // @[RegFile.scala 75:16:@46530.4]
  assign regs_331_io_reset = reset; // @[RegFile.scala 78:19:@46534.4]
  assign regs_331_io_enable = 1'h1; // @[RegFile.scala 74:20:@46528.4]
  assign regs_332_clock = clock; // @[:@46537.4]
  assign regs_332_reset = io_reset; // @[:@46538.4 RegFile.scala 76:16:@46545.4]
  assign regs_332_io_in = 64'h0; // @[RegFile.scala 75:16:@46544.4]
  assign regs_332_io_reset = reset; // @[RegFile.scala 78:19:@46548.4]
  assign regs_332_io_enable = 1'h1; // @[RegFile.scala 74:20:@46542.4]
  assign regs_333_clock = clock; // @[:@46551.4]
  assign regs_333_reset = io_reset; // @[:@46552.4 RegFile.scala 76:16:@46559.4]
  assign regs_333_io_in = 64'h0; // @[RegFile.scala 75:16:@46558.4]
  assign regs_333_io_reset = reset; // @[RegFile.scala 78:19:@46562.4]
  assign regs_333_io_enable = 1'h1; // @[RegFile.scala 74:20:@46556.4]
  assign regs_334_clock = clock; // @[:@46565.4]
  assign regs_334_reset = io_reset; // @[:@46566.4 RegFile.scala 76:16:@46573.4]
  assign regs_334_io_in = 64'h0; // @[RegFile.scala 75:16:@46572.4]
  assign regs_334_io_reset = reset; // @[RegFile.scala 78:19:@46576.4]
  assign regs_334_io_enable = 1'h1; // @[RegFile.scala 74:20:@46570.4]
  assign regs_335_clock = clock; // @[:@46579.4]
  assign regs_335_reset = io_reset; // @[:@46580.4 RegFile.scala 76:16:@46587.4]
  assign regs_335_io_in = 64'h0; // @[RegFile.scala 75:16:@46586.4]
  assign regs_335_io_reset = reset; // @[RegFile.scala 78:19:@46590.4]
  assign regs_335_io_enable = 1'h1; // @[RegFile.scala 74:20:@46584.4]
  assign regs_336_clock = clock; // @[:@46593.4]
  assign regs_336_reset = io_reset; // @[:@46594.4 RegFile.scala 76:16:@46601.4]
  assign regs_336_io_in = 64'h0; // @[RegFile.scala 75:16:@46600.4]
  assign regs_336_io_reset = reset; // @[RegFile.scala 78:19:@46604.4]
  assign regs_336_io_enable = 1'h1; // @[RegFile.scala 74:20:@46598.4]
  assign regs_337_clock = clock; // @[:@46607.4]
  assign regs_337_reset = io_reset; // @[:@46608.4 RegFile.scala 76:16:@46615.4]
  assign regs_337_io_in = 64'h0; // @[RegFile.scala 75:16:@46614.4]
  assign regs_337_io_reset = reset; // @[RegFile.scala 78:19:@46618.4]
  assign regs_337_io_enable = 1'h1; // @[RegFile.scala 74:20:@46612.4]
  assign regs_338_clock = clock; // @[:@46621.4]
  assign regs_338_reset = io_reset; // @[:@46622.4 RegFile.scala 76:16:@46629.4]
  assign regs_338_io_in = 64'h0; // @[RegFile.scala 75:16:@46628.4]
  assign regs_338_io_reset = reset; // @[RegFile.scala 78:19:@46632.4]
  assign regs_338_io_enable = 1'h1; // @[RegFile.scala 74:20:@46626.4]
  assign regs_339_clock = clock; // @[:@46635.4]
  assign regs_339_reset = io_reset; // @[:@46636.4 RegFile.scala 76:16:@46643.4]
  assign regs_339_io_in = 64'h0; // @[RegFile.scala 75:16:@46642.4]
  assign regs_339_io_reset = reset; // @[RegFile.scala 78:19:@46646.4]
  assign regs_339_io_enable = 1'h1; // @[RegFile.scala 74:20:@46640.4]
  assign regs_340_clock = clock; // @[:@46649.4]
  assign regs_340_reset = io_reset; // @[:@46650.4 RegFile.scala 76:16:@46657.4]
  assign regs_340_io_in = 64'h0; // @[RegFile.scala 75:16:@46656.4]
  assign regs_340_io_reset = reset; // @[RegFile.scala 78:19:@46660.4]
  assign regs_340_io_enable = 1'h1; // @[RegFile.scala 74:20:@46654.4]
  assign regs_341_clock = clock; // @[:@46663.4]
  assign regs_341_reset = io_reset; // @[:@46664.4 RegFile.scala 76:16:@46671.4]
  assign regs_341_io_in = 64'h0; // @[RegFile.scala 75:16:@46670.4]
  assign regs_341_io_reset = reset; // @[RegFile.scala 78:19:@46674.4]
  assign regs_341_io_enable = 1'h1; // @[RegFile.scala 74:20:@46668.4]
  assign regs_342_clock = clock; // @[:@46677.4]
  assign regs_342_reset = io_reset; // @[:@46678.4 RegFile.scala 76:16:@46685.4]
  assign regs_342_io_in = 64'h0; // @[RegFile.scala 75:16:@46684.4]
  assign regs_342_io_reset = reset; // @[RegFile.scala 78:19:@46688.4]
  assign regs_342_io_enable = 1'h1; // @[RegFile.scala 74:20:@46682.4]
  assign regs_343_clock = clock; // @[:@46691.4]
  assign regs_343_reset = io_reset; // @[:@46692.4 RegFile.scala 76:16:@46699.4]
  assign regs_343_io_in = 64'h0; // @[RegFile.scala 75:16:@46698.4]
  assign regs_343_io_reset = reset; // @[RegFile.scala 78:19:@46702.4]
  assign regs_343_io_enable = 1'h1; // @[RegFile.scala 74:20:@46696.4]
  assign regs_344_clock = clock; // @[:@46705.4]
  assign regs_344_reset = io_reset; // @[:@46706.4 RegFile.scala 76:16:@46713.4]
  assign regs_344_io_in = 64'h0; // @[RegFile.scala 75:16:@46712.4]
  assign regs_344_io_reset = reset; // @[RegFile.scala 78:19:@46716.4]
  assign regs_344_io_enable = 1'h1; // @[RegFile.scala 74:20:@46710.4]
  assign regs_345_clock = clock; // @[:@46719.4]
  assign regs_345_reset = io_reset; // @[:@46720.4 RegFile.scala 76:16:@46727.4]
  assign regs_345_io_in = 64'h0; // @[RegFile.scala 75:16:@46726.4]
  assign regs_345_io_reset = reset; // @[RegFile.scala 78:19:@46730.4]
  assign regs_345_io_enable = 1'h1; // @[RegFile.scala 74:20:@46724.4]
  assign regs_346_clock = clock; // @[:@46733.4]
  assign regs_346_reset = io_reset; // @[:@46734.4 RegFile.scala 76:16:@46741.4]
  assign regs_346_io_in = 64'h0; // @[RegFile.scala 75:16:@46740.4]
  assign regs_346_io_reset = reset; // @[RegFile.scala 78:19:@46744.4]
  assign regs_346_io_enable = 1'h1; // @[RegFile.scala 74:20:@46738.4]
  assign regs_347_clock = clock; // @[:@46747.4]
  assign regs_347_reset = io_reset; // @[:@46748.4 RegFile.scala 76:16:@46755.4]
  assign regs_347_io_in = 64'h0; // @[RegFile.scala 75:16:@46754.4]
  assign regs_347_io_reset = reset; // @[RegFile.scala 78:19:@46758.4]
  assign regs_347_io_enable = 1'h1; // @[RegFile.scala 74:20:@46752.4]
  assign regs_348_clock = clock; // @[:@46761.4]
  assign regs_348_reset = io_reset; // @[:@46762.4 RegFile.scala 76:16:@46769.4]
  assign regs_348_io_in = 64'h0; // @[RegFile.scala 75:16:@46768.4]
  assign regs_348_io_reset = reset; // @[RegFile.scala 78:19:@46772.4]
  assign regs_348_io_enable = 1'h1; // @[RegFile.scala 74:20:@46766.4]
  assign regs_349_clock = clock; // @[:@46775.4]
  assign regs_349_reset = io_reset; // @[:@46776.4 RegFile.scala 76:16:@46783.4]
  assign regs_349_io_in = 64'h0; // @[RegFile.scala 75:16:@46782.4]
  assign regs_349_io_reset = reset; // @[RegFile.scala 78:19:@46786.4]
  assign regs_349_io_enable = 1'h1; // @[RegFile.scala 74:20:@46780.4]
  assign regs_350_clock = clock; // @[:@46789.4]
  assign regs_350_reset = io_reset; // @[:@46790.4 RegFile.scala 76:16:@46797.4]
  assign regs_350_io_in = 64'h0; // @[RegFile.scala 75:16:@46796.4]
  assign regs_350_io_reset = reset; // @[RegFile.scala 78:19:@46800.4]
  assign regs_350_io_enable = 1'h1; // @[RegFile.scala 74:20:@46794.4]
  assign regs_351_clock = clock; // @[:@46803.4]
  assign regs_351_reset = io_reset; // @[:@46804.4 RegFile.scala 76:16:@46811.4]
  assign regs_351_io_in = 64'h0; // @[RegFile.scala 75:16:@46810.4]
  assign regs_351_io_reset = reset; // @[RegFile.scala 78:19:@46814.4]
  assign regs_351_io_enable = 1'h1; // @[RegFile.scala 74:20:@46808.4]
  assign regs_352_clock = clock; // @[:@46817.4]
  assign regs_352_reset = io_reset; // @[:@46818.4 RegFile.scala 76:16:@46825.4]
  assign regs_352_io_in = 64'h0; // @[RegFile.scala 75:16:@46824.4]
  assign regs_352_io_reset = reset; // @[RegFile.scala 78:19:@46828.4]
  assign regs_352_io_enable = 1'h1; // @[RegFile.scala 74:20:@46822.4]
  assign regs_353_clock = clock; // @[:@46831.4]
  assign regs_353_reset = io_reset; // @[:@46832.4 RegFile.scala 76:16:@46839.4]
  assign regs_353_io_in = 64'h0; // @[RegFile.scala 75:16:@46838.4]
  assign regs_353_io_reset = reset; // @[RegFile.scala 78:19:@46842.4]
  assign regs_353_io_enable = 1'h1; // @[RegFile.scala 74:20:@46836.4]
  assign regs_354_clock = clock; // @[:@46845.4]
  assign regs_354_reset = io_reset; // @[:@46846.4 RegFile.scala 76:16:@46853.4]
  assign regs_354_io_in = 64'h0; // @[RegFile.scala 75:16:@46852.4]
  assign regs_354_io_reset = reset; // @[RegFile.scala 78:19:@46856.4]
  assign regs_354_io_enable = 1'h1; // @[RegFile.scala 74:20:@46850.4]
  assign regs_355_clock = clock; // @[:@46859.4]
  assign regs_355_reset = io_reset; // @[:@46860.4 RegFile.scala 76:16:@46867.4]
  assign regs_355_io_in = 64'h0; // @[RegFile.scala 75:16:@46866.4]
  assign regs_355_io_reset = reset; // @[RegFile.scala 78:19:@46870.4]
  assign regs_355_io_enable = 1'h1; // @[RegFile.scala 74:20:@46864.4]
  assign regs_356_clock = clock; // @[:@46873.4]
  assign regs_356_reset = io_reset; // @[:@46874.4 RegFile.scala 76:16:@46881.4]
  assign regs_356_io_in = 64'h0; // @[RegFile.scala 75:16:@46880.4]
  assign regs_356_io_reset = reset; // @[RegFile.scala 78:19:@46884.4]
  assign regs_356_io_enable = 1'h1; // @[RegFile.scala 74:20:@46878.4]
  assign regs_357_clock = clock; // @[:@46887.4]
  assign regs_357_reset = io_reset; // @[:@46888.4 RegFile.scala 76:16:@46895.4]
  assign regs_357_io_in = 64'h0; // @[RegFile.scala 75:16:@46894.4]
  assign regs_357_io_reset = reset; // @[RegFile.scala 78:19:@46898.4]
  assign regs_357_io_enable = 1'h1; // @[RegFile.scala 74:20:@46892.4]
  assign regs_358_clock = clock; // @[:@46901.4]
  assign regs_358_reset = io_reset; // @[:@46902.4 RegFile.scala 76:16:@46909.4]
  assign regs_358_io_in = 64'h0; // @[RegFile.scala 75:16:@46908.4]
  assign regs_358_io_reset = reset; // @[RegFile.scala 78:19:@46912.4]
  assign regs_358_io_enable = 1'h1; // @[RegFile.scala 74:20:@46906.4]
  assign regs_359_clock = clock; // @[:@46915.4]
  assign regs_359_reset = io_reset; // @[:@46916.4 RegFile.scala 76:16:@46923.4]
  assign regs_359_io_in = 64'h0; // @[RegFile.scala 75:16:@46922.4]
  assign regs_359_io_reset = reset; // @[RegFile.scala 78:19:@46926.4]
  assign regs_359_io_enable = 1'h1; // @[RegFile.scala 74:20:@46920.4]
  assign regs_360_clock = clock; // @[:@46929.4]
  assign regs_360_reset = io_reset; // @[:@46930.4 RegFile.scala 76:16:@46937.4]
  assign regs_360_io_in = 64'h0; // @[RegFile.scala 75:16:@46936.4]
  assign regs_360_io_reset = reset; // @[RegFile.scala 78:19:@46940.4]
  assign regs_360_io_enable = 1'h1; // @[RegFile.scala 74:20:@46934.4]
  assign regs_361_clock = clock; // @[:@46943.4]
  assign regs_361_reset = io_reset; // @[:@46944.4 RegFile.scala 76:16:@46951.4]
  assign regs_361_io_in = 64'h0; // @[RegFile.scala 75:16:@46950.4]
  assign regs_361_io_reset = reset; // @[RegFile.scala 78:19:@46954.4]
  assign regs_361_io_enable = 1'h1; // @[RegFile.scala 74:20:@46948.4]
  assign regs_362_clock = clock; // @[:@46957.4]
  assign regs_362_reset = io_reset; // @[:@46958.4 RegFile.scala 76:16:@46965.4]
  assign regs_362_io_in = 64'h0; // @[RegFile.scala 75:16:@46964.4]
  assign regs_362_io_reset = reset; // @[RegFile.scala 78:19:@46968.4]
  assign regs_362_io_enable = 1'h1; // @[RegFile.scala 74:20:@46962.4]
  assign regs_363_clock = clock; // @[:@46971.4]
  assign regs_363_reset = io_reset; // @[:@46972.4 RegFile.scala 76:16:@46979.4]
  assign regs_363_io_in = 64'h0; // @[RegFile.scala 75:16:@46978.4]
  assign regs_363_io_reset = reset; // @[RegFile.scala 78:19:@46982.4]
  assign regs_363_io_enable = 1'h1; // @[RegFile.scala 74:20:@46976.4]
  assign regs_364_clock = clock; // @[:@46985.4]
  assign regs_364_reset = io_reset; // @[:@46986.4 RegFile.scala 76:16:@46993.4]
  assign regs_364_io_in = 64'h0; // @[RegFile.scala 75:16:@46992.4]
  assign regs_364_io_reset = reset; // @[RegFile.scala 78:19:@46996.4]
  assign regs_364_io_enable = 1'h1; // @[RegFile.scala 74:20:@46990.4]
  assign regs_365_clock = clock; // @[:@46999.4]
  assign regs_365_reset = io_reset; // @[:@47000.4 RegFile.scala 76:16:@47007.4]
  assign regs_365_io_in = 64'h0; // @[RegFile.scala 75:16:@47006.4]
  assign regs_365_io_reset = reset; // @[RegFile.scala 78:19:@47010.4]
  assign regs_365_io_enable = 1'h1; // @[RegFile.scala 74:20:@47004.4]
  assign regs_366_clock = clock; // @[:@47013.4]
  assign regs_366_reset = io_reset; // @[:@47014.4 RegFile.scala 76:16:@47021.4]
  assign regs_366_io_in = 64'h0; // @[RegFile.scala 75:16:@47020.4]
  assign regs_366_io_reset = reset; // @[RegFile.scala 78:19:@47024.4]
  assign regs_366_io_enable = 1'h1; // @[RegFile.scala 74:20:@47018.4]
  assign regs_367_clock = clock; // @[:@47027.4]
  assign regs_367_reset = io_reset; // @[:@47028.4 RegFile.scala 76:16:@47035.4]
  assign regs_367_io_in = 64'h0; // @[RegFile.scala 75:16:@47034.4]
  assign regs_367_io_reset = reset; // @[RegFile.scala 78:19:@47038.4]
  assign regs_367_io_enable = 1'h1; // @[RegFile.scala 74:20:@47032.4]
  assign regs_368_clock = clock; // @[:@47041.4]
  assign regs_368_reset = io_reset; // @[:@47042.4 RegFile.scala 76:16:@47049.4]
  assign regs_368_io_in = 64'h0; // @[RegFile.scala 75:16:@47048.4]
  assign regs_368_io_reset = reset; // @[RegFile.scala 78:19:@47052.4]
  assign regs_368_io_enable = 1'h1; // @[RegFile.scala 74:20:@47046.4]
  assign regs_369_clock = clock; // @[:@47055.4]
  assign regs_369_reset = io_reset; // @[:@47056.4 RegFile.scala 76:16:@47063.4]
  assign regs_369_io_in = 64'h0; // @[RegFile.scala 75:16:@47062.4]
  assign regs_369_io_reset = reset; // @[RegFile.scala 78:19:@47066.4]
  assign regs_369_io_enable = 1'h1; // @[RegFile.scala 74:20:@47060.4]
  assign regs_370_clock = clock; // @[:@47069.4]
  assign regs_370_reset = io_reset; // @[:@47070.4 RegFile.scala 76:16:@47077.4]
  assign regs_370_io_in = 64'h0; // @[RegFile.scala 75:16:@47076.4]
  assign regs_370_io_reset = reset; // @[RegFile.scala 78:19:@47080.4]
  assign regs_370_io_enable = 1'h1; // @[RegFile.scala 74:20:@47074.4]
  assign regs_371_clock = clock; // @[:@47083.4]
  assign regs_371_reset = io_reset; // @[:@47084.4 RegFile.scala 76:16:@47091.4]
  assign regs_371_io_in = 64'h0; // @[RegFile.scala 75:16:@47090.4]
  assign regs_371_io_reset = reset; // @[RegFile.scala 78:19:@47094.4]
  assign regs_371_io_enable = 1'h1; // @[RegFile.scala 74:20:@47088.4]
  assign regs_372_clock = clock; // @[:@47097.4]
  assign regs_372_reset = io_reset; // @[:@47098.4 RegFile.scala 76:16:@47105.4]
  assign regs_372_io_in = 64'h0; // @[RegFile.scala 75:16:@47104.4]
  assign regs_372_io_reset = reset; // @[RegFile.scala 78:19:@47108.4]
  assign regs_372_io_enable = 1'h1; // @[RegFile.scala 74:20:@47102.4]
  assign regs_373_clock = clock; // @[:@47111.4]
  assign regs_373_reset = io_reset; // @[:@47112.4 RegFile.scala 76:16:@47119.4]
  assign regs_373_io_in = 64'h0; // @[RegFile.scala 75:16:@47118.4]
  assign regs_373_io_reset = reset; // @[RegFile.scala 78:19:@47122.4]
  assign regs_373_io_enable = 1'h1; // @[RegFile.scala 74:20:@47116.4]
  assign regs_374_clock = clock; // @[:@47125.4]
  assign regs_374_reset = io_reset; // @[:@47126.4 RegFile.scala 76:16:@47133.4]
  assign regs_374_io_in = 64'h0; // @[RegFile.scala 75:16:@47132.4]
  assign regs_374_io_reset = reset; // @[RegFile.scala 78:19:@47136.4]
  assign regs_374_io_enable = 1'h1; // @[RegFile.scala 74:20:@47130.4]
  assign regs_375_clock = clock; // @[:@47139.4]
  assign regs_375_reset = io_reset; // @[:@47140.4 RegFile.scala 76:16:@47147.4]
  assign regs_375_io_in = 64'h0; // @[RegFile.scala 75:16:@47146.4]
  assign regs_375_io_reset = reset; // @[RegFile.scala 78:19:@47150.4]
  assign regs_375_io_enable = 1'h1; // @[RegFile.scala 74:20:@47144.4]
  assign regs_376_clock = clock; // @[:@47153.4]
  assign regs_376_reset = io_reset; // @[:@47154.4 RegFile.scala 76:16:@47161.4]
  assign regs_376_io_in = 64'h0; // @[RegFile.scala 75:16:@47160.4]
  assign regs_376_io_reset = reset; // @[RegFile.scala 78:19:@47164.4]
  assign regs_376_io_enable = 1'h1; // @[RegFile.scala 74:20:@47158.4]
  assign regs_377_clock = clock; // @[:@47167.4]
  assign regs_377_reset = io_reset; // @[:@47168.4 RegFile.scala 76:16:@47175.4]
  assign regs_377_io_in = 64'h0; // @[RegFile.scala 75:16:@47174.4]
  assign regs_377_io_reset = reset; // @[RegFile.scala 78:19:@47178.4]
  assign regs_377_io_enable = 1'h1; // @[RegFile.scala 74:20:@47172.4]
  assign regs_378_clock = clock; // @[:@47181.4]
  assign regs_378_reset = io_reset; // @[:@47182.4 RegFile.scala 76:16:@47189.4]
  assign regs_378_io_in = 64'h0; // @[RegFile.scala 75:16:@47188.4]
  assign regs_378_io_reset = reset; // @[RegFile.scala 78:19:@47192.4]
  assign regs_378_io_enable = 1'h1; // @[RegFile.scala 74:20:@47186.4]
  assign regs_379_clock = clock; // @[:@47195.4]
  assign regs_379_reset = io_reset; // @[:@47196.4 RegFile.scala 76:16:@47203.4]
  assign regs_379_io_in = 64'h0; // @[RegFile.scala 75:16:@47202.4]
  assign regs_379_io_reset = reset; // @[RegFile.scala 78:19:@47206.4]
  assign regs_379_io_enable = 1'h1; // @[RegFile.scala 74:20:@47200.4]
  assign regs_380_clock = clock; // @[:@47209.4]
  assign regs_380_reset = io_reset; // @[:@47210.4 RegFile.scala 76:16:@47217.4]
  assign regs_380_io_in = 64'h0; // @[RegFile.scala 75:16:@47216.4]
  assign regs_380_io_reset = reset; // @[RegFile.scala 78:19:@47220.4]
  assign regs_380_io_enable = 1'h1; // @[RegFile.scala 74:20:@47214.4]
  assign regs_381_clock = clock; // @[:@47223.4]
  assign regs_381_reset = io_reset; // @[:@47224.4 RegFile.scala 76:16:@47231.4]
  assign regs_381_io_in = 64'h0; // @[RegFile.scala 75:16:@47230.4]
  assign regs_381_io_reset = reset; // @[RegFile.scala 78:19:@47234.4]
  assign regs_381_io_enable = 1'h1; // @[RegFile.scala 74:20:@47228.4]
  assign regs_382_clock = clock; // @[:@47237.4]
  assign regs_382_reset = io_reset; // @[:@47238.4 RegFile.scala 76:16:@47245.4]
  assign regs_382_io_in = 64'h0; // @[RegFile.scala 75:16:@47244.4]
  assign regs_382_io_reset = reset; // @[RegFile.scala 78:19:@47248.4]
  assign regs_382_io_enable = 1'h1; // @[RegFile.scala 74:20:@47242.4]
  assign regs_383_clock = clock; // @[:@47251.4]
  assign regs_383_reset = io_reset; // @[:@47252.4 RegFile.scala 76:16:@47259.4]
  assign regs_383_io_in = 64'h0; // @[RegFile.scala 75:16:@47258.4]
  assign regs_383_io_reset = reset; // @[RegFile.scala 78:19:@47262.4]
  assign regs_383_io_enable = 1'h1; // @[RegFile.scala 74:20:@47256.4]
  assign regs_384_clock = clock; // @[:@47265.4]
  assign regs_384_reset = io_reset; // @[:@47266.4 RegFile.scala 76:16:@47273.4]
  assign regs_384_io_in = 64'h0; // @[RegFile.scala 75:16:@47272.4]
  assign regs_384_io_reset = reset; // @[RegFile.scala 78:19:@47276.4]
  assign regs_384_io_enable = 1'h1; // @[RegFile.scala 74:20:@47270.4]
  assign regs_385_clock = clock; // @[:@47279.4]
  assign regs_385_reset = io_reset; // @[:@47280.4 RegFile.scala 76:16:@47287.4]
  assign regs_385_io_in = 64'h0; // @[RegFile.scala 75:16:@47286.4]
  assign regs_385_io_reset = reset; // @[RegFile.scala 78:19:@47290.4]
  assign regs_385_io_enable = 1'h1; // @[RegFile.scala 74:20:@47284.4]
  assign regs_386_clock = clock; // @[:@47293.4]
  assign regs_386_reset = io_reset; // @[:@47294.4 RegFile.scala 76:16:@47301.4]
  assign regs_386_io_in = 64'h0; // @[RegFile.scala 75:16:@47300.4]
  assign regs_386_io_reset = reset; // @[RegFile.scala 78:19:@47304.4]
  assign regs_386_io_enable = 1'h1; // @[RegFile.scala 74:20:@47298.4]
  assign regs_387_clock = clock; // @[:@47307.4]
  assign regs_387_reset = io_reset; // @[:@47308.4 RegFile.scala 76:16:@47315.4]
  assign regs_387_io_in = 64'h0; // @[RegFile.scala 75:16:@47314.4]
  assign regs_387_io_reset = reset; // @[RegFile.scala 78:19:@47318.4]
  assign regs_387_io_enable = 1'h1; // @[RegFile.scala 74:20:@47312.4]
  assign regs_388_clock = clock; // @[:@47321.4]
  assign regs_388_reset = io_reset; // @[:@47322.4 RegFile.scala 76:16:@47329.4]
  assign regs_388_io_in = 64'h0; // @[RegFile.scala 75:16:@47328.4]
  assign regs_388_io_reset = reset; // @[RegFile.scala 78:19:@47332.4]
  assign regs_388_io_enable = 1'h1; // @[RegFile.scala 74:20:@47326.4]
  assign regs_389_clock = clock; // @[:@47335.4]
  assign regs_389_reset = io_reset; // @[:@47336.4 RegFile.scala 76:16:@47343.4]
  assign regs_389_io_in = 64'h0; // @[RegFile.scala 75:16:@47342.4]
  assign regs_389_io_reset = reset; // @[RegFile.scala 78:19:@47346.4]
  assign regs_389_io_enable = 1'h1; // @[RegFile.scala 74:20:@47340.4]
  assign regs_390_clock = clock; // @[:@47349.4]
  assign regs_390_reset = io_reset; // @[:@47350.4 RegFile.scala 76:16:@47357.4]
  assign regs_390_io_in = 64'h0; // @[RegFile.scala 75:16:@47356.4]
  assign regs_390_io_reset = reset; // @[RegFile.scala 78:19:@47360.4]
  assign regs_390_io_enable = 1'h1; // @[RegFile.scala 74:20:@47354.4]
  assign regs_391_clock = clock; // @[:@47363.4]
  assign regs_391_reset = io_reset; // @[:@47364.4 RegFile.scala 76:16:@47371.4]
  assign regs_391_io_in = 64'h0; // @[RegFile.scala 75:16:@47370.4]
  assign regs_391_io_reset = reset; // @[RegFile.scala 78:19:@47374.4]
  assign regs_391_io_enable = 1'h1; // @[RegFile.scala 74:20:@47368.4]
  assign regs_392_clock = clock; // @[:@47377.4]
  assign regs_392_reset = io_reset; // @[:@47378.4 RegFile.scala 76:16:@47385.4]
  assign regs_392_io_in = 64'h0; // @[RegFile.scala 75:16:@47384.4]
  assign regs_392_io_reset = reset; // @[RegFile.scala 78:19:@47388.4]
  assign regs_392_io_enable = 1'h1; // @[RegFile.scala 74:20:@47382.4]
  assign regs_393_clock = clock; // @[:@47391.4]
  assign regs_393_reset = io_reset; // @[:@47392.4 RegFile.scala 76:16:@47399.4]
  assign regs_393_io_in = 64'h0; // @[RegFile.scala 75:16:@47398.4]
  assign regs_393_io_reset = reset; // @[RegFile.scala 78:19:@47402.4]
  assign regs_393_io_enable = 1'h1; // @[RegFile.scala 74:20:@47396.4]
  assign regs_394_clock = clock; // @[:@47405.4]
  assign regs_394_reset = io_reset; // @[:@47406.4 RegFile.scala 76:16:@47413.4]
  assign regs_394_io_in = 64'h0; // @[RegFile.scala 75:16:@47412.4]
  assign regs_394_io_reset = reset; // @[RegFile.scala 78:19:@47416.4]
  assign regs_394_io_enable = 1'h1; // @[RegFile.scala 74:20:@47410.4]
  assign regs_395_clock = clock; // @[:@47419.4]
  assign regs_395_reset = io_reset; // @[:@47420.4 RegFile.scala 76:16:@47427.4]
  assign regs_395_io_in = 64'h0; // @[RegFile.scala 75:16:@47426.4]
  assign regs_395_io_reset = reset; // @[RegFile.scala 78:19:@47430.4]
  assign regs_395_io_enable = 1'h1; // @[RegFile.scala 74:20:@47424.4]
  assign regs_396_clock = clock; // @[:@47433.4]
  assign regs_396_reset = io_reset; // @[:@47434.4 RegFile.scala 76:16:@47441.4]
  assign regs_396_io_in = 64'h0; // @[RegFile.scala 75:16:@47440.4]
  assign regs_396_io_reset = reset; // @[RegFile.scala 78:19:@47444.4]
  assign regs_396_io_enable = 1'h1; // @[RegFile.scala 74:20:@47438.4]
  assign regs_397_clock = clock; // @[:@47447.4]
  assign regs_397_reset = io_reset; // @[:@47448.4 RegFile.scala 76:16:@47455.4]
  assign regs_397_io_in = 64'h0; // @[RegFile.scala 75:16:@47454.4]
  assign regs_397_io_reset = reset; // @[RegFile.scala 78:19:@47458.4]
  assign regs_397_io_enable = 1'h1; // @[RegFile.scala 74:20:@47452.4]
  assign regs_398_clock = clock; // @[:@47461.4]
  assign regs_398_reset = io_reset; // @[:@47462.4 RegFile.scala 76:16:@47469.4]
  assign regs_398_io_in = 64'h0; // @[RegFile.scala 75:16:@47468.4]
  assign regs_398_io_reset = reset; // @[RegFile.scala 78:19:@47472.4]
  assign regs_398_io_enable = 1'h1; // @[RegFile.scala 74:20:@47466.4]
  assign regs_399_clock = clock; // @[:@47475.4]
  assign regs_399_reset = io_reset; // @[:@47476.4 RegFile.scala 76:16:@47483.4]
  assign regs_399_io_in = 64'h0; // @[RegFile.scala 75:16:@47482.4]
  assign regs_399_io_reset = reset; // @[RegFile.scala 78:19:@47486.4]
  assign regs_399_io_enable = 1'h1; // @[RegFile.scala 74:20:@47480.4]
  assign regs_400_clock = clock; // @[:@47489.4]
  assign regs_400_reset = io_reset; // @[:@47490.4 RegFile.scala 76:16:@47497.4]
  assign regs_400_io_in = 64'h0; // @[RegFile.scala 75:16:@47496.4]
  assign regs_400_io_reset = reset; // @[RegFile.scala 78:19:@47500.4]
  assign regs_400_io_enable = 1'h1; // @[RegFile.scala 74:20:@47494.4]
  assign regs_401_clock = clock; // @[:@47503.4]
  assign regs_401_reset = io_reset; // @[:@47504.4 RegFile.scala 76:16:@47511.4]
  assign regs_401_io_in = 64'h0; // @[RegFile.scala 75:16:@47510.4]
  assign regs_401_io_reset = reset; // @[RegFile.scala 78:19:@47514.4]
  assign regs_401_io_enable = 1'h1; // @[RegFile.scala 74:20:@47508.4]
  assign regs_402_clock = clock; // @[:@47517.4]
  assign regs_402_reset = io_reset; // @[:@47518.4 RegFile.scala 76:16:@47525.4]
  assign regs_402_io_in = 64'h0; // @[RegFile.scala 75:16:@47524.4]
  assign regs_402_io_reset = reset; // @[RegFile.scala 78:19:@47528.4]
  assign regs_402_io_enable = 1'h1; // @[RegFile.scala 74:20:@47522.4]
  assign regs_403_clock = clock; // @[:@47531.4]
  assign regs_403_reset = io_reset; // @[:@47532.4 RegFile.scala 76:16:@47539.4]
  assign regs_403_io_in = 64'h0; // @[RegFile.scala 75:16:@47538.4]
  assign regs_403_io_reset = reset; // @[RegFile.scala 78:19:@47542.4]
  assign regs_403_io_enable = 1'h1; // @[RegFile.scala 74:20:@47536.4]
  assign regs_404_clock = clock; // @[:@47545.4]
  assign regs_404_reset = io_reset; // @[:@47546.4 RegFile.scala 76:16:@47553.4]
  assign regs_404_io_in = 64'h0; // @[RegFile.scala 75:16:@47552.4]
  assign regs_404_io_reset = reset; // @[RegFile.scala 78:19:@47556.4]
  assign regs_404_io_enable = 1'h1; // @[RegFile.scala 74:20:@47550.4]
  assign regs_405_clock = clock; // @[:@47559.4]
  assign regs_405_reset = io_reset; // @[:@47560.4 RegFile.scala 76:16:@47567.4]
  assign regs_405_io_in = 64'h0; // @[RegFile.scala 75:16:@47566.4]
  assign regs_405_io_reset = reset; // @[RegFile.scala 78:19:@47570.4]
  assign regs_405_io_enable = 1'h1; // @[RegFile.scala 74:20:@47564.4]
  assign regs_406_clock = clock; // @[:@47573.4]
  assign regs_406_reset = io_reset; // @[:@47574.4 RegFile.scala 76:16:@47581.4]
  assign regs_406_io_in = 64'h0; // @[RegFile.scala 75:16:@47580.4]
  assign regs_406_io_reset = reset; // @[RegFile.scala 78:19:@47584.4]
  assign regs_406_io_enable = 1'h1; // @[RegFile.scala 74:20:@47578.4]
  assign regs_407_clock = clock; // @[:@47587.4]
  assign regs_407_reset = io_reset; // @[:@47588.4 RegFile.scala 76:16:@47595.4]
  assign regs_407_io_in = 64'h0; // @[RegFile.scala 75:16:@47594.4]
  assign regs_407_io_reset = reset; // @[RegFile.scala 78:19:@47598.4]
  assign regs_407_io_enable = 1'h1; // @[RegFile.scala 74:20:@47592.4]
  assign regs_408_clock = clock; // @[:@47601.4]
  assign regs_408_reset = io_reset; // @[:@47602.4 RegFile.scala 76:16:@47609.4]
  assign regs_408_io_in = 64'h0; // @[RegFile.scala 75:16:@47608.4]
  assign regs_408_io_reset = reset; // @[RegFile.scala 78:19:@47612.4]
  assign regs_408_io_enable = 1'h1; // @[RegFile.scala 74:20:@47606.4]
  assign regs_409_clock = clock; // @[:@47615.4]
  assign regs_409_reset = io_reset; // @[:@47616.4 RegFile.scala 76:16:@47623.4]
  assign regs_409_io_in = 64'h0; // @[RegFile.scala 75:16:@47622.4]
  assign regs_409_io_reset = reset; // @[RegFile.scala 78:19:@47626.4]
  assign regs_409_io_enable = 1'h1; // @[RegFile.scala 74:20:@47620.4]
  assign regs_410_clock = clock; // @[:@47629.4]
  assign regs_410_reset = io_reset; // @[:@47630.4 RegFile.scala 76:16:@47637.4]
  assign regs_410_io_in = 64'h0; // @[RegFile.scala 75:16:@47636.4]
  assign regs_410_io_reset = reset; // @[RegFile.scala 78:19:@47640.4]
  assign regs_410_io_enable = 1'h1; // @[RegFile.scala 74:20:@47634.4]
  assign regs_411_clock = clock; // @[:@47643.4]
  assign regs_411_reset = io_reset; // @[:@47644.4 RegFile.scala 76:16:@47651.4]
  assign regs_411_io_in = 64'h0; // @[RegFile.scala 75:16:@47650.4]
  assign regs_411_io_reset = reset; // @[RegFile.scala 78:19:@47654.4]
  assign regs_411_io_enable = 1'h1; // @[RegFile.scala 74:20:@47648.4]
  assign regs_412_clock = clock; // @[:@47657.4]
  assign regs_412_reset = io_reset; // @[:@47658.4 RegFile.scala 76:16:@47665.4]
  assign regs_412_io_in = 64'h0; // @[RegFile.scala 75:16:@47664.4]
  assign regs_412_io_reset = reset; // @[RegFile.scala 78:19:@47668.4]
  assign regs_412_io_enable = 1'h1; // @[RegFile.scala 74:20:@47662.4]
  assign regs_413_clock = clock; // @[:@47671.4]
  assign regs_413_reset = io_reset; // @[:@47672.4 RegFile.scala 76:16:@47679.4]
  assign regs_413_io_in = 64'h0; // @[RegFile.scala 75:16:@47678.4]
  assign regs_413_io_reset = reset; // @[RegFile.scala 78:19:@47682.4]
  assign regs_413_io_enable = 1'h1; // @[RegFile.scala 74:20:@47676.4]
  assign regs_414_clock = clock; // @[:@47685.4]
  assign regs_414_reset = io_reset; // @[:@47686.4 RegFile.scala 76:16:@47693.4]
  assign regs_414_io_in = 64'h0; // @[RegFile.scala 75:16:@47692.4]
  assign regs_414_io_reset = reset; // @[RegFile.scala 78:19:@47696.4]
  assign regs_414_io_enable = 1'h1; // @[RegFile.scala 74:20:@47690.4]
  assign regs_415_clock = clock; // @[:@47699.4]
  assign regs_415_reset = io_reset; // @[:@47700.4 RegFile.scala 76:16:@47707.4]
  assign regs_415_io_in = 64'h0; // @[RegFile.scala 75:16:@47706.4]
  assign regs_415_io_reset = reset; // @[RegFile.scala 78:19:@47710.4]
  assign regs_415_io_enable = 1'h1; // @[RegFile.scala 74:20:@47704.4]
  assign regs_416_clock = clock; // @[:@47713.4]
  assign regs_416_reset = io_reset; // @[:@47714.4 RegFile.scala 76:16:@47721.4]
  assign regs_416_io_in = 64'h0; // @[RegFile.scala 75:16:@47720.4]
  assign regs_416_io_reset = reset; // @[RegFile.scala 78:19:@47724.4]
  assign regs_416_io_enable = 1'h1; // @[RegFile.scala 74:20:@47718.4]
  assign regs_417_clock = clock; // @[:@47727.4]
  assign regs_417_reset = io_reset; // @[:@47728.4 RegFile.scala 76:16:@47735.4]
  assign regs_417_io_in = 64'h0; // @[RegFile.scala 75:16:@47734.4]
  assign regs_417_io_reset = reset; // @[RegFile.scala 78:19:@47738.4]
  assign regs_417_io_enable = 1'h1; // @[RegFile.scala 74:20:@47732.4]
  assign regs_418_clock = clock; // @[:@47741.4]
  assign regs_418_reset = io_reset; // @[:@47742.4 RegFile.scala 76:16:@47749.4]
  assign regs_418_io_in = 64'h0; // @[RegFile.scala 75:16:@47748.4]
  assign regs_418_io_reset = reset; // @[RegFile.scala 78:19:@47752.4]
  assign regs_418_io_enable = 1'h1; // @[RegFile.scala 74:20:@47746.4]
  assign regs_419_clock = clock; // @[:@47755.4]
  assign regs_419_reset = io_reset; // @[:@47756.4 RegFile.scala 76:16:@47763.4]
  assign regs_419_io_in = 64'h0; // @[RegFile.scala 75:16:@47762.4]
  assign regs_419_io_reset = reset; // @[RegFile.scala 78:19:@47766.4]
  assign regs_419_io_enable = 1'h1; // @[RegFile.scala 74:20:@47760.4]
  assign regs_420_clock = clock; // @[:@47769.4]
  assign regs_420_reset = io_reset; // @[:@47770.4 RegFile.scala 76:16:@47777.4]
  assign regs_420_io_in = 64'h0; // @[RegFile.scala 75:16:@47776.4]
  assign regs_420_io_reset = reset; // @[RegFile.scala 78:19:@47780.4]
  assign regs_420_io_enable = 1'h1; // @[RegFile.scala 74:20:@47774.4]
  assign regs_421_clock = clock; // @[:@47783.4]
  assign regs_421_reset = io_reset; // @[:@47784.4 RegFile.scala 76:16:@47791.4]
  assign regs_421_io_in = 64'h0; // @[RegFile.scala 75:16:@47790.4]
  assign regs_421_io_reset = reset; // @[RegFile.scala 78:19:@47794.4]
  assign regs_421_io_enable = 1'h1; // @[RegFile.scala 74:20:@47788.4]
  assign regs_422_clock = clock; // @[:@47797.4]
  assign regs_422_reset = io_reset; // @[:@47798.4 RegFile.scala 76:16:@47805.4]
  assign regs_422_io_in = 64'h0; // @[RegFile.scala 75:16:@47804.4]
  assign regs_422_io_reset = reset; // @[RegFile.scala 78:19:@47808.4]
  assign regs_422_io_enable = 1'h1; // @[RegFile.scala 74:20:@47802.4]
  assign regs_423_clock = clock; // @[:@47811.4]
  assign regs_423_reset = io_reset; // @[:@47812.4 RegFile.scala 76:16:@47819.4]
  assign regs_423_io_in = 64'h0; // @[RegFile.scala 75:16:@47818.4]
  assign regs_423_io_reset = reset; // @[RegFile.scala 78:19:@47822.4]
  assign regs_423_io_enable = 1'h1; // @[RegFile.scala 74:20:@47816.4]
  assign regs_424_clock = clock; // @[:@47825.4]
  assign regs_424_reset = io_reset; // @[:@47826.4 RegFile.scala 76:16:@47833.4]
  assign regs_424_io_in = 64'h0; // @[RegFile.scala 75:16:@47832.4]
  assign regs_424_io_reset = reset; // @[RegFile.scala 78:19:@47836.4]
  assign regs_424_io_enable = 1'h1; // @[RegFile.scala 74:20:@47830.4]
  assign regs_425_clock = clock; // @[:@47839.4]
  assign regs_425_reset = io_reset; // @[:@47840.4 RegFile.scala 76:16:@47847.4]
  assign regs_425_io_in = 64'h0; // @[RegFile.scala 75:16:@47846.4]
  assign regs_425_io_reset = reset; // @[RegFile.scala 78:19:@47850.4]
  assign regs_425_io_enable = 1'h1; // @[RegFile.scala 74:20:@47844.4]
  assign regs_426_clock = clock; // @[:@47853.4]
  assign regs_426_reset = io_reset; // @[:@47854.4 RegFile.scala 76:16:@47861.4]
  assign regs_426_io_in = 64'h0; // @[RegFile.scala 75:16:@47860.4]
  assign regs_426_io_reset = reset; // @[RegFile.scala 78:19:@47864.4]
  assign regs_426_io_enable = 1'h1; // @[RegFile.scala 74:20:@47858.4]
  assign regs_427_clock = clock; // @[:@47867.4]
  assign regs_427_reset = io_reset; // @[:@47868.4 RegFile.scala 76:16:@47875.4]
  assign regs_427_io_in = 64'h0; // @[RegFile.scala 75:16:@47874.4]
  assign regs_427_io_reset = reset; // @[RegFile.scala 78:19:@47878.4]
  assign regs_427_io_enable = 1'h1; // @[RegFile.scala 74:20:@47872.4]
  assign regs_428_clock = clock; // @[:@47881.4]
  assign regs_428_reset = io_reset; // @[:@47882.4 RegFile.scala 76:16:@47889.4]
  assign regs_428_io_in = 64'h0; // @[RegFile.scala 75:16:@47888.4]
  assign regs_428_io_reset = reset; // @[RegFile.scala 78:19:@47892.4]
  assign regs_428_io_enable = 1'h1; // @[RegFile.scala 74:20:@47886.4]
  assign regs_429_clock = clock; // @[:@47895.4]
  assign regs_429_reset = io_reset; // @[:@47896.4 RegFile.scala 76:16:@47903.4]
  assign regs_429_io_in = 64'h0; // @[RegFile.scala 75:16:@47902.4]
  assign regs_429_io_reset = reset; // @[RegFile.scala 78:19:@47906.4]
  assign regs_429_io_enable = 1'h1; // @[RegFile.scala 74:20:@47900.4]
  assign regs_430_clock = clock; // @[:@47909.4]
  assign regs_430_reset = io_reset; // @[:@47910.4 RegFile.scala 76:16:@47917.4]
  assign regs_430_io_in = 64'h0; // @[RegFile.scala 75:16:@47916.4]
  assign regs_430_io_reset = reset; // @[RegFile.scala 78:19:@47920.4]
  assign regs_430_io_enable = 1'h1; // @[RegFile.scala 74:20:@47914.4]
  assign regs_431_clock = clock; // @[:@47923.4]
  assign regs_431_reset = io_reset; // @[:@47924.4 RegFile.scala 76:16:@47931.4]
  assign regs_431_io_in = 64'h0; // @[RegFile.scala 75:16:@47930.4]
  assign regs_431_io_reset = reset; // @[RegFile.scala 78:19:@47934.4]
  assign regs_431_io_enable = 1'h1; // @[RegFile.scala 74:20:@47928.4]
  assign regs_432_clock = clock; // @[:@47937.4]
  assign regs_432_reset = io_reset; // @[:@47938.4 RegFile.scala 76:16:@47945.4]
  assign regs_432_io_in = 64'h0; // @[RegFile.scala 75:16:@47944.4]
  assign regs_432_io_reset = reset; // @[RegFile.scala 78:19:@47948.4]
  assign regs_432_io_enable = 1'h1; // @[RegFile.scala 74:20:@47942.4]
  assign regs_433_clock = clock; // @[:@47951.4]
  assign regs_433_reset = io_reset; // @[:@47952.4 RegFile.scala 76:16:@47959.4]
  assign regs_433_io_in = 64'h0; // @[RegFile.scala 75:16:@47958.4]
  assign regs_433_io_reset = reset; // @[RegFile.scala 78:19:@47962.4]
  assign regs_433_io_enable = 1'h1; // @[RegFile.scala 74:20:@47956.4]
  assign regs_434_clock = clock; // @[:@47965.4]
  assign regs_434_reset = io_reset; // @[:@47966.4 RegFile.scala 76:16:@47973.4]
  assign regs_434_io_in = 64'h0; // @[RegFile.scala 75:16:@47972.4]
  assign regs_434_io_reset = reset; // @[RegFile.scala 78:19:@47976.4]
  assign regs_434_io_enable = 1'h1; // @[RegFile.scala 74:20:@47970.4]
  assign regs_435_clock = clock; // @[:@47979.4]
  assign regs_435_reset = io_reset; // @[:@47980.4 RegFile.scala 76:16:@47987.4]
  assign regs_435_io_in = 64'h0; // @[RegFile.scala 75:16:@47986.4]
  assign regs_435_io_reset = reset; // @[RegFile.scala 78:19:@47990.4]
  assign regs_435_io_enable = 1'h1; // @[RegFile.scala 74:20:@47984.4]
  assign regs_436_clock = clock; // @[:@47993.4]
  assign regs_436_reset = io_reset; // @[:@47994.4 RegFile.scala 76:16:@48001.4]
  assign regs_436_io_in = 64'h0; // @[RegFile.scala 75:16:@48000.4]
  assign regs_436_io_reset = reset; // @[RegFile.scala 78:19:@48004.4]
  assign regs_436_io_enable = 1'h1; // @[RegFile.scala 74:20:@47998.4]
  assign regs_437_clock = clock; // @[:@48007.4]
  assign regs_437_reset = io_reset; // @[:@48008.4 RegFile.scala 76:16:@48015.4]
  assign regs_437_io_in = 64'h0; // @[RegFile.scala 75:16:@48014.4]
  assign regs_437_io_reset = reset; // @[RegFile.scala 78:19:@48018.4]
  assign regs_437_io_enable = 1'h1; // @[RegFile.scala 74:20:@48012.4]
  assign regs_438_clock = clock; // @[:@48021.4]
  assign regs_438_reset = io_reset; // @[:@48022.4 RegFile.scala 76:16:@48029.4]
  assign regs_438_io_in = 64'h0; // @[RegFile.scala 75:16:@48028.4]
  assign regs_438_io_reset = reset; // @[RegFile.scala 78:19:@48032.4]
  assign regs_438_io_enable = 1'h1; // @[RegFile.scala 74:20:@48026.4]
  assign regs_439_clock = clock; // @[:@48035.4]
  assign regs_439_reset = io_reset; // @[:@48036.4 RegFile.scala 76:16:@48043.4]
  assign regs_439_io_in = 64'h0; // @[RegFile.scala 75:16:@48042.4]
  assign regs_439_io_reset = reset; // @[RegFile.scala 78:19:@48046.4]
  assign regs_439_io_enable = 1'h1; // @[RegFile.scala 74:20:@48040.4]
  assign regs_440_clock = clock; // @[:@48049.4]
  assign regs_440_reset = io_reset; // @[:@48050.4 RegFile.scala 76:16:@48057.4]
  assign regs_440_io_in = 64'h0; // @[RegFile.scala 75:16:@48056.4]
  assign regs_440_io_reset = reset; // @[RegFile.scala 78:19:@48060.4]
  assign regs_440_io_enable = 1'h1; // @[RegFile.scala 74:20:@48054.4]
  assign regs_441_clock = clock; // @[:@48063.4]
  assign regs_441_reset = io_reset; // @[:@48064.4 RegFile.scala 76:16:@48071.4]
  assign regs_441_io_in = 64'h0; // @[RegFile.scala 75:16:@48070.4]
  assign regs_441_io_reset = reset; // @[RegFile.scala 78:19:@48074.4]
  assign regs_441_io_enable = 1'h1; // @[RegFile.scala 74:20:@48068.4]
  assign regs_442_clock = clock; // @[:@48077.4]
  assign regs_442_reset = io_reset; // @[:@48078.4 RegFile.scala 76:16:@48085.4]
  assign regs_442_io_in = 64'h0; // @[RegFile.scala 75:16:@48084.4]
  assign regs_442_io_reset = reset; // @[RegFile.scala 78:19:@48088.4]
  assign regs_442_io_enable = 1'h1; // @[RegFile.scala 74:20:@48082.4]
  assign regs_443_clock = clock; // @[:@48091.4]
  assign regs_443_reset = io_reset; // @[:@48092.4 RegFile.scala 76:16:@48099.4]
  assign regs_443_io_in = 64'h0; // @[RegFile.scala 75:16:@48098.4]
  assign regs_443_io_reset = reset; // @[RegFile.scala 78:19:@48102.4]
  assign regs_443_io_enable = 1'h1; // @[RegFile.scala 74:20:@48096.4]
  assign regs_444_clock = clock; // @[:@48105.4]
  assign regs_444_reset = io_reset; // @[:@48106.4 RegFile.scala 76:16:@48113.4]
  assign regs_444_io_in = 64'h0; // @[RegFile.scala 75:16:@48112.4]
  assign regs_444_io_reset = reset; // @[RegFile.scala 78:19:@48116.4]
  assign regs_444_io_enable = 1'h1; // @[RegFile.scala 74:20:@48110.4]
  assign regs_445_clock = clock; // @[:@48119.4]
  assign regs_445_reset = io_reset; // @[:@48120.4 RegFile.scala 76:16:@48127.4]
  assign regs_445_io_in = 64'h0; // @[RegFile.scala 75:16:@48126.4]
  assign regs_445_io_reset = reset; // @[RegFile.scala 78:19:@48130.4]
  assign regs_445_io_enable = 1'h1; // @[RegFile.scala 74:20:@48124.4]
  assign regs_446_clock = clock; // @[:@48133.4]
  assign regs_446_reset = io_reset; // @[:@48134.4 RegFile.scala 76:16:@48141.4]
  assign regs_446_io_in = 64'h0; // @[RegFile.scala 75:16:@48140.4]
  assign regs_446_io_reset = reset; // @[RegFile.scala 78:19:@48144.4]
  assign regs_446_io_enable = 1'h1; // @[RegFile.scala 74:20:@48138.4]
  assign regs_447_clock = clock; // @[:@48147.4]
  assign regs_447_reset = io_reset; // @[:@48148.4 RegFile.scala 76:16:@48155.4]
  assign regs_447_io_in = 64'h0; // @[RegFile.scala 75:16:@48154.4]
  assign regs_447_io_reset = reset; // @[RegFile.scala 78:19:@48158.4]
  assign regs_447_io_enable = 1'h1; // @[RegFile.scala 74:20:@48152.4]
  assign regs_448_clock = clock; // @[:@48161.4]
  assign regs_448_reset = io_reset; // @[:@48162.4 RegFile.scala 76:16:@48169.4]
  assign regs_448_io_in = 64'h0; // @[RegFile.scala 75:16:@48168.4]
  assign regs_448_io_reset = reset; // @[RegFile.scala 78:19:@48172.4]
  assign regs_448_io_enable = 1'h1; // @[RegFile.scala 74:20:@48166.4]
  assign regs_449_clock = clock; // @[:@48175.4]
  assign regs_449_reset = io_reset; // @[:@48176.4 RegFile.scala 76:16:@48183.4]
  assign regs_449_io_in = 64'h0; // @[RegFile.scala 75:16:@48182.4]
  assign regs_449_io_reset = reset; // @[RegFile.scala 78:19:@48186.4]
  assign regs_449_io_enable = 1'h1; // @[RegFile.scala 74:20:@48180.4]
  assign regs_450_clock = clock; // @[:@48189.4]
  assign regs_450_reset = io_reset; // @[:@48190.4 RegFile.scala 76:16:@48197.4]
  assign regs_450_io_in = 64'h0; // @[RegFile.scala 75:16:@48196.4]
  assign regs_450_io_reset = reset; // @[RegFile.scala 78:19:@48200.4]
  assign regs_450_io_enable = 1'h1; // @[RegFile.scala 74:20:@48194.4]
  assign regs_451_clock = clock; // @[:@48203.4]
  assign regs_451_reset = io_reset; // @[:@48204.4 RegFile.scala 76:16:@48211.4]
  assign regs_451_io_in = 64'h0; // @[RegFile.scala 75:16:@48210.4]
  assign regs_451_io_reset = reset; // @[RegFile.scala 78:19:@48214.4]
  assign regs_451_io_enable = 1'h1; // @[RegFile.scala 74:20:@48208.4]
  assign regs_452_clock = clock; // @[:@48217.4]
  assign regs_452_reset = io_reset; // @[:@48218.4 RegFile.scala 76:16:@48225.4]
  assign regs_452_io_in = 64'h0; // @[RegFile.scala 75:16:@48224.4]
  assign regs_452_io_reset = reset; // @[RegFile.scala 78:19:@48228.4]
  assign regs_452_io_enable = 1'h1; // @[RegFile.scala 74:20:@48222.4]
  assign regs_453_clock = clock; // @[:@48231.4]
  assign regs_453_reset = io_reset; // @[:@48232.4 RegFile.scala 76:16:@48239.4]
  assign regs_453_io_in = 64'h0; // @[RegFile.scala 75:16:@48238.4]
  assign regs_453_io_reset = reset; // @[RegFile.scala 78:19:@48242.4]
  assign regs_453_io_enable = 1'h1; // @[RegFile.scala 74:20:@48236.4]
  assign regs_454_clock = clock; // @[:@48245.4]
  assign regs_454_reset = io_reset; // @[:@48246.4 RegFile.scala 76:16:@48253.4]
  assign regs_454_io_in = 64'h0; // @[RegFile.scala 75:16:@48252.4]
  assign regs_454_io_reset = reset; // @[RegFile.scala 78:19:@48256.4]
  assign regs_454_io_enable = 1'h1; // @[RegFile.scala 74:20:@48250.4]
  assign regs_455_clock = clock; // @[:@48259.4]
  assign regs_455_reset = io_reset; // @[:@48260.4 RegFile.scala 76:16:@48267.4]
  assign regs_455_io_in = 64'h0; // @[RegFile.scala 75:16:@48266.4]
  assign regs_455_io_reset = reset; // @[RegFile.scala 78:19:@48270.4]
  assign regs_455_io_enable = 1'h1; // @[RegFile.scala 74:20:@48264.4]
  assign regs_456_clock = clock; // @[:@48273.4]
  assign regs_456_reset = io_reset; // @[:@48274.4 RegFile.scala 76:16:@48281.4]
  assign regs_456_io_in = 64'h0; // @[RegFile.scala 75:16:@48280.4]
  assign regs_456_io_reset = reset; // @[RegFile.scala 78:19:@48284.4]
  assign regs_456_io_enable = 1'h1; // @[RegFile.scala 74:20:@48278.4]
  assign regs_457_clock = clock; // @[:@48287.4]
  assign regs_457_reset = io_reset; // @[:@48288.4 RegFile.scala 76:16:@48295.4]
  assign regs_457_io_in = 64'h0; // @[RegFile.scala 75:16:@48294.4]
  assign regs_457_io_reset = reset; // @[RegFile.scala 78:19:@48298.4]
  assign regs_457_io_enable = 1'h1; // @[RegFile.scala 74:20:@48292.4]
  assign regs_458_clock = clock; // @[:@48301.4]
  assign regs_458_reset = io_reset; // @[:@48302.4 RegFile.scala 76:16:@48309.4]
  assign regs_458_io_in = 64'h0; // @[RegFile.scala 75:16:@48308.4]
  assign regs_458_io_reset = reset; // @[RegFile.scala 78:19:@48312.4]
  assign regs_458_io_enable = 1'h1; // @[RegFile.scala 74:20:@48306.4]
  assign regs_459_clock = clock; // @[:@48315.4]
  assign regs_459_reset = io_reset; // @[:@48316.4 RegFile.scala 76:16:@48323.4]
  assign regs_459_io_in = 64'h0; // @[RegFile.scala 75:16:@48322.4]
  assign regs_459_io_reset = reset; // @[RegFile.scala 78:19:@48326.4]
  assign regs_459_io_enable = 1'h1; // @[RegFile.scala 74:20:@48320.4]
  assign regs_460_clock = clock; // @[:@48329.4]
  assign regs_460_reset = io_reset; // @[:@48330.4 RegFile.scala 76:16:@48337.4]
  assign regs_460_io_in = 64'h0; // @[RegFile.scala 75:16:@48336.4]
  assign regs_460_io_reset = reset; // @[RegFile.scala 78:19:@48340.4]
  assign regs_460_io_enable = 1'h1; // @[RegFile.scala 74:20:@48334.4]
  assign regs_461_clock = clock; // @[:@48343.4]
  assign regs_461_reset = io_reset; // @[:@48344.4 RegFile.scala 76:16:@48351.4]
  assign regs_461_io_in = 64'h0; // @[RegFile.scala 75:16:@48350.4]
  assign regs_461_io_reset = reset; // @[RegFile.scala 78:19:@48354.4]
  assign regs_461_io_enable = 1'h1; // @[RegFile.scala 74:20:@48348.4]
  assign regs_462_clock = clock; // @[:@48357.4]
  assign regs_462_reset = io_reset; // @[:@48358.4 RegFile.scala 76:16:@48365.4]
  assign regs_462_io_in = 64'h0; // @[RegFile.scala 75:16:@48364.4]
  assign regs_462_io_reset = reset; // @[RegFile.scala 78:19:@48368.4]
  assign regs_462_io_enable = 1'h1; // @[RegFile.scala 74:20:@48362.4]
  assign regs_463_clock = clock; // @[:@48371.4]
  assign regs_463_reset = io_reset; // @[:@48372.4 RegFile.scala 76:16:@48379.4]
  assign regs_463_io_in = 64'h0; // @[RegFile.scala 75:16:@48378.4]
  assign regs_463_io_reset = reset; // @[RegFile.scala 78:19:@48382.4]
  assign regs_463_io_enable = 1'h1; // @[RegFile.scala 74:20:@48376.4]
  assign regs_464_clock = clock; // @[:@48385.4]
  assign regs_464_reset = io_reset; // @[:@48386.4 RegFile.scala 76:16:@48393.4]
  assign regs_464_io_in = 64'h0; // @[RegFile.scala 75:16:@48392.4]
  assign regs_464_io_reset = reset; // @[RegFile.scala 78:19:@48396.4]
  assign regs_464_io_enable = 1'h1; // @[RegFile.scala 74:20:@48390.4]
  assign regs_465_clock = clock; // @[:@48399.4]
  assign regs_465_reset = io_reset; // @[:@48400.4 RegFile.scala 76:16:@48407.4]
  assign regs_465_io_in = 64'h0; // @[RegFile.scala 75:16:@48406.4]
  assign regs_465_io_reset = reset; // @[RegFile.scala 78:19:@48410.4]
  assign regs_465_io_enable = 1'h1; // @[RegFile.scala 74:20:@48404.4]
  assign regs_466_clock = clock; // @[:@48413.4]
  assign regs_466_reset = io_reset; // @[:@48414.4 RegFile.scala 76:16:@48421.4]
  assign regs_466_io_in = 64'h0; // @[RegFile.scala 75:16:@48420.4]
  assign regs_466_io_reset = reset; // @[RegFile.scala 78:19:@48424.4]
  assign regs_466_io_enable = 1'h1; // @[RegFile.scala 74:20:@48418.4]
  assign regs_467_clock = clock; // @[:@48427.4]
  assign regs_467_reset = io_reset; // @[:@48428.4 RegFile.scala 76:16:@48435.4]
  assign regs_467_io_in = 64'h0; // @[RegFile.scala 75:16:@48434.4]
  assign regs_467_io_reset = reset; // @[RegFile.scala 78:19:@48438.4]
  assign regs_467_io_enable = 1'h1; // @[RegFile.scala 74:20:@48432.4]
  assign regs_468_clock = clock; // @[:@48441.4]
  assign regs_468_reset = io_reset; // @[:@48442.4 RegFile.scala 76:16:@48449.4]
  assign regs_468_io_in = 64'h0; // @[RegFile.scala 75:16:@48448.4]
  assign regs_468_io_reset = reset; // @[RegFile.scala 78:19:@48452.4]
  assign regs_468_io_enable = 1'h1; // @[RegFile.scala 74:20:@48446.4]
  assign regs_469_clock = clock; // @[:@48455.4]
  assign regs_469_reset = io_reset; // @[:@48456.4 RegFile.scala 76:16:@48463.4]
  assign regs_469_io_in = 64'h0; // @[RegFile.scala 75:16:@48462.4]
  assign regs_469_io_reset = reset; // @[RegFile.scala 78:19:@48466.4]
  assign regs_469_io_enable = 1'h1; // @[RegFile.scala 74:20:@48460.4]
  assign regs_470_clock = clock; // @[:@48469.4]
  assign regs_470_reset = io_reset; // @[:@48470.4 RegFile.scala 76:16:@48477.4]
  assign regs_470_io_in = 64'h0; // @[RegFile.scala 75:16:@48476.4]
  assign regs_470_io_reset = reset; // @[RegFile.scala 78:19:@48480.4]
  assign regs_470_io_enable = 1'h1; // @[RegFile.scala 74:20:@48474.4]
  assign regs_471_clock = clock; // @[:@48483.4]
  assign regs_471_reset = io_reset; // @[:@48484.4 RegFile.scala 76:16:@48491.4]
  assign regs_471_io_in = 64'h0; // @[RegFile.scala 75:16:@48490.4]
  assign regs_471_io_reset = reset; // @[RegFile.scala 78:19:@48494.4]
  assign regs_471_io_enable = 1'h1; // @[RegFile.scala 74:20:@48488.4]
  assign regs_472_clock = clock; // @[:@48497.4]
  assign regs_472_reset = io_reset; // @[:@48498.4 RegFile.scala 76:16:@48505.4]
  assign regs_472_io_in = 64'h0; // @[RegFile.scala 75:16:@48504.4]
  assign regs_472_io_reset = reset; // @[RegFile.scala 78:19:@48508.4]
  assign regs_472_io_enable = 1'h1; // @[RegFile.scala 74:20:@48502.4]
  assign regs_473_clock = clock; // @[:@48511.4]
  assign regs_473_reset = io_reset; // @[:@48512.4 RegFile.scala 76:16:@48519.4]
  assign regs_473_io_in = 64'h0; // @[RegFile.scala 75:16:@48518.4]
  assign regs_473_io_reset = reset; // @[RegFile.scala 78:19:@48522.4]
  assign regs_473_io_enable = 1'h1; // @[RegFile.scala 74:20:@48516.4]
  assign regs_474_clock = clock; // @[:@48525.4]
  assign regs_474_reset = io_reset; // @[:@48526.4 RegFile.scala 76:16:@48533.4]
  assign regs_474_io_in = 64'h0; // @[RegFile.scala 75:16:@48532.4]
  assign regs_474_io_reset = reset; // @[RegFile.scala 78:19:@48536.4]
  assign regs_474_io_enable = 1'h1; // @[RegFile.scala 74:20:@48530.4]
  assign regs_475_clock = clock; // @[:@48539.4]
  assign regs_475_reset = io_reset; // @[:@48540.4 RegFile.scala 76:16:@48547.4]
  assign regs_475_io_in = 64'h0; // @[RegFile.scala 75:16:@48546.4]
  assign regs_475_io_reset = reset; // @[RegFile.scala 78:19:@48550.4]
  assign regs_475_io_enable = 1'h1; // @[RegFile.scala 74:20:@48544.4]
  assign regs_476_clock = clock; // @[:@48553.4]
  assign regs_476_reset = io_reset; // @[:@48554.4 RegFile.scala 76:16:@48561.4]
  assign regs_476_io_in = 64'h0; // @[RegFile.scala 75:16:@48560.4]
  assign regs_476_io_reset = reset; // @[RegFile.scala 78:19:@48564.4]
  assign regs_476_io_enable = 1'h1; // @[RegFile.scala 74:20:@48558.4]
  assign regs_477_clock = clock; // @[:@48567.4]
  assign regs_477_reset = io_reset; // @[:@48568.4 RegFile.scala 76:16:@48575.4]
  assign regs_477_io_in = 64'h0; // @[RegFile.scala 75:16:@48574.4]
  assign regs_477_io_reset = reset; // @[RegFile.scala 78:19:@48578.4]
  assign regs_477_io_enable = 1'h1; // @[RegFile.scala 74:20:@48572.4]
  assign regs_478_clock = clock; // @[:@48581.4]
  assign regs_478_reset = io_reset; // @[:@48582.4 RegFile.scala 76:16:@48589.4]
  assign regs_478_io_in = 64'h0; // @[RegFile.scala 75:16:@48588.4]
  assign regs_478_io_reset = reset; // @[RegFile.scala 78:19:@48592.4]
  assign regs_478_io_enable = 1'h1; // @[RegFile.scala 74:20:@48586.4]
  assign regs_479_clock = clock; // @[:@48595.4]
  assign regs_479_reset = io_reset; // @[:@48596.4 RegFile.scala 76:16:@48603.4]
  assign regs_479_io_in = 64'h0; // @[RegFile.scala 75:16:@48602.4]
  assign regs_479_io_reset = reset; // @[RegFile.scala 78:19:@48606.4]
  assign regs_479_io_enable = 1'h1; // @[RegFile.scala 74:20:@48600.4]
  assign regs_480_clock = clock; // @[:@48609.4]
  assign regs_480_reset = io_reset; // @[:@48610.4 RegFile.scala 76:16:@48617.4]
  assign regs_480_io_in = 64'h0; // @[RegFile.scala 75:16:@48616.4]
  assign regs_480_io_reset = reset; // @[RegFile.scala 78:19:@48620.4]
  assign regs_480_io_enable = 1'h1; // @[RegFile.scala 74:20:@48614.4]
  assign regs_481_clock = clock; // @[:@48623.4]
  assign regs_481_reset = io_reset; // @[:@48624.4 RegFile.scala 76:16:@48631.4]
  assign regs_481_io_in = 64'h0; // @[RegFile.scala 75:16:@48630.4]
  assign regs_481_io_reset = reset; // @[RegFile.scala 78:19:@48634.4]
  assign regs_481_io_enable = 1'h1; // @[RegFile.scala 74:20:@48628.4]
  assign regs_482_clock = clock; // @[:@48637.4]
  assign regs_482_reset = io_reset; // @[:@48638.4 RegFile.scala 76:16:@48645.4]
  assign regs_482_io_in = 64'h0; // @[RegFile.scala 75:16:@48644.4]
  assign regs_482_io_reset = reset; // @[RegFile.scala 78:19:@48648.4]
  assign regs_482_io_enable = 1'h1; // @[RegFile.scala 74:20:@48642.4]
  assign regs_483_clock = clock; // @[:@48651.4]
  assign regs_483_reset = io_reset; // @[:@48652.4 RegFile.scala 76:16:@48659.4]
  assign regs_483_io_in = 64'h0; // @[RegFile.scala 75:16:@48658.4]
  assign regs_483_io_reset = reset; // @[RegFile.scala 78:19:@48662.4]
  assign regs_483_io_enable = 1'h1; // @[RegFile.scala 74:20:@48656.4]
  assign regs_484_clock = clock; // @[:@48665.4]
  assign regs_484_reset = io_reset; // @[:@48666.4 RegFile.scala 76:16:@48673.4]
  assign regs_484_io_in = 64'h0; // @[RegFile.scala 75:16:@48672.4]
  assign regs_484_io_reset = reset; // @[RegFile.scala 78:19:@48676.4]
  assign regs_484_io_enable = 1'h1; // @[RegFile.scala 74:20:@48670.4]
  assign regs_485_clock = clock; // @[:@48679.4]
  assign regs_485_reset = io_reset; // @[:@48680.4 RegFile.scala 76:16:@48687.4]
  assign regs_485_io_in = 64'h0; // @[RegFile.scala 75:16:@48686.4]
  assign regs_485_io_reset = reset; // @[RegFile.scala 78:19:@48690.4]
  assign regs_485_io_enable = 1'h1; // @[RegFile.scala 74:20:@48684.4]
  assign regs_486_clock = clock; // @[:@48693.4]
  assign regs_486_reset = io_reset; // @[:@48694.4 RegFile.scala 76:16:@48701.4]
  assign regs_486_io_in = 64'h0; // @[RegFile.scala 75:16:@48700.4]
  assign regs_486_io_reset = reset; // @[RegFile.scala 78:19:@48704.4]
  assign regs_486_io_enable = 1'h1; // @[RegFile.scala 74:20:@48698.4]
  assign regs_487_clock = clock; // @[:@48707.4]
  assign regs_487_reset = io_reset; // @[:@48708.4 RegFile.scala 76:16:@48715.4]
  assign regs_487_io_in = 64'h0; // @[RegFile.scala 75:16:@48714.4]
  assign regs_487_io_reset = reset; // @[RegFile.scala 78:19:@48718.4]
  assign regs_487_io_enable = 1'h1; // @[RegFile.scala 74:20:@48712.4]
  assign regs_488_clock = clock; // @[:@48721.4]
  assign regs_488_reset = io_reset; // @[:@48722.4 RegFile.scala 76:16:@48729.4]
  assign regs_488_io_in = 64'h0; // @[RegFile.scala 75:16:@48728.4]
  assign regs_488_io_reset = reset; // @[RegFile.scala 78:19:@48732.4]
  assign regs_488_io_enable = 1'h1; // @[RegFile.scala 74:20:@48726.4]
  assign regs_489_clock = clock; // @[:@48735.4]
  assign regs_489_reset = io_reset; // @[:@48736.4 RegFile.scala 76:16:@48743.4]
  assign regs_489_io_in = 64'h0; // @[RegFile.scala 75:16:@48742.4]
  assign regs_489_io_reset = reset; // @[RegFile.scala 78:19:@48746.4]
  assign regs_489_io_enable = 1'h1; // @[RegFile.scala 74:20:@48740.4]
  assign regs_490_clock = clock; // @[:@48749.4]
  assign regs_490_reset = io_reset; // @[:@48750.4 RegFile.scala 76:16:@48757.4]
  assign regs_490_io_in = 64'h0; // @[RegFile.scala 75:16:@48756.4]
  assign regs_490_io_reset = reset; // @[RegFile.scala 78:19:@48760.4]
  assign regs_490_io_enable = 1'h1; // @[RegFile.scala 74:20:@48754.4]
  assign regs_491_clock = clock; // @[:@48763.4]
  assign regs_491_reset = io_reset; // @[:@48764.4 RegFile.scala 76:16:@48771.4]
  assign regs_491_io_in = 64'h0; // @[RegFile.scala 75:16:@48770.4]
  assign regs_491_io_reset = reset; // @[RegFile.scala 78:19:@48774.4]
  assign regs_491_io_enable = 1'h1; // @[RegFile.scala 74:20:@48768.4]
  assign regs_492_clock = clock; // @[:@48777.4]
  assign regs_492_reset = io_reset; // @[:@48778.4 RegFile.scala 76:16:@48785.4]
  assign regs_492_io_in = 64'h0; // @[RegFile.scala 75:16:@48784.4]
  assign regs_492_io_reset = reset; // @[RegFile.scala 78:19:@48788.4]
  assign regs_492_io_enable = 1'h1; // @[RegFile.scala 74:20:@48782.4]
  assign regs_493_clock = clock; // @[:@48791.4]
  assign regs_493_reset = io_reset; // @[:@48792.4 RegFile.scala 76:16:@48799.4]
  assign regs_493_io_in = 64'h0; // @[RegFile.scala 75:16:@48798.4]
  assign regs_493_io_reset = reset; // @[RegFile.scala 78:19:@48802.4]
  assign regs_493_io_enable = 1'h1; // @[RegFile.scala 74:20:@48796.4]
  assign regs_494_clock = clock; // @[:@48805.4]
  assign regs_494_reset = io_reset; // @[:@48806.4 RegFile.scala 76:16:@48813.4]
  assign regs_494_io_in = 64'h0; // @[RegFile.scala 75:16:@48812.4]
  assign regs_494_io_reset = reset; // @[RegFile.scala 78:19:@48816.4]
  assign regs_494_io_enable = 1'h1; // @[RegFile.scala 74:20:@48810.4]
  assign regs_495_clock = clock; // @[:@48819.4]
  assign regs_495_reset = io_reset; // @[:@48820.4 RegFile.scala 76:16:@48827.4]
  assign regs_495_io_in = 64'h0; // @[RegFile.scala 75:16:@48826.4]
  assign regs_495_io_reset = reset; // @[RegFile.scala 78:19:@48830.4]
  assign regs_495_io_enable = 1'h1; // @[RegFile.scala 74:20:@48824.4]
  assign regs_496_clock = clock; // @[:@48833.4]
  assign regs_496_reset = io_reset; // @[:@48834.4 RegFile.scala 76:16:@48841.4]
  assign regs_496_io_in = 64'h0; // @[RegFile.scala 75:16:@48840.4]
  assign regs_496_io_reset = reset; // @[RegFile.scala 78:19:@48844.4]
  assign regs_496_io_enable = 1'h1; // @[RegFile.scala 74:20:@48838.4]
  assign regs_497_clock = clock; // @[:@48847.4]
  assign regs_497_reset = io_reset; // @[:@48848.4 RegFile.scala 76:16:@48855.4]
  assign regs_497_io_in = 64'h0; // @[RegFile.scala 75:16:@48854.4]
  assign regs_497_io_reset = reset; // @[RegFile.scala 78:19:@48858.4]
  assign regs_497_io_enable = 1'h1; // @[RegFile.scala 74:20:@48852.4]
  assign regs_498_clock = clock; // @[:@48861.4]
  assign regs_498_reset = io_reset; // @[:@48862.4 RegFile.scala 76:16:@48869.4]
  assign regs_498_io_in = 64'h0; // @[RegFile.scala 75:16:@48868.4]
  assign regs_498_io_reset = reset; // @[RegFile.scala 78:19:@48872.4]
  assign regs_498_io_enable = 1'h1; // @[RegFile.scala 74:20:@48866.4]
  assign regs_499_clock = clock; // @[:@48875.4]
  assign regs_499_reset = io_reset; // @[:@48876.4 RegFile.scala 76:16:@48883.4]
  assign regs_499_io_in = 64'h0; // @[RegFile.scala 75:16:@48882.4]
  assign regs_499_io_reset = reset; // @[RegFile.scala 78:19:@48886.4]
  assign regs_499_io_enable = 1'h1; // @[RegFile.scala 74:20:@48880.4]
  assign regs_500_clock = clock; // @[:@48889.4]
  assign regs_500_reset = io_reset; // @[:@48890.4 RegFile.scala 76:16:@48897.4]
  assign regs_500_io_in = 64'h0; // @[RegFile.scala 75:16:@48896.4]
  assign regs_500_io_reset = reset; // @[RegFile.scala 78:19:@48900.4]
  assign regs_500_io_enable = 1'h1; // @[RegFile.scala 74:20:@48894.4]
  assign regs_501_clock = clock; // @[:@48903.4]
  assign regs_501_reset = io_reset; // @[:@48904.4 RegFile.scala 76:16:@48911.4]
  assign regs_501_io_in = 64'h0; // @[RegFile.scala 75:16:@48910.4]
  assign regs_501_io_reset = reset; // @[RegFile.scala 78:19:@48914.4]
  assign regs_501_io_enable = 1'h1; // @[RegFile.scala 74:20:@48908.4]
  assign regs_502_clock = clock; // @[:@48917.4]
  assign regs_502_reset = io_reset; // @[:@48918.4 RegFile.scala 76:16:@48925.4]
  assign regs_502_io_in = 64'h0; // @[RegFile.scala 75:16:@48924.4]
  assign regs_502_io_reset = reset; // @[RegFile.scala 78:19:@48928.4]
  assign regs_502_io_enable = 1'h1; // @[RegFile.scala 74:20:@48922.4]
  assign regs_503_clock = clock; // @[:@48931.4]
  assign regs_503_reset = io_reset; // @[:@48932.4 RegFile.scala 76:16:@48939.4]
  assign regs_503_io_in = 64'h0; // @[RegFile.scala 75:16:@48938.4]
  assign regs_503_io_reset = reset; // @[RegFile.scala 78:19:@48942.4]
  assign regs_503_io_enable = 1'h1; // @[RegFile.scala 74:20:@48936.4]
  assign regs_504_clock = clock; // @[:@48945.4]
  assign regs_504_reset = io_reset; // @[:@48946.4 RegFile.scala 76:16:@48953.4]
  assign regs_504_io_in = 64'h0; // @[RegFile.scala 75:16:@48952.4]
  assign regs_504_io_reset = reset; // @[RegFile.scala 78:19:@48956.4]
  assign regs_504_io_enable = 1'h1; // @[RegFile.scala 74:20:@48950.4]
  assign regs_505_clock = clock; // @[:@48959.4]
  assign regs_505_reset = io_reset; // @[:@48960.4 RegFile.scala 76:16:@48967.4]
  assign regs_505_io_in = 64'h0; // @[RegFile.scala 75:16:@48966.4]
  assign regs_505_io_reset = reset; // @[RegFile.scala 78:19:@48970.4]
  assign regs_505_io_enable = 1'h1; // @[RegFile.scala 74:20:@48964.4]
  assign regs_506_clock = clock; // @[:@48973.4]
  assign regs_506_reset = io_reset; // @[:@48974.4 RegFile.scala 76:16:@48981.4]
  assign regs_506_io_in = 64'h0; // @[RegFile.scala 75:16:@48980.4]
  assign regs_506_io_reset = reset; // @[RegFile.scala 78:19:@48984.4]
  assign regs_506_io_enable = 1'h1; // @[RegFile.scala 74:20:@48978.4]
  assign regs_507_clock = clock; // @[:@48987.4]
  assign regs_507_reset = io_reset; // @[:@48988.4 RegFile.scala 76:16:@48995.4]
  assign regs_507_io_in = 64'h0; // @[RegFile.scala 75:16:@48994.4]
  assign regs_507_io_reset = reset; // @[RegFile.scala 78:19:@48998.4]
  assign regs_507_io_enable = 1'h1; // @[RegFile.scala 74:20:@48992.4]
  assign regs_508_clock = clock; // @[:@49001.4]
  assign regs_508_reset = io_reset; // @[:@49002.4 RegFile.scala 76:16:@49009.4]
  assign regs_508_io_in = 64'h0; // @[RegFile.scala 75:16:@49008.4]
  assign regs_508_io_reset = reset; // @[RegFile.scala 78:19:@49012.4]
  assign regs_508_io_enable = 1'h1; // @[RegFile.scala 74:20:@49006.4]
  assign regs_509_clock = clock; // @[:@49015.4]
  assign regs_509_reset = io_reset; // @[:@49016.4 RegFile.scala 76:16:@49023.4]
  assign regs_509_io_in = 64'h0; // @[RegFile.scala 75:16:@49022.4]
  assign regs_509_io_reset = reset; // @[RegFile.scala 78:19:@49026.4]
  assign regs_509_io_enable = 1'h1; // @[RegFile.scala 74:20:@49020.4]
  assign regs_510_clock = clock; // @[:@49029.4]
  assign regs_510_reset = io_reset; // @[:@49030.4 RegFile.scala 76:16:@49037.4]
  assign regs_510_io_in = 64'h0; // @[RegFile.scala 75:16:@49036.4]
  assign regs_510_io_reset = reset; // @[RegFile.scala 78:19:@49040.4]
  assign regs_510_io_enable = 1'h1; // @[RegFile.scala 74:20:@49034.4]
  assign regs_511_clock = clock; // @[:@49043.4]
  assign regs_511_reset = io_reset; // @[:@49044.4 RegFile.scala 76:16:@49051.4]
  assign regs_511_io_in = 64'h0; // @[RegFile.scala 75:16:@49050.4]
  assign regs_511_io_reset = reset; // @[RegFile.scala 78:19:@49054.4]
  assign regs_511_io_enable = 1'h1; // @[RegFile.scala 74:20:@49048.4]
  assign regs_512_clock = clock; // @[:@49057.4]
  assign regs_512_reset = io_reset; // @[:@49058.4 RegFile.scala 76:16:@49065.4]
  assign regs_512_io_in = 64'h0; // @[RegFile.scala 75:16:@49064.4]
  assign regs_512_io_reset = reset; // @[RegFile.scala 78:19:@49068.4]
  assign regs_512_io_enable = 1'h1; // @[RegFile.scala 74:20:@49062.4]
  assign regs_513_clock = clock; // @[:@49071.4]
  assign regs_513_reset = io_reset; // @[:@49072.4 RegFile.scala 76:16:@49079.4]
  assign regs_513_io_in = 64'h0; // @[RegFile.scala 75:16:@49078.4]
  assign regs_513_io_reset = reset; // @[RegFile.scala 78:19:@49082.4]
  assign regs_513_io_enable = 1'h1; // @[RegFile.scala 74:20:@49076.4]
  assign regs_514_clock = clock; // @[:@49085.4]
  assign regs_514_reset = io_reset; // @[:@49086.4 RegFile.scala 76:16:@49093.4]
  assign regs_514_io_in = 64'h0; // @[RegFile.scala 75:16:@49092.4]
  assign regs_514_io_reset = reset; // @[RegFile.scala 78:19:@49096.4]
  assign regs_514_io_enable = 1'h1; // @[RegFile.scala 74:20:@49090.4]
  assign regs_515_clock = clock; // @[:@49099.4]
  assign regs_515_reset = io_reset; // @[:@49100.4 RegFile.scala 76:16:@49107.4]
  assign regs_515_io_in = 64'h0; // @[RegFile.scala 75:16:@49106.4]
  assign regs_515_io_reset = reset; // @[RegFile.scala 78:19:@49110.4]
  assign regs_515_io_enable = 1'h1; // @[RegFile.scala 74:20:@49104.4]
  assign regs_516_clock = clock; // @[:@49113.4]
  assign regs_516_reset = io_reset; // @[:@49114.4 RegFile.scala 76:16:@49121.4]
  assign regs_516_io_in = 64'h0; // @[RegFile.scala 75:16:@49120.4]
  assign regs_516_io_reset = reset; // @[RegFile.scala 78:19:@49124.4]
  assign regs_516_io_enable = 1'h1; // @[RegFile.scala 74:20:@49118.4]
  assign regs_517_clock = clock; // @[:@49127.4]
  assign regs_517_reset = io_reset; // @[:@49128.4 RegFile.scala 76:16:@49135.4]
  assign regs_517_io_in = 64'h0; // @[RegFile.scala 75:16:@49134.4]
  assign regs_517_io_reset = reset; // @[RegFile.scala 78:19:@49138.4]
  assign regs_517_io_enable = 1'h1; // @[RegFile.scala 74:20:@49132.4]
  assign regs_518_clock = clock; // @[:@49141.4]
  assign regs_518_reset = io_reset; // @[:@49142.4 RegFile.scala 76:16:@49149.4]
  assign regs_518_io_in = 64'h0; // @[RegFile.scala 75:16:@49148.4]
  assign regs_518_io_reset = reset; // @[RegFile.scala 78:19:@49152.4]
  assign regs_518_io_enable = 1'h1; // @[RegFile.scala 74:20:@49146.4]
  assign regs_519_clock = clock; // @[:@49155.4]
  assign regs_519_reset = io_reset; // @[:@49156.4 RegFile.scala 76:16:@49163.4]
  assign regs_519_io_in = 64'h0; // @[RegFile.scala 75:16:@49162.4]
  assign regs_519_io_reset = reset; // @[RegFile.scala 78:19:@49166.4]
  assign regs_519_io_enable = 1'h1; // @[RegFile.scala 74:20:@49160.4]
  assign regs_520_clock = clock; // @[:@49169.4]
  assign regs_520_reset = io_reset; // @[:@49170.4 RegFile.scala 76:16:@49177.4]
  assign regs_520_io_in = 64'h0; // @[RegFile.scala 75:16:@49176.4]
  assign regs_520_io_reset = reset; // @[RegFile.scala 78:19:@49180.4]
  assign regs_520_io_enable = 1'h1; // @[RegFile.scala 74:20:@49174.4]
  assign regs_521_clock = clock; // @[:@49183.4]
  assign regs_521_reset = io_reset; // @[:@49184.4 RegFile.scala 76:16:@49191.4]
  assign regs_521_io_in = 64'h0; // @[RegFile.scala 75:16:@49190.4]
  assign regs_521_io_reset = reset; // @[RegFile.scala 78:19:@49194.4]
  assign regs_521_io_enable = 1'h1; // @[RegFile.scala 74:20:@49188.4]
  assign rport_io_ins_0 = regs_0_io_out; // @[RegFile.scala 97:16:@49722.4]
  assign rport_io_ins_1 = regs_1_io_out; // @[RegFile.scala 97:16:@49723.4]
  assign rport_io_ins_2 = regs_2_io_out; // @[RegFile.scala 97:16:@49724.4]
  assign rport_io_ins_3 = regs_3_io_out; // @[RegFile.scala 97:16:@49725.4]
  assign rport_io_ins_4 = regs_4_io_out; // @[RegFile.scala 97:16:@49726.4]
  assign rport_io_ins_5 = regs_5_io_out; // @[RegFile.scala 97:16:@49727.4]
  assign rport_io_ins_6 = regs_6_io_out; // @[RegFile.scala 97:16:@49728.4]
  assign rport_io_ins_7 = regs_7_io_out; // @[RegFile.scala 97:16:@49729.4]
  assign rport_io_ins_8 = regs_8_io_out; // @[RegFile.scala 97:16:@49730.4]
  assign rport_io_ins_9 = regs_9_io_out; // @[RegFile.scala 97:16:@49731.4]
  assign rport_io_ins_10 = regs_10_io_out; // @[RegFile.scala 97:16:@49732.4]
  assign rport_io_ins_11 = regs_11_io_out; // @[RegFile.scala 97:16:@49733.4]
  assign rport_io_ins_12 = regs_12_io_out; // @[RegFile.scala 97:16:@49734.4]
  assign rport_io_ins_13 = regs_13_io_out; // @[RegFile.scala 97:16:@49735.4]
  assign rport_io_ins_14 = regs_14_io_out; // @[RegFile.scala 97:16:@49736.4]
  assign rport_io_ins_15 = regs_15_io_out; // @[RegFile.scala 97:16:@49737.4]
  assign rport_io_ins_16 = regs_16_io_out; // @[RegFile.scala 97:16:@49738.4]
  assign rport_io_ins_17 = regs_17_io_out; // @[RegFile.scala 97:16:@49739.4]
  assign rport_io_ins_18 = regs_18_io_out; // @[RegFile.scala 97:16:@49740.4]
  assign rport_io_ins_19 = regs_19_io_out; // @[RegFile.scala 97:16:@49741.4]
  assign rport_io_ins_20 = regs_20_io_out; // @[RegFile.scala 97:16:@49742.4]
  assign rport_io_ins_21 = regs_21_io_out; // @[RegFile.scala 97:16:@49743.4]
  assign rport_io_ins_22 = regs_22_io_out; // @[RegFile.scala 97:16:@49744.4]
  assign rport_io_ins_23 = regs_23_io_out; // @[RegFile.scala 97:16:@49745.4]
  assign rport_io_ins_24 = regs_24_io_out; // @[RegFile.scala 97:16:@49746.4]
  assign rport_io_ins_25 = regs_25_io_out; // @[RegFile.scala 97:16:@49747.4]
  assign rport_io_ins_26 = regs_26_io_out; // @[RegFile.scala 97:16:@49748.4]
  assign rport_io_ins_27 = regs_27_io_out; // @[RegFile.scala 97:16:@49749.4]
  assign rport_io_ins_28 = regs_28_io_out; // @[RegFile.scala 97:16:@49750.4]
  assign rport_io_ins_29 = regs_29_io_out; // @[RegFile.scala 97:16:@49751.4]
  assign rport_io_ins_30 = regs_30_io_out; // @[RegFile.scala 97:16:@49752.4]
  assign rport_io_ins_31 = regs_31_io_out; // @[RegFile.scala 97:16:@49753.4]
  assign rport_io_ins_32 = regs_32_io_out; // @[RegFile.scala 97:16:@49754.4]
  assign rport_io_ins_33 = regs_33_io_out; // @[RegFile.scala 97:16:@49755.4]
  assign rport_io_ins_34 = regs_34_io_out; // @[RegFile.scala 97:16:@49756.4]
  assign rport_io_ins_35 = regs_35_io_out; // @[RegFile.scala 97:16:@49757.4]
  assign rport_io_ins_36 = regs_36_io_out; // @[RegFile.scala 97:16:@49758.4]
  assign rport_io_ins_37 = regs_37_io_out; // @[RegFile.scala 97:16:@49759.4]
  assign rport_io_ins_38 = regs_38_io_out; // @[RegFile.scala 97:16:@49760.4]
  assign rport_io_ins_39 = regs_39_io_out; // @[RegFile.scala 97:16:@49761.4]
  assign rport_io_ins_40 = regs_40_io_out; // @[RegFile.scala 97:16:@49762.4]
  assign rport_io_ins_41 = regs_41_io_out; // @[RegFile.scala 97:16:@49763.4]
  assign rport_io_ins_42 = regs_42_io_out; // @[RegFile.scala 97:16:@49764.4]
  assign rport_io_ins_43 = regs_43_io_out; // @[RegFile.scala 97:16:@49765.4]
  assign rport_io_ins_44 = regs_44_io_out; // @[RegFile.scala 97:16:@49766.4]
  assign rport_io_ins_45 = regs_45_io_out; // @[RegFile.scala 97:16:@49767.4]
  assign rport_io_ins_46 = regs_46_io_out; // @[RegFile.scala 97:16:@49768.4]
  assign rport_io_ins_47 = regs_47_io_out; // @[RegFile.scala 97:16:@49769.4]
  assign rport_io_ins_48 = regs_48_io_out; // @[RegFile.scala 97:16:@49770.4]
  assign rport_io_ins_49 = regs_49_io_out; // @[RegFile.scala 97:16:@49771.4]
  assign rport_io_ins_50 = regs_50_io_out; // @[RegFile.scala 97:16:@49772.4]
  assign rport_io_ins_51 = regs_51_io_out; // @[RegFile.scala 97:16:@49773.4]
  assign rport_io_ins_52 = regs_52_io_out; // @[RegFile.scala 97:16:@49774.4]
  assign rport_io_ins_53 = regs_53_io_out; // @[RegFile.scala 97:16:@49775.4]
  assign rport_io_ins_54 = regs_54_io_out; // @[RegFile.scala 97:16:@49776.4]
  assign rport_io_ins_55 = regs_55_io_out; // @[RegFile.scala 97:16:@49777.4]
  assign rport_io_ins_56 = regs_56_io_out; // @[RegFile.scala 97:16:@49778.4]
  assign rport_io_ins_57 = regs_57_io_out; // @[RegFile.scala 97:16:@49779.4]
  assign rport_io_ins_58 = regs_58_io_out; // @[RegFile.scala 97:16:@49780.4]
  assign rport_io_ins_59 = regs_59_io_out; // @[RegFile.scala 97:16:@49781.4]
  assign rport_io_ins_60 = regs_60_io_out; // @[RegFile.scala 97:16:@49782.4]
  assign rport_io_ins_61 = regs_61_io_out; // @[RegFile.scala 97:16:@49783.4]
  assign rport_io_ins_62 = regs_62_io_out; // @[RegFile.scala 97:16:@49784.4]
  assign rport_io_ins_63 = regs_63_io_out; // @[RegFile.scala 97:16:@49785.4]
  assign rport_io_ins_64 = regs_64_io_out; // @[RegFile.scala 97:16:@49786.4]
  assign rport_io_ins_65 = regs_65_io_out; // @[RegFile.scala 97:16:@49787.4]
  assign rport_io_ins_66 = regs_66_io_out; // @[RegFile.scala 97:16:@49788.4]
  assign rport_io_ins_67 = regs_67_io_out; // @[RegFile.scala 97:16:@49789.4]
  assign rport_io_ins_68 = regs_68_io_out; // @[RegFile.scala 97:16:@49790.4]
  assign rport_io_ins_69 = regs_69_io_out; // @[RegFile.scala 97:16:@49791.4]
  assign rport_io_ins_70 = regs_70_io_out; // @[RegFile.scala 97:16:@49792.4]
  assign rport_io_ins_71 = regs_71_io_out; // @[RegFile.scala 97:16:@49793.4]
  assign rport_io_ins_72 = regs_72_io_out; // @[RegFile.scala 97:16:@49794.4]
  assign rport_io_ins_73 = regs_73_io_out; // @[RegFile.scala 97:16:@49795.4]
  assign rport_io_ins_74 = regs_74_io_out; // @[RegFile.scala 97:16:@49796.4]
  assign rport_io_ins_75 = regs_75_io_out; // @[RegFile.scala 97:16:@49797.4]
  assign rport_io_ins_76 = regs_76_io_out; // @[RegFile.scala 97:16:@49798.4]
  assign rport_io_ins_77 = regs_77_io_out; // @[RegFile.scala 97:16:@49799.4]
  assign rport_io_ins_78 = regs_78_io_out; // @[RegFile.scala 97:16:@49800.4]
  assign rport_io_ins_79 = regs_79_io_out; // @[RegFile.scala 97:16:@49801.4]
  assign rport_io_ins_80 = regs_80_io_out; // @[RegFile.scala 97:16:@49802.4]
  assign rport_io_ins_81 = regs_81_io_out; // @[RegFile.scala 97:16:@49803.4]
  assign rport_io_ins_82 = regs_82_io_out; // @[RegFile.scala 97:16:@49804.4]
  assign rport_io_ins_83 = regs_83_io_out; // @[RegFile.scala 97:16:@49805.4]
  assign rport_io_ins_84 = regs_84_io_out; // @[RegFile.scala 97:16:@49806.4]
  assign rport_io_ins_85 = regs_85_io_out; // @[RegFile.scala 97:16:@49807.4]
  assign rport_io_ins_86 = regs_86_io_out; // @[RegFile.scala 97:16:@49808.4]
  assign rport_io_ins_87 = regs_87_io_out; // @[RegFile.scala 97:16:@49809.4]
  assign rport_io_ins_88 = regs_88_io_out; // @[RegFile.scala 97:16:@49810.4]
  assign rport_io_ins_89 = regs_89_io_out; // @[RegFile.scala 97:16:@49811.4]
  assign rport_io_ins_90 = regs_90_io_out; // @[RegFile.scala 97:16:@49812.4]
  assign rport_io_ins_91 = regs_91_io_out; // @[RegFile.scala 97:16:@49813.4]
  assign rport_io_ins_92 = regs_92_io_out; // @[RegFile.scala 97:16:@49814.4]
  assign rport_io_ins_93 = regs_93_io_out; // @[RegFile.scala 97:16:@49815.4]
  assign rport_io_ins_94 = regs_94_io_out; // @[RegFile.scala 97:16:@49816.4]
  assign rport_io_ins_95 = regs_95_io_out; // @[RegFile.scala 97:16:@49817.4]
  assign rport_io_ins_96 = regs_96_io_out; // @[RegFile.scala 97:16:@49818.4]
  assign rport_io_ins_97 = regs_97_io_out; // @[RegFile.scala 97:16:@49819.4]
  assign rport_io_ins_98 = regs_98_io_out; // @[RegFile.scala 97:16:@49820.4]
  assign rport_io_ins_99 = regs_99_io_out; // @[RegFile.scala 97:16:@49821.4]
  assign rport_io_ins_100 = regs_100_io_out; // @[RegFile.scala 97:16:@49822.4]
  assign rport_io_ins_101 = regs_101_io_out; // @[RegFile.scala 97:16:@49823.4]
  assign rport_io_ins_102 = regs_102_io_out; // @[RegFile.scala 97:16:@49824.4]
  assign rport_io_ins_103 = regs_103_io_out; // @[RegFile.scala 97:16:@49825.4]
  assign rport_io_ins_104 = regs_104_io_out; // @[RegFile.scala 97:16:@49826.4]
  assign rport_io_ins_105 = regs_105_io_out; // @[RegFile.scala 97:16:@49827.4]
  assign rport_io_ins_106 = regs_106_io_out; // @[RegFile.scala 97:16:@49828.4]
  assign rport_io_ins_107 = regs_107_io_out; // @[RegFile.scala 97:16:@49829.4]
  assign rport_io_ins_108 = regs_108_io_out; // @[RegFile.scala 97:16:@49830.4]
  assign rport_io_ins_109 = regs_109_io_out; // @[RegFile.scala 97:16:@49831.4]
  assign rport_io_ins_110 = regs_110_io_out; // @[RegFile.scala 97:16:@49832.4]
  assign rport_io_ins_111 = regs_111_io_out; // @[RegFile.scala 97:16:@49833.4]
  assign rport_io_ins_112 = regs_112_io_out; // @[RegFile.scala 97:16:@49834.4]
  assign rport_io_ins_113 = regs_113_io_out; // @[RegFile.scala 97:16:@49835.4]
  assign rport_io_ins_114 = regs_114_io_out; // @[RegFile.scala 97:16:@49836.4]
  assign rport_io_ins_115 = regs_115_io_out; // @[RegFile.scala 97:16:@49837.4]
  assign rport_io_ins_116 = regs_116_io_out; // @[RegFile.scala 97:16:@49838.4]
  assign rport_io_ins_117 = regs_117_io_out; // @[RegFile.scala 97:16:@49839.4]
  assign rport_io_ins_118 = regs_118_io_out; // @[RegFile.scala 97:16:@49840.4]
  assign rport_io_ins_119 = regs_119_io_out; // @[RegFile.scala 97:16:@49841.4]
  assign rport_io_ins_120 = regs_120_io_out; // @[RegFile.scala 97:16:@49842.4]
  assign rport_io_ins_121 = regs_121_io_out; // @[RegFile.scala 97:16:@49843.4]
  assign rport_io_ins_122 = regs_122_io_out; // @[RegFile.scala 97:16:@49844.4]
  assign rport_io_ins_123 = regs_123_io_out; // @[RegFile.scala 97:16:@49845.4]
  assign rport_io_ins_124 = regs_124_io_out; // @[RegFile.scala 97:16:@49846.4]
  assign rport_io_ins_125 = regs_125_io_out; // @[RegFile.scala 97:16:@49847.4]
  assign rport_io_ins_126 = regs_126_io_out; // @[RegFile.scala 97:16:@49848.4]
  assign rport_io_ins_127 = regs_127_io_out; // @[RegFile.scala 97:16:@49849.4]
  assign rport_io_ins_128 = regs_128_io_out; // @[RegFile.scala 97:16:@49850.4]
  assign rport_io_ins_129 = regs_129_io_out; // @[RegFile.scala 97:16:@49851.4]
  assign rport_io_ins_130 = regs_130_io_out; // @[RegFile.scala 97:16:@49852.4]
  assign rport_io_ins_131 = regs_131_io_out; // @[RegFile.scala 97:16:@49853.4]
  assign rport_io_ins_132 = regs_132_io_out; // @[RegFile.scala 97:16:@49854.4]
  assign rport_io_ins_133 = regs_133_io_out; // @[RegFile.scala 97:16:@49855.4]
  assign rport_io_ins_134 = regs_134_io_out; // @[RegFile.scala 97:16:@49856.4]
  assign rport_io_ins_135 = regs_135_io_out; // @[RegFile.scala 97:16:@49857.4]
  assign rport_io_ins_136 = regs_136_io_out; // @[RegFile.scala 97:16:@49858.4]
  assign rport_io_ins_137 = regs_137_io_out; // @[RegFile.scala 97:16:@49859.4]
  assign rport_io_ins_138 = regs_138_io_out; // @[RegFile.scala 97:16:@49860.4]
  assign rport_io_ins_139 = regs_139_io_out; // @[RegFile.scala 97:16:@49861.4]
  assign rport_io_ins_140 = regs_140_io_out; // @[RegFile.scala 97:16:@49862.4]
  assign rport_io_ins_141 = regs_141_io_out; // @[RegFile.scala 97:16:@49863.4]
  assign rport_io_ins_142 = regs_142_io_out; // @[RegFile.scala 97:16:@49864.4]
  assign rport_io_ins_143 = regs_143_io_out; // @[RegFile.scala 97:16:@49865.4]
  assign rport_io_ins_144 = regs_144_io_out; // @[RegFile.scala 97:16:@49866.4]
  assign rport_io_ins_145 = regs_145_io_out; // @[RegFile.scala 97:16:@49867.4]
  assign rport_io_ins_146 = regs_146_io_out; // @[RegFile.scala 97:16:@49868.4]
  assign rport_io_ins_147 = regs_147_io_out; // @[RegFile.scala 97:16:@49869.4]
  assign rport_io_ins_148 = regs_148_io_out; // @[RegFile.scala 97:16:@49870.4]
  assign rport_io_ins_149 = regs_149_io_out; // @[RegFile.scala 97:16:@49871.4]
  assign rport_io_ins_150 = regs_150_io_out; // @[RegFile.scala 97:16:@49872.4]
  assign rport_io_ins_151 = regs_151_io_out; // @[RegFile.scala 97:16:@49873.4]
  assign rport_io_ins_152 = regs_152_io_out; // @[RegFile.scala 97:16:@49874.4]
  assign rport_io_ins_153 = regs_153_io_out; // @[RegFile.scala 97:16:@49875.4]
  assign rport_io_ins_154 = regs_154_io_out; // @[RegFile.scala 97:16:@49876.4]
  assign rport_io_ins_155 = regs_155_io_out; // @[RegFile.scala 97:16:@49877.4]
  assign rport_io_ins_156 = regs_156_io_out; // @[RegFile.scala 97:16:@49878.4]
  assign rport_io_ins_157 = regs_157_io_out; // @[RegFile.scala 97:16:@49879.4]
  assign rport_io_ins_158 = regs_158_io_out; // @[RegFile.scala 97:16:@49880.4]
  assign rport_io_ins_159 = regs_159_io_out; // @[RegFile.scala 97:16:@49881.4]
  assign rport_io_ins_160 = regs_160_io_out; // @[RegFile.scala 97:16:@49882.4]
  assign rport_io_ins_161 = regs_161_io_out; // @[RegFile.scala 97:16:@49883.4]
  assign rport_io_ins_162 = regs_162_io_out; // @[RegFile.scala 97:16:@49884.4]
  assign rport_io_ins_163 = regs_163_io_out; // @[RegFile.scala 97:16:@49885.4]
  assign rport_io_ins_164 = regs_164_io_out; // @[RegFile.scala 97:16:@49886.4]
  assign rport_io_ins_165 = regs_165_io_out; // @[RegFile.scala 97:16:@49887.4]
  assign rport_io_ins_166 = regs_166_io_out; // @[RegFile.scala 97:16:@49888.4]
  assign rport_io_ins_167 = regs_167_io_out; // @[RegFile.scala 97:16:@49889.4]
  assign rport_io_ins_168 = regs_168_io_out; // @[RegFile.scala 97:16:@49890.4]
  assign rport_io_ins_169 = regs_169_io_out; // @[RegFile.scala 97:16:@49891.4]
  assign rport_io_ins_170 = regs_170_io_out; // @[RegFile.scala 97:16:@49892.4]
  assign rport_io_ins_171 = regs_171_io_out; // @[RegFile.scala 97:16:@49893.4]
  assign rport_io_ins_172 = regs_172_io_out; // @[RegFile.scala 97:16:@49894.4]
  assign rport_io_ins_173 = regs_173_io_out; // @[RegFile.scala 97:16:@49895.4]
  assign rport_io_ins_174 = regs_174_io_out; // @[RegFile.scala 97:16:@49896.4]
  assign rport_io_ins_175 = regs_175_io_out; // @[RegFile.scala 97:16:@49897.4]
  assign rport_io_ins_176 = regs_176_io_out; // @[RegFile.scala 97:16:@49898.4]
  assign rport_io_ins_177 = regs_177_io_out; // @[RegFile.scala 97:16:@49899.4]
  assign rport_io_ins_178 = regs_178_io_out; // @[RegFile.scala 97:16:@49900.4]
  assign rport_io_ins_179 = regs_179_io_out; // @[RegFile.scala 97:16:@49901.4]
  assign rport_io_ins_180 = regs_180_io_out; // @[RegFile.scala 97:16:@49902.4]
  assign rport_io_ins_181 = regs_181_io_out; // @[RegFile.scala 97:16:@49903.4]
  assign rport_io_ins_182 = regs_182_io_out; // @[RegFile.scala 97:16:@49904.4]
  assign rport_io_ins_183 = regs_183_io_out; // @[RegFile.scala 97:16:@49905.4]
  assign rport_io_ins_184 = regs_184_io_out; // @[RegFile.scala 97:16:@49906.4]
  assign rport_io_ins_185 = regs_185_io_out; // @[RegFile.scala 97:16:@49907.4]
  assign rport_io_ins_186 = regs_186_io_out; // @[RegFile.scala 97:16:@49908.4]
  assign rport_io_ins_187 = regs_187_io_out; // @[RegFile.scala 97:16:@49909.4]
  assign rport_io_ins_188 = regs_188_io_out; // @[RegFile.scala 97:16:@49910.4]
  assign rport_io_ins_189 = regs_189_io_out; // @[RegFile.scala 97:16:@49911.4]
  assign rport_io_ins_190 = regs_190_io_out; // @[RegFile.scala 97:16:@49912.4]
  assign rport_io_ins_191 = regs_191_io_out; // @[RegFile.scala 97:16:@49913.4]
  assign rport_io_ins_192 = regs_192_io_out; // @[RegFile.scala 97:16:@49914.4]
  assign rport_io_ins_193 = regs_193_io_out; // @[RegFile.scala 97:16:@49915.4]
  assign rport_io_ins_194 = regs_194_io_out; // @[RegFile.scala 97:16:@49916.4]
  assign rport_io_ins_195 = regs_195_io_out; // @[RegFile.scala 97:16:@49917.4]
  assign rport_io_ins_196 = regs_196_io_out; // @[RegFile.scala 97:16:@49918.4]
  assign rport_io_ins_197 = regs_197_io_out; // @[RegFile.scala 97:16:@49919.4]
  assign rport_io_ins_198 = regs_198_io_out; // @[RegFile.scala 97:16:@49920.4]
  assign rport_io_ins_199 = regs_199_io_out; // @[RegFile.scala 97:16:@49921.4]
  assign rport_io_ins_200 = regs_200_io_out; // @[RegFile.scala 97:16:@49922.4]
  assign rport_io_ins_201 = regs_201_io_out; // @[RegFile.scala 97:16:@49923.4]
  assign rport_io_ins_202 = regs_202_io_out; // @[RegFile.scala 97:16:@49924.4]
  assign rport_io_ins_203 = regs_203_io_out; // @[RegFile.scala 97:16:@49925.4]
  assign rport_io_ins_204 = regs_204_io_out; // @[RegFile.scala 97:16:@49926.4]
  assign rport_io_ins_205 = regs_205_io_out; // @[RegFile.scala 97:16:@49927.4]
  assign rport_io_ins_206 = regs_206_io_out; // @[RegFile.scala 97:16:@49928.4]
  assign rport_io_ins_207 = regs_207_io_out; // @[RegFile.scala 97:16:@49929.4]
  assign rport_io_ins_208 = regs_208_io_out; // @[RegFile.scala 97:16:@49930.4]
  assign rport_io_ins_209 = regs_209_io_out; // @[RegFile.scala 97:16:@49931.4]
  assign rport_io_ins_210 = regs_210_io_out; // @[RegFile.scala 97:16:@49932.4]
  assign rport_io_ins_211 = regs_211_io_out; // @[RegFile.scala 97:16:@49933.4]
  assign rport_io_ins_212 = regs_212_io_out; // @[RegFile.scala 97:16:@49934.4]
  assign rport_io_ins_213 = regs_213_io_out; // @[RegFile.scala 97:16:@49935.4]
  assign rport_io_ins_214 = regs_214_io_out; // @[RegFile.scala 97:16:@49936.4]
  assign rport_io_ins_215 = regs_215_io_out; // @[RegFile.scala 97:16:@49937.4]
  assign rport_io_ins_216 = regs_216_io_out; // @[RegFile.scala 97:16:@49938.4]
  assign rport_io_ins_217 = regs_217_io_out; // @[RegFile.scala 97:16:@49939.4]
  assign rport_io_ins_218 = regs_218_io_out; // @[RegFile.scala 97:16:@49940.4]
  assign rport_io_ins_219 = regs_219_io_out; // @[RegFile.scala 97:16:@49941.4]
  assign rport_io_ins_220 = regs_220_io_out; // @[RegFile.scala 97:16:@49942.4]
  assign rport_io_ins_221 = regs_221_io_out; // @[RegFile.scala 97:16:@49943.4]
  assign rport_io_ins_222 = regs_222_io_out; // @[RegFile.scala 97:16:@49944.4]
  assign rport_io_ins_223 = regs_223_io_out; // @[RegFile.scala 97:16:@49945.4]
  assign rport_io_ins_224 = regs_224_io_out; // @[RegFile.scala 97:16:@49946.4]
  assign rport_io_ins_225 = regs_225_io_out; // @[RegFile.scala 97:16:@49947.4]
  assign rport_io_ins_226 = regs_226_io_out; // @[RegFile.scala 97:16:@49948.4]
  assign rport_io_ins_227 = regs_227_io_out; // @[RegFile.scala 97:16:@49949.4]
  assign rport_io_ins_228 = regs_228_io_out; // @[RegFile.scala 97:16:@49950.4]
  assign rport_io_ins_229 = regs_229_io_out; // @[RegFile.scala 97:16:@49951.4]
  assign rport_io_ins_230 = regs_230_io_out; // @[RegFile.scala 97:16:@49952.4]
  assign rport_io_ins_231 = regs_231_io_out; // @[RegFile.scala 97:16:@49953.4]
  assign rport_io_ins_232 = regs_232_io_out; // @[RegFile.scala 97:16:@49954.4]
  assign rport_io_ins_233 = regs_233_io_out; // @[RegFile.scala 97:16:@49955.4]
  assign rport_io_ins_234 = regs_234_io_out; // @[RegFile.scala 97:16:@49956.4]
  assign rport_io_ins_235 = regs_235_io_out; // @[RegFile.scala 97:16:@49957.4]
  assign rport_io_ins_236 = regs_236_io_out; // @[RegFile.scala 97:16:@49958.4]
  assign rport_io_ins_237 = regs_237_io_out; // @[RegFile.scala 97:16:@49959.4]
  assign rport_io_ins_238 = regs_238_io_out; // @[RegFile.scala 97:16:@49960.4]
  assign rport_io_ins_239 = regs_239_io_out; // @[RegFile.scala 97:16:@49961.4]
  assign rport_io_ins_240 = regs_240_io_out; // @[RegFile.scala 97:16:@49962.4]
  assign rport_io_ins_241 = regs_241_io_out; // @[RegFile.scala 97:16:@49963.4]
  assign rport_io_ins_242 = regs_242_io_out; // @[RegFile.scala 97:16:@49964.4]
  assign rport_io_ins_243 = regs_243_io_out; // @[RegFile.scala 97:16:@49965.4]
  assign rport_io_ins_244 = regs_244_io_out; // @[RegFile.scala 97:16:@49966.4]
  assign rport_io_ins_245 = regs_245_io_out; // @[RegFile.scala 97:16:@49967.4]
  assign rport_io_ins_246 = regs_246_io_out; // @[RegFile.scala 97:16:@49968.4]
  assign rport_io_ins_247 = regs_247_io_out; // @[RegFile.scala 97:16:@49969.4]
  assign rport_io_ins_248 = regs_248_io_out; // @[RegFile.scala 97:16:@49970.4]
  assign rport_io_ins_249 = regs_249_io_out; // @[RegFile.scala 97:16:@49971.4]
  assign rport_io_ins_250 = regs_250_io_out; // @[RegFile.scala 97:16:@49972.4]
  assign rport_io_ins_251 = regs_251_io_out; // @[RegFile.scala 97:16:@49973.4]
  assign rport_io_ins_252 = regs_252_io_out; // @[RegFile.scala 97:16:@49974.4]
  assign rport_io_ins_253 = regs_253_io_out; // @[RegFile.scala 97:16:@49975.4]
  assign rport_io_ins_254 = regs_254_io_out; // @[RegFile.scala 97:16:@49976.4]
  assign rport_io_ins_255 = regs_255_io_out; // @[RegFile.scala 97:16:@49977.4]
  assign rport_io_ins_256 = regs_256_io_out; // @[RegFile.scala 97:16:@49978.4]
  assign rport_io_ins_257 = regs_257_io_out; // @[RegFile.scala 97:16:@49979.4]
  assign rport_io_ins_258 = regs_258_io_out; // @[RegFile.scala 97:16:@49980.4]
  assign rport_io_ins_259 = regs_259_io_out; // @[RegFile.scala 97:16:@49981.4]
  assign rport_io_ins_260 = regs_260_io_out; // @[RegFile.scala 97:16:@49982.4]
  assign rport_io_ins_261 = regs_261_io_out; // @[RegFile.scala 97:16:@49983.4]
  assign rport_io_ins_262 = regs_262_io_out; // @[RegFile.scala 97:16:@49984.4]
  assign rport_io_ins_263 = regs_263_io_out; // @[RegFile.scala 97:16:@49985.4]
  assign rport_io_ins_264 = regs_264_io_out; // @[RegFile.scala 97:16:@49986.4]
  assign rport_io_ins_265 = regs_265_io_out; // @[RegFile.scala 97:16:@49987.4]
  assign rport_io_ins_266 = regs_266_io_out; // @[RegFile.scala 97:16:@49988.4]
  assign rport_io_ins_267 = regs_267_io_out; // @[RegFile.scala 97:16:@49989.4]
  assign rport_io_ins_268 = regs_268_io_out; // @[RegFile.scala 97:16:@49990.4]
  assign rport_io_ins_269 = regs_269_io_out; // @[RegFile.scala 97:16:@49991.4]
  assign rport_io_ins_270 = regs_270_io_out; // @[RegFile.scala 97:16:@49992.4]
  assign rport_io_ins_271 = regs_271_io_out; // @[RegFile.scala 97:16:@49993.4]
  assign rport_io_ins_272 = regs_272_io_out; // @[RegFile.scala 97:16:@49994.4]
  assign rport_io_ins_273 = regs_273_io_out; // @[RegFile.scala 97:16:@49995.4]
  assign rport_io_ins_274 = regs_274_io_out; // @[RegFile.scala 97:16:@49996.4]
  assign rport_io_ins_275 = regs_275_io_out; // @[RegFile.scala 97:16:@49997.4]
  assign rport_io_ins_276 = regs_276_io_out; // @[RegFile.scala 97:16:@49998.4]
  assign rport_io_ins_277 = regs_277_io_out; // @[RegFile.scala 97:16:@49999.4]
  assign rport_io_ins_278 = regs_278_io_out; // @[RegFile.scala 97:16:@50000.4]
  assign rport_io_ins_279 = regs_279_io_out; // @[RegFile.scala 97:16:@50001.4]
  assign rport_io_ins_280 = regs_280_io_out; // @[RegFile.scala 97:16:@50002.4]
  assign rport_io_ins_281 = regs_281_io_out; // @[RegFile.scala 97:16:@50003.4]
  assign rport_io_ins_282 = regs_282_io_out; // @[RegFile.scala 97:16:@50004.4]
  assign rport_io_ins_283 = regs_283_io_out; // @[RegFile.scala 97:16:@50005.4]
  assign rport_io_ins_284 = regs_284_io_out; // @[RegFile.scala 97:16:@50006.4]
  assign rport_io_ins_285 = regs_285_io_out; // @[RegFile.scala 97:16:@50007.4]
  assign rport_io_ins_286 = regs_286_io_out; // @[RegFile.scala 97:16:@50008.4]
  assign rport_io_ins_287 = regs_287_io_out; // @[RegFile.scala 97:16:@50009.4]
  assign rport_io_ins_288 = regs_288_io_out; // @[RegFile.scala 97:16:@50010.4]
  assign rport_io_ins_289 = regs_289_io_out; // @[RegFile.scala 97:16:@50011.4]
  assign rport_io_ins_290 = regs_290_io_out; // @[RegFile.scala 97:16:@50012.4]
  assign rport_io_ins_291 = regs_291_io_out; // @[RegFile.scala 97:16:@50013.4]
  assign rport_io_ins_292 = regs_292_io_out; // @[RegFile.scala 97:16:@50014.4]
  assign rport_io_ins_293 = regs_293_io_out; // @[RegFile.scala 97:16:@50015.4]
  assign rport_io_ins_294 = regs_294_io_out; // @[RegFile.scala 97:16:@50016.4]
  assign rport_io_ins_295 = regs_295_io_out; // @[RegFile.scala 97:16:@50017.4]
  assign rport_io_ins_296 = regs_296_io_out; // @[RegFile.scala 97:16:@50018.4]
  assign rport_io_ins_297 = regs_297_io_out; // @[RegFile.scala 97:16:@50019.4]
  assign rport_io_ins_298 = regs_298_io_out; // @[RegFile.scala 97:16:@50020.4]
  assign rport_io_ins_299 = regs_299_io_out; // @[RegFile.scala 97:16:@50021.4]
  assign rport_io_ins_300 = regs_300_io_out; // @[RegFile.scala 97:16:@50022.4]
  assign rport_io_ins_301 = regs_301_io_out; // @[RegFile.scala 97:16:@50023.4]
  assign rport_io_ins_302 = regs_302_io_out; // @[RegFile.scala 97:16:@50024.4]
  assign rport_io_ins_303 = regs_303_io_out; // @[RegFile.scala 97:16:@50025.4]
  assign rport_io_ins_304 = regs_304_io_out; // @[RegFile.scala 97:16:@50026.4]
  assign rport_io_ins_305 = regs_305_io_out; // @[RegFile.scala 97:16:@50027.4]
  assign rport_io_ins_306 = regs_306_io_out; // @[RegFile.scala 97:16:@50028.4]
  assign rport_io_ins_307 = regs_307_io_out; // @[RegFile.scala 97:16:@50029.4]
  assign rport_io_ins_308 = regs_308_io_out; // @[RegFile.scala 97:16:@50030.4]
  assign rport_io_ins_309 = regs_309_io_out; // @[RegFile.scala 97:16:@50031.4]
  assign rport_io_ins_310 = regs_310_io_out; // @[RegFile.scala 97:16:@50032.4]
  assign rport_io_ins_311 = regs_311_io_out; // @[RegFile.scala 97:16:@50033.4]
  assign rport_io_ins_312 = regs_312_io_out; // @[RegFile.scala 97:16:@50034.4]
  assign rport_io_ins_313 = regs_313_io_out; // @[RegFile.scala 97:16:@50035.4]
  assign rport_io_ins_314 = regs_314_io_out; // @[RegFile.scala 97:16:@50036.4]
  assign rport_io_ins_315 = regs_315_io_out; // @[RegFile.scala 97:16:@50037.4]
  assign rport_io_ins_316 = regs_316_io_out; // @[RegFile.scala 97:16:@50038.4]
  assign rport_io_ins_317 = regs_317_io_out; // @[RegFile.scala 97:16:@50039.4]
  assign rport_io_ins_318 = regs_318_io_out; // @[RegFile.scala 97:16:@50040.4]
  assign rport_io_ins_319 = regs_319_io_out; // @[RegFile.scala 97:16:@50041.4]
  assign rport_io_ins_320 = regs_320_io_out; // @[RegFile.scala 97:16:@50042.4]
  assign rport_io_ins_321 = regs_321_io_out; // @[RegFile.scala 97:16:@50043.4]
  assign rport_io_ins_322 = regs_322_io_out; // @[RegFile.scala 97:16:@50044.4]
  assign rport_io_ins_323 = regs_323_io_out; // @[RegFile.scala 97:16:@50045.4]
  assign rport_io_ins_324 = regs_324_io_out; // @[RegFile.scala 97:16:@50046.4]
  assign rport_io_ins_325 = regs_325_io_out; // @[RegFile.scala 97:16:@50047.4]
  assign rport_io_ins_326 = regs_326_io_out; // @[RegFile.scala 97:16:@50048.4]
  assign rport_io_ins_327 = regs_327_io_out; // @[RegFile.scala 97:16:@50049.4]
  assign rport_io_ins_328 = regs_328_io_out; // @[RegFile.scala 97:16:@50050.4]
  assign rport_io_ins_329 = regs_329_io_out; // @[RegFile.scala 97:16:@50051.4]
  assign rport_io_ins_330 = regs_330_io_out; // @[RegFile.scala 97:16:@50052.4]
  assign rport_io_ins_331 = regs_331_io_out; // @[RegFile.scala 97:16:@50053.4]
  assign rport_io_ins_332 = regs_332_io_out; // @[RegFile.scala 97:16:@50054.4]
  assign rport_io_ins_333 = regs_333_io_out; // @[RegFile.scala 97:16:@50055.4]
  assign rport_io_ins_334 = regs_334_io_out; // @[RegFile.scala 97:16:@50056.4]
  assign rport_io_ins_335 = regs_335_io_out; // @[RegFile.scala 97:16:@50057.4]
  assign rport_io_ins_336 = regs_336_io_out; // @[RegFile.scala 97:16:@50058.4]
  assign rport_io_ins_337 = regs_337_io_out; // @[RegFile.scala 97:16:@50059.4]
  assign rport_io_ins_338 = regs_338_io_out; // @[RegFile.scala 97:16:@50060.4]
  assign rport_io_ins_339 = regs_339_io_out; // @[RegFile.scala 97:16:@50061.4]
  assign rport_io_ins_340 = regs_340_io_out; // @[RegFile.scala 97:16:@50062.4]
  assign rport_io_ins_341 = regs_341_io_out; // @[RegFile.scala 97:16:@50063.4]
  assign rport_io_ins_342 = regs_342_io_out; // @[RegFile.scala 97:16:@50064.4]
  assign rport_io_ins_343 = regs_343_io_out; // @[RegFile.scala 97:16:@50065.4]
  assign rport_io_ins_344 = regs_344_io_out; // @[RegFile.scala 97:16:@50066.4]
  assign rport_io_ins_345 = regs_345_io_out; // @[RegFile.scala 97:16:@50067.4]
  assign rport_io_ins_346 = regs_346_io_out; // @[RegFile.scala 97:16:@50068.4]
  assign rport_io_ins_347 = regs_347_io_out; // @[RegFile.scala 97:16:@50069.4]
  assign rport_io_ins_348 = regs_348_io_out; // @[RegFile.scala 97:16:@50070.4]
  assign rport_io_ins_349 = regs_349_io_out; // @[RegFile.scala 97:16:@50071.4]
  assign rport_io_ins_350 = regs_350_io_out; // @[RegFile.scala 97:16:@50072.4]
  assign rport_io_ins_351 = regs_351_io_out; // @[RegFile.scala 97:16:@50073.4]
  assign rport_io_ins_352 = regs_352_io_out; // @[RegFile.scala 97:16:@50074.4]
  assign rport_io_ins_353 = regs_353_io_out; // @[RegFile.scala 97:16:@50075.4]
  assign rport_io_ins_354 = regs_354_io_out; // @[RegFile.scala 97:16:@50076.4]
  assign rport_io_ins_355 = regs_355_io_out; // @[RegFile.scala 97:16:@50077.4]
  assign rport_io_ins_356 = regs_356_io_out; // @[RegFile.scala 97:16:@50078.4]
  assign rport_io_ins_357 = regs_357_io_out; // @[RegFile.scala 97:16:@50079.4]
  assign rport_io_ins_358 = regs_358_io_out; // @[RegFile.scala 97:16:@50080.4]
  assign rport_io_ins_359 = regs_359_io_out; // @[RegFile.scala 97:16:@50081.4]
  assign rport_io_ins_360 = regs_360_io_out; // @[RegFile.scala 97:16:@50082.4]
  assign rport_io_ins_361 = regs_361_io_out; // @[RegFile.scala 97:16:@50083.4]
  assign rport_io_ins_362 = regs_362_io_out; // @[RegFile.scala 97:16:@50084.4]
  assign rport_io_ins_363 = regs_363_io_out; // @[RegFile.scala 97:16:@50085.4]
  assign rport_io_ins_364 = regs_364_io_out; // @[RegFile.scala 97:16:@50086.4]
  assign rport_io_ins_365 = regs_365_io_out; // @[RegFile.scala 97:16:@50087.4]
  assign rport_io_ins_366 = regs_366_io_out; // @[RegFile.scala 97:16:@50088.4]
  assign rport_io_ins_367 = regs_367_io_out; // @[RegFile.scala 97:16:@50089.4]
  assign rport_io_ins_368 = regs_368_io_out; // @[RegFile.scala 97:16:@50090.4]
  assign rport_io_ins_369 = regs_369_io_out; // @[RegFile.scala 97:16:@50091.4]
  assign rport_io_ins_370 = regs_370_io_out; // @[RegFile.scala 97:16:@50092.4]
  assign rport_io_ins_371 = regs_371_io_out; // @[RegFile.scala 97:16:@50093.4]
  assign rport_io_ins_372 = regs_372_io_out; // @[RegFile.scala 97:16:@50094.4]
  assign rport_io_ins_373 = regs_373_io_out; // @[RegFile.scala 97:16:@50095.4]
  assign rport_io_ins_374 = regs_374_io_out; // @[RegFile.scala 97:16:@50096.4]
  assign rport_io_ins_375 = regs_375_io_out; // @[RegFile.scala 97:16:@50097.4]
  assign rport_io_ins_376 = regs_376_io_out; // @[RegFile.scala 97:16:@50098.4]
  assign rport_io_ins_377 = regs_377_io_out; // @[RegFile.scala 97:16:@50099.4]
  assign rport_io_ins_378 = regs_378_io_out; // @[RegFile.scala 97:16:@50100.4]
  assign rport_io_ins_379 = regs_379_io_out; // @[RegFile.scala 97:16:@50101.4]
  assign rport_io_ins_380 = regs_380_io_out; // @[RegFile.scala 97:16:@50102.4]
  assign rport_io_ins_381 = regs_381_io_out; // @[RegFile.scala 97:16:@50103.4]
  assign rport_io_ins_382 = regs_382_io_out; // @[RegFile.scala 97:16:@50104.4]
  assign rport_io_ins_383 = regs_383_io_out; // @[RegFile.scala 97:16:@50105.4]
  assign rport_io_ins_384 = regs_384_io_out; // @[RegFile.scala 97:16:@50106.4]
  assign rport_io_ins_385 = regs_385_io_out; // @[RegFile.scala 97:16:@50107.4]
  assign rport_io_ins_386 = regs_386_io_out; // @[RegFile.scala 97:16:@50108.4]
  assign rport_io_ins_387 = regs_387_io_out; // @[RegFile.scala 97:16:@50109.4]
  assign rport_io_ins_388 = regs_388_io_out; // @[RegFile.scala 97:16:@50110.4]
  assign rport_io_ins_389 = regs_389_io_out; // @[RegFile.scala 97:16:@50111.4]
  assign rport_io_ins_390 = regs_390_io_out; // @[RegFile.scala 97:16:@50112.4]
  assign rport_io_ins_391 = regs_391_io_out; // @[RegFile.scala 97:16:@50113.4]
  assign rport_io_ins_392 = regs_392_io_out; // @[RegFile.scala 97:16:@50114.4]
  assign rport_io_ins_393 = regs_393_io_out; // @[RegFile.scala 97:16:@50115.4]
  assign rport_io_ins_394 = regs_394_io_out; // @[RegFile.scala 97:16:@50116.4]
  assign rport_io_ins_395 = regs_395_io_out; // @[RegFile.scala 97:16:@50117.4]
  assign rport_io_ins_396 = regs_396_io_out; // @[RegFile.scala 97:16:@50118.4]
  assign rport_io_ins_397 = regs_397_io_out; // @[RegFile.scala 97:16:@50119.4]
  assign rport_io_ins_398 = regs_398_io_out; // @[RegFile.scala 97:16:@50120.4]
  assign rport_io_ins_399 = regs_399_io_out; // @[RegFile.scala 97:16:@50121.4]
  assign rport_io_ins_400 = regs_400_io_out; // @[RegFile.scala 97:16:@50122.4]
  assign rport_io_ins_401 = regs_401_io_out; // @[RegFile.scala 97:16:@50123.4]
  assign rport_io_ins_402 = regs_402_io_out; // @[RegFile.scala 97:16:@50124.4]
  assign rport_io_ins_403 = regs_403_io_out; // @[RegFile.scala 97:16:@50125.4]
  assign rport_io_ins_404 = regs_404_io_out; // @[RegFile.scala 97:16:@50126.4]
  assign rport_io_ins_405 = regs_405_io_out; // @[RegFile.scala 97:16:@50127.4]
  assign rport_io_ins_406 = regs_406_io_out; // @[RegFile.scala 97:16:@50128.4]
  assign rport_io_ins_407 = regs_407_io_out; // @[RegFile.scala 97:16:@50129.4]
  assign rport_io_ins_408 = regs_408_io_out; // @[RegFile.scala 97:16:@50130.4]
  assign rport_io_ins_409 = regs_409_io_out; // @[RegFile.scala 97:16:@50131.4]
  assign rport_io_ins_410 = regs_410_io_out; // @[RegFile.scala 97:16:@50132.4]
  assign rport_io_ins_411 = regs_411_io_out; // @[RegFile.scala 97:16:@50133.4]
  assign rport_io_ins_412 = regs_412_io_out; // @[RegFile.scala 97:16:@50134.4]
  assign rport_io_ins_413 = regs_413_io_out; // @[RegFile.scala 97:16:@50135.4]
  assign rport_io_ins_414 = regs_414_io_out; // @[RegFile.scala 97:16:@50136.4]
  assign rport_io_ins_415 = regs_415_io_out; // @[RegFile.scala 97:16:@50137.4]
  assign rport_io_ins_416 = regs_416_io_out; // @[RegFile.scala 97:16:@50138.4]
  assign rport_io_ins_417 = regs_417_io_out; // @[RegFile.scala 97:16:@50139.4]
  assign rport_io_ins_418 = regs_418_io_out; // @[RegFile.scala 97:16:@50140.4]
  assign rport_io_ins_419 = regs_419_io_out; // @[RegFile.scala 97:16:@50141.4]
  assign rport_io_ins_420 = regs_420_io_out; // @[RegFile.scala 97:16:@50142.4]
  assign rport_io_ins_421 = regs_421_io_out; // @[RegFile.scala 97:16:@50143.4]
  assign rport_io_ins_422 = regs_422_io_out; // @[RegFile.scala 97:16:@50144.4]
  assign rport_io_ins_423 = regs_423_io_out; // @[RegFile.scala 97:16:@50145.4]
  assign rport_io_ins_424 = regs_424_io_out; // @[RegFile.scala 97:16:@50146.4]
  assign rport_io_ins_425 = regs_425_io_out; // @[RegFile.scala 97:16:@50147.4]
  assign rport_io_ins_426 = regs_426_io_out; // @[RegFile.scala 97:16:@50148.4]
  assign rport_io_ins_427 = regs_427_io_out; // @[RegFile.scala 97:16:@50149.4]
  assign rport_io_ins_428 = regs_428_io_out; // @[RegFile.scala 97:16:@50150.4]
  assign rport_io_ins_429 = regs_429_io_out; // @[RegFile.scala 97:16:@50151.4]
  assign rport_io_ins_430 = regs_430_io_out; // @[RegFile.scala 97:16:@50152.4]
  assign rport_io_ins_431 = regs_431_io_out; // @[RegFile.scala 97:16:@50153.4]
  assign rport_io_ins_432 = regs_432_io_out; // @[RegFile.scala 97:16:@50154.4]
  assign rport_io_ins_433 = regs_433_io_out; // @[RegFile.scala 97:16:@50155.4]
  assign rport_io_ins_434 = regs_434_io_out; // @[RegFile.scala 97:16:@50156.4]
  assign rport_io_ins_435 = regs_435_io_out; // @[RegFile.scala 97:16:@50157.4]
  assign rport_io_ins_436 = regs_436_io_out; // @[RegFile.scala 97:16:@50158.4]
  assign rport_io_ins_437 = regs_437_io_out; // @[RegFile.scala 97:16:@50159.4]
  assign rport_io_ins_438 = regs_438_io_out; // @[RegFile.scala 97:16:@50160.4]
  assign rport_io_ins_439 = regs_439_io_out; // @[RegFile.scala 97:16:@50161.4]
  assign rport_io_ins_440 = regs_440_io_out; // @[RegFile.scala 97:16:@50162.4]
  assign rport_io_ins_441 = regs_441_io_out; // @[RegFile.scala 97:16:@50163.4]
  assign rport_io_ins_442 = regs_442_io_out; // @[RegFile.scala 97:16:@50164.4]
  assign rport_io_ins_443 = regs_443_io_out; // @[RegFile.scala 97:16:@50165.4]
  assign rport_io_ins_444 = regs_444_io_out; // @[RegFile.scala 97:16:@50166.4]
  assign rport_io_ins_445 = regs_445_io_out; // @[RegFile.scala 97:16:@50167.4]
  assign rport_io_ins_446 = regs_446_io_out; // @[RegFile.scala 97:16:@50168.4]
  assign rport_io_ins_447 = regs_447_io_out; // @[RegFile.scala 97:16:@50169.4]
  assign rport_io_ins_448 = regs_448_io_out; // @[RegFile.scala 97:16:@50170.4]
  assign rport_io_ins_449 = regs_449_io_out; // @[RegFile.scala 97:16:@50171.4]
  assign rport_io_ins_450 = regs_450_io_out; // @[RegFile.scala 97:16:@50172.4]
  assign rport_io_ins_451 = regs_451_io_out; // @[RegFile.scala 97:16:@50173.4]
  assign rport_io_ins_452 = regs_452_io_out; // @[RegFile.scala 97:16:@50174.4]
  assign rport_io_ins_453 = regs_453_io_out; // @[RegFile.scala 97:16:@50175.4]
  assign rport_io_ins_454 = regs_454_io_out; // @[RegFile.scala 97:16:@50176.4]
  assign rport_io_ins_455 = regs_455_io_out; // @[RegFile.scala 97:16:@50177.4]
  assign rport_io_ins_456 = regs_456_io_out; // @[RegFile.scala 97:16:@50178.4]
  assign rport_io_ins_457 = regs_457_io_out; // @[RegFile.scala 97:16:@50179.4]
  assign rport_io_ins_458 = regs_458_io_out; // @[RegFile.scala 97:16:@50180.4]
  assign rport_io_ins_459 = regs_459_io_out; // @[RegFile.scala 97:16:@50181.4]
  assign rport_io_ins_460 = regs_460_io_out; // @[RegFile.scala 97:16:@50182.4]
  assign rport_io_ins_461 = regs_461_io_out; // @[RegFile.scala 97:16:@50183.4]
  assign rport_io_ins_462 = regs_462_io_out; // @[RegFile.scala 97:16:@50184.4]
  assign rport_io_ins_463 = regs_463_io_out; // @[RegFile.scala 97:16:@50185.4]
  assign rport_io_ins_464 = regs_464_io_out; // @[RegFile.scala 97:16:@50186.4]
  assign rport_io_ins_465 = regs_465_io_out; // @[RegFile.scala 97:16:@50187.4]
  assign rport_io_ins_466 = regs_466_io_out; // @[RegFile.scala 97:16:@50188.4]
  assign rport_io_ins_467 = regs_467_io_out; // @[RegFile.scala 97:16:@50189.4]
  assign rport_io_ins_468 = regs_468_io_out; // @[RegFile.scala 97:16:@50190.4]
  assign rport_io_ins_469 = regs_469_io_out; // @[RegFile.scala 97:16:@50191.4]
  assign rport_io_ins_470 = regs_470_io_out; // @[RegFile.scala 97:16:@50192.4]
  assign rport_io_ins_471 = regs_471_io_out; // @[RegFile.scala 97:16:@50193.4]
  assign rport_io_ins_472 = regs_472_io_out; // @[RegFile.scala 97:16:@50194.4]
  assign rport_io_ins_473 = regs_473_io_out; // @[RegFile.scala 97:16:@50195.4]
  assign rport_io_ins_474 = regs_474_io_out; // @[RegFile.scala 97:16:@50196.4]
  assign rport_io_ins_475 = regs_475_io_out; // @[RegFile.scala 97:16:@50197.4]
  assign rport_io_ins_476 = regs_476_io_out; // @[RegFile.scala 97:16:@50198.4]
  assign rport_io_ins_477 = regs_477_io_out; // @[RegFile.scala 97:16:@50199.4]
  assign rport_io_ins_478 = regs_478_io_out; // @[RegFile.scala 97:16:@50200.4]
  assign rport_io_ins_479 = regs_479_io_out; // @[RegFile.scala 97:16:@50201.4]
  assign rport_io_ins_480 = regs_480_io_out; // @[RegFile.scala 97:16:@50202.4]
  assign rport_io_ins_481 = regs_481_io_out; // @[RegFile.scala 97:16:@50203.4]
  assign rport_io_ins_482 = regs_482_io_out; // @[RegFile.scala 97:16:@50204.4]
  assign rport_io_ins_483 = regs_483_io_out; // @[RegFile.scala 97:16:@50205.4]
  assign rport_io_ins_484 = regs_484_io_out; // @[RegFile.scala 97:16:@50206.4]
  assign rport_io_ins_485 = regs_485_io_out; // @[RegFile.scala 97:16:@50207.4]
  assign rport_io_ins_486 = regs_486_io_out; // @[RegFile.scala 97:16:@50208.4]
  assign rport_io_ins_487 = regs_487_io_out; // @[RegFile.scala 97:16:@50209.4]
  assign rport_io_ins_488 = regs_488_io_out; // @[RegFile.scala 97:16:@50210.4]
  assign rport_io_ins_489 = regs_489_io_out; // @[RegFile.scala 97:16:@50211.4]
  assign rport_io_ins_490 = regs_490_io_out; // @[RegFile.scala 97:16:@50212.4]
  assign rport_io_ins_491 = regs_491_io_out; // @[RegFile.scala 97:16:@50213.4]
  assign rport_io_ins_492 = regs_492_io_out; // @[RegFile.scala 97:16:@50214.4]
  assign rport_io_ins_493 = regs_493_io_out; // @[RegFile.scala 97:16:@50215.4]
  assign rport_io_ins_494 = regs_494_io_out; // @[RegFile.scala 97:16:@50216.4]
  assign rport_io_ins_495 = regs_495_io_out; // @[RegFile.scala 97:16:@50217.4]
  assign rport_io_ins_496 = regs_496_io_out; // @[RegFile.scala 97:16:@50218.4]
  assign rport_io_ins_497 = regs_497_io_out; // @[RegFile.scala 97:16:@50219.4]
  assign rport_io_ins_498 = regs_498_io_out; // @[RegFile.scala 97:16:@50220.4]
  assign rport_io_ins_499 = regs_499_io_out; // @[RegFile.scala 97:16:@50221.4]
  assign rport_io_ins_500 = regs_500_io_out; // @[RegFile.scala 97:16:@50222.4]
  assign rport_io_ins_501 = regs_501_io_out; // @[RegFile.scala 97:16:@50223.4]
  assign rport_io_ins_502 = regs_502_io_out; // @[RegFile.scala 97:16:@50224.4]
  assign rport_io_ins_503 = regs_503_io_out; // @[RegFile.scala 97:16:@50225.4]
  assign rport_io_ins_504 = regs_504_io_out; // @[RegFile.scala 97:16:@50226.4]
  assign rport_io_ins_505 = regs_505_io_out; // @[RegFile.scala 97:16:@50227.4]
  assign rport_io_ins_506 = regs_506_io_out; // @[RegFile.scala 97:16:@50228.4]
  assign rport_io_ins_507 = regs_507_io_out; // @[RegFile.scala 97:16:@50229.4]
  assign rport_io_ins_508 = regs_508_io_out; // @[RegFile.scala 97:16:@50230.4]
  assign rport_io_ins_509 = regs_509_io_out; // @[RegFile.scala 97:16:@50231.4]
  assign rport_io_ins_510 = regs_510_io_out; // @[RegFile.scala 97:16:@50232.4]
  assign rport_io_ins_511 = regs_511_io_out; // @[RegFile.scala 97:16:@50233.4]
  assign rport_io_ins_512 = regs_512_io_out; // @[RegFile.scala 97:16:@50234.4]
  assign rport_io_ins_513 = regs_513_io_out; // @[RegFile.scala 97:16:@50235.4]
  assign rport_io_ins_514 = regs_514_io_out; // @[RegFile.scala 97:16:@50236.4]
  assign rport_io_ins_515 = regs_515_io_out; // @[RegFile.scala 97:16:@50237.4]
  assign rport_io_ins_516 = regs_516_io_out; // @[RegFile.scala 97:16:@50238.4]
  assign rport_io_ins_517 = regs_517_io_out; // @[RegFile.scala 97:16:@50239.4]
  assign rport_io_ins_518 = regs_518_io_out; // @[RegFile.scala 97:16:@50240.4]
  assign rport_io_ins_519 = regs_519_io_out; // @[RegFile.scala 97:16:@50241.4]
  assign rport_io_ins_520 = regs_520_io_out; // @[RegFile.scala 97:16:@50242.4]
  assign rport_io_ins_521 = regs_521_io_out; // @[RegFile.scala 97:16:@50243.4]
  assign rport_io_sel = io_raddr[9:0]; // @[RegFile.scala 106:18:@50244.4]
endmodule
module RetimeWrapper_590( // @[:@50266.2]
  input         clock, // @[:@50267.4]
  input         reset, // @[:@50268.4]
  input  [39:0] io_in, // @[:@50269.4]
  output [39:0] io_out // @[:@50269.4]
);
  wire [39:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@50271.4]
  wire [39:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@50271.4]
  wire [39:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@50271.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@50271.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@50271.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@50271.4]
  RetimeShiftRegister #(.WIDTH(40), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@50271.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@50284.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@50283.4]
  assign sr_init = 40'h0; // @[RetimeShiftRegister.scala 19:16:@50282.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@50281.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@50280.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@50278.4]
endmodule
module FringeFF_522( // @[:@50286.2]
  input         clock, // @[:@50287.4]
  input         reset, // @[:@50288.4]
  input  [39:0] io_in, // @[:@50289.4]
  output [39:0] io_out, // @[:@50289.4]
  input         io_enable // @[:@50289.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@50292.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@50292.4]
  wire [39:0] RetimeWrapper_io_in; // @[package.scala 93:22:@50292.4]
  wire [39:0] RetimeWrapper_io_out; // @[package.scala 93:22:@50292.4]
  wire [39:0] _T_18; // @[package.scala 96:25:@50297.4 package.scala 96:25:@50298.4]
  RetimeWrapper_590 RetimeWrapper ( // @[package.scala 93:22:@50292.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@50297.4 package.scala 96:25:@50298.4]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@50309.4]
  assign RetimeWrapper_clock = clock; // @[:@50293.4]
  assign RetimeWrapper_reset = reset; // @[:@50294.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _T_18; // @[package.scala 94:16:@50295.4]
endmodule
module FringeCounter( // @[:@50311.2]
  input   clock, // @[:@50312.4]
  input   reset, // @[:@50313.4]
  input   io_enable, // @[:@50314.4]
  output  io_done // @[:@50314.4]
);
  wire  reg$_clock; // @[FringeCounter.scala 24:19:@50316.4]
  wire  reg$_reset; // @[FringeCounter.scala 24:19:@50316.4]
  wire [39:0] reg$_io_in; // @[FringeCounter.scala 24:19:@50316.4]
  wire [39:0] reg$_io_out; // @[FringeCounter.scala 24:19:@50316.4]
  wire  reg$_io_enable; // @[FringeCounter.scala 24:19:@50316.4]
  wire [40:0] count; // @[Cat.scala 30:58:@50323.4]
  wire [41:0] _T_25; // @[FringeCounter.scala 31:22:@50324.4]
  wire [40:0] newval; // @[FringeCounter.scala 31:22:@50325.4]
  wire  isMax; // @[FringeCounter.scala 32:22:@50326.4]
  wire [40:0] next; // @[FringeCounter.scala 33:17:@50328.4]
  FringeFF_522 reg$ ( // @[FringeCounter.scala 24:19:@50316.4]
    .clock(reg$_clock),
    .reset(reg$_reset),
    .io_in(reg$_io_in),
    .io_out(reg$_io_out),
    .io_enable(reg$_io_enable)
  );
  assign count = {1'h0,reg$_io_out}; // @[Cat.scala 30:58:@50323.4]
  assign _T_25 = count + 41'h1; // @[FringeCounter.scala 31:22:@50324.4]
  assign newval = count + 41'h1; // @[FringeCounter.scala 31:22:@50325.4]
  assign isMax = newval >= 41'h2cb417800; // @[FringeCounter.scala 32:22:@50326.4]
  assign next = isMax ? count : newval; // @[FringeCounter.scala 33:17:@50328.4]
  assign io_done = io_enable & isMax; // @[FringeCounter.scala 43:11:@50339.4]
  assign reg$_clock = clock; // @[:@50317.4]
  assign reg$_reset = reset; // @[:@50318.4]
  assign reg$_io_in = next[39:0]; // @[FringeCounter.scala 35:15:@50330.6 FringeCounter.scala 37:15:@50333.6]
  assign reg$_io_enable = io_enable; // @[FringeCounter.scala 27:17:@50321.4]
endmodule
module FringeFF_523( // @[:@50373.2]
  input   clock, // @[:@50374.4]
  input   reset, // @[:@50375.4]
  input   io_in, // @[:@50376.4]
  input   io_reset, // @[:@50376.4]
  output  io_out, // @[:@50376.4]
  input   io_enable // @[:@50376.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@50379.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@50379.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@50379.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@50379.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@50379.4]
  wire  _T_18; // @[package.scala 96:25:@50384.4 package.scala 96:25:@50385.4]
  wire  _GEN_0; // @[FringeFF.scala 21:27:@50390.6]
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@50379.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@50384.4 package.scala 96:25:@50385.4]
  assign _GEN_0 = io_reset ? 1'h0 : _T_18; // @[FringeFF.scala 21:27:@50390.6]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@50396.4]
  assign RetimeWrapper_clock = clock; // @[:@50380.4]
  assign RetimeWrapper_reset = reset; // @[:@50381.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@50383.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _GEN_0; // @[package.scala 94:16:@50382.4]
endmodule
module Depulser( // @[:@50398.2]
  input   clock, // @[:@50399.4]
  input   reset, // @[:@50400.4]
  input   io_in, // @[:@50401.4]
  input   io_rst, // @[:@50401.4]
  output  io_out // @[:@50401.4]
);
  wire  r_clock; // @[Depulser.scala 14:17:@50403.4]
  wire  r_reset; // @[Depulser.scala 14:17:@50403.4]
  wire  r_io_in; // @[Depulser.scala 14:17:@50403.4]
  wire  r_io_reset; // @[Depulser.scala 14:17:@50403.4]
  wire  r_io_out; // @[Depulser.scala 14:17:@50403.4]
  wire  r_io_enable; // @[Depulser.scala 14:17:@50403.4]
  FringeFF_523 r ( // @[Depulser.scala 14:17:@50403.4]
    .clock(r_clock),
    .reset(r_reset),
    .io_in(r_io_in),
    .io_reset(r_io_reset),
    .io_out(r_io_out),
    .io_enable(r_io_enable)
  );
  assign io_out = r_io_out; // @[Depulser.scala 19:10:@50412.4]
  assign r_clock = clock; // @[:@50404.4]
  assign r_reset = reset; // @[:@50405.4]
  assign r_io_in = io_rst ? 1'h0 : io_in; // @[Depulser.scala 15:11:@50407.4]
  assign r_io_reset = io_rst; // @[Depulser.scala 18:14:@50411.4]
  assign r_io_enable = io_in | io_rst; // @[Depulser.scala 17:15:@50410.4]
endmodule
module Fringe( // @[:@50414.2]
  input         clock, // @[:@50415.4]
  input         reset, // @[:@50416.4]
  input  [31:0] io_raddr, // @[:@50417.4]
  input         io_wen, // @[:@50417.4]
  input  [31:0] io_waddr, // @[:@50417.4]
  input  [63:0] io_wdata, // @[:@50417.4]
  output [63:0] io_rdata, // @[:@50417.4]
  output        io_enable, // @[:@50417.4]
  input         io_done, // @[:@50417.4]
  output        io_reset, // @[:@50417.4]
  output [63:0] io_argIns_0, // @[:@50417.4]
  input         io_argOuts_0_valid, // @[:@50417.4]
  input  [63:0] io_argOuts_0_bits, // @[:@50417.4]
  input         io_argOuts_1_valid, // @[:@50417.4]
  input  [63:0] io_argOuts_1_bits, // @[:@50417.4]
  input         io_argOuts_2_valid, // @[:@50417.4]
  input  [63:0] io_argOuts_2_bits, // @[:@50417.4]
  input         io_argOuts_3_valid, // @[:@50417.4]
  input  [63:0] io_argOuts_3_bits, // @[:@50417.4]
  input         io_argOuts_4_valid, // @[:@50417.4]
  input  [63:0] io_argOuts_4_bits, // @[:@50417.4]
  input         io_argOuts_5_valid, // @[:@50417.4]
  input  [63:0] io_argOuts_5_bits, // @[:@50417.4]
  input         io_argOuts_6_valid, // @[:@50417.4]
  input  [63:0] io_argOuts_6_bits, // @[:@50417.4]
  input         io_argOuts_7_valid, // @[:@50417.4]
  input  [63:0] io_argOuts_7_bits, // @[:@50417.4]
  input         io_argOuts_8_valid, // @[:@50417.4]
  input  [63:0] io_argOuts_8_bits, // @[:@50417.4]
  input         io_argOuts_9_valid, // @[:@50417.4]
  input  [63:0] io_argOuts_9_bits, // @[:@50417.4]
  input         io_argOuts_10_valid, // @[:@50417.4]
  input  [63:0] io_argOuts_10_bits, // @[:@50417.4]
  input         io_argOuts_11_valid, // @[:@50417.4]
  input  [63:0] io_argOuts_11_bits, // @[:@50417.4]
  input         io_argOuts_12_valid, // @[:@50417.4]
  input  [63:0] io_argOuts_12_bits, // @[:@50417.4]
  input         io_argOuts_13_valid, // @[:@50417.4]
  input  [63:0] io_argOuts_13_bits, // @[:@50417.4]
  input         io_argOuts_14_valid, // @[:@50417.4]
  input  [63:0] io_argOuts_14_bits, // @[:@50417.4]
  input         io_argOuts_15_valid, // @[:@50417.4]
  input  [63:0] io_argOuts_15_bits, // @[:@50417.4]
  input         io_argOuts_16_valid, // @[:@50417.4]
  input  [63:0] io_argOuts_16_bits, // @[:@50417.4]
  input         io_argOuts_17_valid, // @[:@50417.4]
  input  [63:0] io_argOuts_17_bits, // @[:@50417.4]
  input         io_argOuts_18_valid, // @[:@50417.4]
  input  [63:0] io_argOuts_18_bits, // @[:@50417.4]
  input         io_argOuts_19_valid, // @[:@50417.4]
  input  [63:0] io_argOuts_19_bits, // @[:@50417.4]
  input         io_heap_0_req_valid, // @[:@50417.4]
  input         io_heap_0_req_bits_allocDealloc, // @[:@50417.4]
  input  [63:0] io_heap_0_req_bits_sizeAddr, // @[:@50417.4]
  output        io_heap_0_resp_valid, // @[:@50417.4]
  output        io_heap_0_resp_bits_allocDealloc, // @[:@50417.4]
  output [63:0] io_heap_0_resp_bits_sizeAddr // @[:@50417.4]
);
  wire  heap_io_accel_0_req_valid; // @[Fringe.scala 107:20:@51522.4]
  wire  heap_io_accel_0_req_bits_allocDealloc; // @[Fringe.scala 107:20:@51522.4]
  wire [63:0] heap_io_accel_0_req_bits_sizeAddr; // @[Fringe.scala 107:20:@51522.4]
  wire  heap_io_accel_0_resp_valid; // @[Fringe.scala 107:20:@51522.4]
  wire  heap_io_accel_0_resp_bits_allocDealloc; // @[Fringe.scala 107:20:@51522.4]
  wire [63:0] heap_io_accel_0_resp_bits_sizeAddr; // @[Fringe.scala 107:20:@51522.4]
  wire  heap_io_host_0_req_valid; // @[Fringe.scala 107:20:@51522.4]
  wire  heap_io_host_0_req_bits_allocDealloc; // @[Fringe.scala 107:20:@51522.4]
  wire [63:0] heap_io_host_0_req_bits_sizeAddr; // @[Fringe.scala 107:20:@51522.4]
  wire  heap_io_host_0_resp_valid; // @[Fringe.scala 107:20:@51522.4]
  wire  heap_io_host_0_resp_bits_allocDealloc; // @[Fringe.scala 107:20:@51522.4]
  wire [63:0] heap_io_host_0_resp_bits_sizeAddr; // @[Fringe.scala 107:20:@51522.4]
  wire  regs_clock; // @[Fringe.scala 116:20:@51531.4]
  wire  regs_reset; // @[Fringe.scala 116:20:@51531.4]
  wire [31:0] regs_io_raddr; // @[Fringe.scala 116:20:@51531.4]
  wire  regs_io_wen; // @[Fringe.scala 116:20:@51531.4]
  wire [31:0] regs_io_waddr; // @[Fringe.scala 116:20:@51531.4]
  wire [63:0] regs_io_wdata; // @[Fringe.scala 116:20:@51531.4]
  wire [63:0] regs_io_rdata; // @[Fringe.scala 116:20:@51531.4]
  wire  regs_io_reset; // @[Fringe.scala 116:20:@51531.4]
  wire [63:0] regs_io_argIns_0; // @[Fringe.scala 116:20:@51531.4]
  wire [63:0] regs_io_argIns_1; // @[Fringe.scala 116:20:@51531.4]
  wire [63:0] regs_io_argIns_2; // @[Fringe.scala 116:20:@51531.4]
  wire  regs_io_argOuts_0_valid; // @[Fringe.scala 116:20:@51531.4]
  wire [63:0] regs_io_argOuts_0_bits; // @[Fringe.scala 116:20:@51531.4]
  wire  regs_io_argOuts_1_valid; // @[Fringe.scala 116:20:@51531.4]
  wire [63:0] regs_io_argOuts_1_bits; // @[Fringe.scala 116:20:@51531.4]
  wire  regs_io_argOuts_2_valid; // @[Fringe.scala 116:20:@51531.4]
  wire [63:0] regs_io_argOuts_2_bits; // @[Fringe.scala 116:20:@51531.4]
  wire  regs_io_argOuts_3_valid; // @[Fringe.scala 116:20:@51531.4]
  wire [63:0] regs_io_argOuts_3_bits; // @[Fringe.scala 116:20:@51531.4]
  wire  regs_io_argOuts_4_valid; // @[Fringe.scala 116:20:@51531.4]
  wire [63:0] regs_io_argOuts_4_bits; // @[Fringe.scala 116:20:@51531.4]
  wire  regs_io_argOuts_5_valid; // @[Fringe.scala 116:20:@51531.4]
  wire [63:0] regs_io_argOuts_5_bits; // @[Fringe.scala 116:20:@51531.4]
  wire  regs_io_argOuts_6_valid; // @[Fringe.scala 116:20:@51531.4]
  wire [63:0] regs_io_argOuts_6_bits; // @[Fringe.scala 116:20:@51531.4]
  wire  regs_io_argOuts_7_valid; // @[Fringe.scala 116:20:@51531.4]
  wire [63:0] regs_io_argOuts_7_bits; // @[Fringe.scala 116:20:@51531.4]
  wire  regs_io_argOuts_8_valid; // @[Fringe.scala 116:20:@51531.4]
  wire [63:0] regs_io_argOuts_8_bits; // @[Fringe.scala 116:20:@51531.4]
  wire  regs_io_argOuts_9_valid; // @[Fringe.scala 116:20:@51531.4]
  wire [63:0] regs_io_argOuts_9_bits; // @[Fringe.scala 116:20:@51531.4]
  wire  regs_io_argOuts_10_valid; // @[Fringe.scala 116:20:@51531.4]
  wire [63:0] regs_io_argOuts_10_bits; // @[Fringe.scala 116:20:@51531.4]
  wire  regs_io_argOuts_11_valid; // @[Fringe.scala 116:20:@51531.4]
  wire [63:0] regs_io_argOuts_11_bits; // @[Fringe.scala 116:20:@51531.4]
  wire  regs_io_argOuts_12_valid; // @[Fringe.scala 116:20:@51531.4]
  wire [63:0] regs_io_argOuts_12_bits; // @[Fringe.scala 116:20:@51531.4]
  wire  regs_io_argOuts_13_valid; // @[Fringe.scala 116:20:@51531.4]
  wire [63:0] regs_io_argOuts_13_bits; // @[Fringe.scala 116:20:@51531.4]
  wire  regs_io_argOuts_14_valid; // @[Fringe.scala 116:20:@51531.4]
  wire [63:0] regs_io_argOuts_14_bits; // @[Fringe.scala 116:20:@51531.4]
  wire  regs_io_argOuts_15_valid; // @[Fringe.scala 116:20:@51531.4]
  wire [63:0] regs_io_argOuts_15_bits; // @[Fringe.scala 116:20:@51531.4]
  wire  regs_io_argOuts_16_valid; // @[Fringe.scala 116:20:@51531.4]
  wire [63:0] regs_io_argOuts_16_bits; // @[Fringe.scala 116:20:@51531.4]
  wire  regs_io_argOuts_17_valid; // @[Fringe.scala 116:20:@51531.4]
  wire [63:0] regs_io_argOuts_17_bits; // @[Fringe.scala 116:20:@51531.4]
  wire  regs_io_argOuts_18_valid; // @[Fringe.scala 116:20:@51531.4]
  wire [63:0] regs_io_argOuts_18_bits; // @[Fringe.scala 116:20:@51531.4]
  wire  regs_io_argOuts_19_valid; // @[Fringe.scala 116:20:@51531.4]
  wire [63:0] regs_io_argOuts_19_bits; // @[Fringe.scala 116:20:@51531.4]
  wire  regs_io_argOuts_20_valid; // @[Fringe.scala 116:20:@51531.4]
  wire [63:0] regs_io_argOuts_20_bits; // @[Fringe.scala 116:20:@51531.4]
  wire  timeoutCtr_clock; // @[Fringe.scala 143:26:@53656.4]
  wire  timeoutCtr_reset; // @[Fringe.scala 143:26:@53656.4]
  wire  timeoutCtr_io_enable; // @[Fringe.scala 143:26:@53656.4]
  wire  timeoutCtr_io_done; // @[Fringe.scala 143:26:@53656.4]
  wire  depulser_clock; // @[Fringe.scala 153:24:@53674.4]
  wire  depulser_reset; // @[Fringe.scala 153:24:@53674.4]
  wire  depulser_io_in; // @[Fringe.scala 153:24:@53674.4]
  wire  depulser_io_rst; // @[Fringe.scala 153:24:@53674.4]
  wire  depulser_io_out; // @[Fringe.scala 153:24:@53674.4]
  wire [63:0] _T_940; // @[:@53633.4 :@53634.4]
  wire  curStatus_done; // @[Fringe.scala 133:45:@53635.4]
  wire  curStatus_timeout; // @[Fringe.scala 133:45:@53637.4]
  wire [2:0] curStatus_allocDealloc; // @[Fringe.scala 133:45:@53639.4]
  wire [58:0] curStatus_sizeAddr; // @[Fringe.scala 133:45:@53641.4]
  wire  _T_945; // @[Fringe.scala 134:28:@53643.4]
  wire  _T_949; // @[Fringe.scala 134:42:@53645.4]
  wire  _T_950; // @[Fringe.scala 135:27:@53647.4]
  wire [63:0] _T_960; // @[Fringe.scala 156:22:@53682.4]
  reg  _T_967; // @[package.scala 152:20:@53685.4]
  reg [31:0] _RAND_0;
  wire  _T_968; // @[package.scala 153:13:@53687.4]
  wire  _T_969; // @[package.scala 153:8:@53688.4]
  wire  _T_972; // @[Fringe.scala 160:55:@53692.4]
  wire  status_bits_done; // @[Fringe.scala 160:26:@53693.4]
  wire  _T_975; // @[Fringe.scala 161:58:@53696.4]
  wire  status_bits_timeout; // @[Fringe.scala 161:29:@53697.4]
  wire [1:0] _T_979; // @[Fringe.scala 162:57:@53699.4]
  wire [1:0] _T_981; // @[Fringe.scala 162:34:@53700.4]
  wire [63:0] _T_983; // @[Fringe.scala 163:30:@53702.4]
  wire [1:0] _T_984; // @[Fringe.scala 171:37:@53705.4]
  wire [58:0] status_bits_sizeAddr; // @[Fringe.scala 158:20:@53684.4 Fringe.scala 163:24:@53703.4]
  wire [2:0] status_bits_allocDealloc; // @[Fringe.scala 158:20:@53684.4 Fringe.scala 162:28:@53701.4]
  wire [61:0] _T_985; // @[Fringe.scala 171:37:@53706.4]
  wire  alloc; // @[Fringe.scala 202:38:@55048.4]
  wire  dealloc; // @[Fringe.scala 203:40:@55049.4]
  wire  _T_1489; // @[Fringe.scala 204:37:@55050.4]
  reg  _T_1492; // @[package.scala 152:20:@55051.4]
  reg [31:0] _RAND_1;
  wire  _T_1493; // @[package.scala 153:13:@55053.4]
  DRAMHeap heap ( // @[Fringe.scala 107:20:@51522.4]
    .io_accel_0_req_valid(heap_io_accel_0_req_valid),
    .io_accel_0_req_bits_allocDealloc(heap_io_accel_0_req_bits_allocDealloc),
    .io_accel_0_req_bits_sizeAddr(heap_io_accel_0_req_bits_sizeAddr),
    .io_accel_0_resp_valid(heap_io_accel_0_resp_valid),
    .io_accel_0_resp_bits_allocDealloc(heap_io_accel_0_resp_bits_allocDealloc),
    .io_accel_0_resp_bits_sizeAddr(heap_io_accel_0_resp_bits_sizeAddr),
    .io_host_0_req_valid(heap_io_host_0_req_valid),
    .io_host_0_req_bits_allocDealloc(heap_io_host_0_req_bits_allocDealloc),
    .io_host_0_req_bits_sizeAddr(heap_io_host_0_req_bits_sizeAddr),
    .io_host_0_resp_valid(heap_io_host_0_resp_valid),
    .io_host_0_resp_bits_allocDealloc(heap_io_host_0_resp_bits_allocDealloc),
    .io_host_0_resp_bits_sizeAddr(heap_io_host_0_resp_bits_sizeAddr)
  );
  RegFile regs ( // @[Fringe.scala 116:20:@51531.4]
    .clock(regs_clock),
    .reset(regs_reset),
    .io_raddr(regs_io_raddr),
    .io_wen(regs_io_wen),
    .io_waddr(regs_io_waddr),
    .io_wdata(regs_io_wdata),
    .io_rdata(regs_io_rdata),
    .io_reset(regs_io_reset),
    .io_argIns_0(regs_io_argIns_0),
    .io_argIns_1(regs_io_argIns_1),
    .io_argIns_2(regs_io_argIns_2),
    .io_argOuts_0_valid(regs_io_argOuts_0_valid),
    .io_argOuts_0_bits(regs_io_argOuts_0_bits),
    .io_argOuts_1_valid(regs_io_argOuts_1_valid),
    .io_argOuts_1_bits(regs_io_argOuts_1_bits),
    .io_argOuts_2_valid(regs_io_argOuts_2_valid),
    .io_argOuts_2_bits(regs_io_argOuts_2_bits),
    .io_argOuts_3_valid(regs_io_argOuts_3_valid),
    .io_argOuts_3_bits(regs_io_argOuts_3_bits),
    .io_argOuts_4_valid(regs_io_argOuts_4_valid),
    .io_argOuts_4_bits(regs_io_argOuts_4_bits),
    .io_argOuts_5_valid(regs_io_argOuts_5_valid),
    .io_argOuts_5_bits(regs_io_argOuts_5_bits),
    .io_argOuts_6_valid(regs_io_argOuts_6_valid),
    .io_argOuts_6_bits(regs_io_argOuts_6_bits),
    .io_argOuts_7_valid(regs_io_argOuts_7_valid),
    .io_argOuts_7_bits(regs_io_argOuts_7_bits),
    .io_argOuts_8_valid(regs_io_argOuts_8_valid),
    .io_argOuts_8_bits(regs_io_argOuts_8_bits),
    .io_argOuts_9_valid(regs_io_argOuts_9_valid),
    .io_argOuts_9_bits(regs_io_argOuts_9_bits),
    .io_argOuts_10_valid(regs_io_argOuts_10_valid),
    .io_argOuts_10_bits(regs_io_argOuts_10_bits),
    .io_argOuts_11_valid(regs_io_argOuts_11_valid),
    .io_argOuts_11_bits(regs_io_argOuts_11_bits),
    .io_argOuts_12_valid(regs_io_argOuts_12_valid),
    .io_argOuts_12_bits(regs_io_argOuts_12_bits),
    .io_argOuts_13_valid(regs_io_argOuts_13_valid),
    .io_argOuts_13_bits(regs_io_argOuts_13_bits),
    .io_argOuts_14_valid(regs_io_argOuts_14_valid),
    .io_argOuts_14_bits(regs_io_argOuts_14_bits),
    .io_argOuts_15_valid(regs_io_argOuts_15_valid),
    .io_argOuts_15_bits(regs_io_argOuts_15_bits),
    .io_argOuts_16_valid(regs_io_argOuts_16_valid),
    .io_argOuts_16_bits(regs_io_argOuts_16_bits),
    .io_argOuts_17_valid(regs_io_argOuts_17_valid),
    .io_argOuts_17_bits(regs_io_argOuts_17_bits),
    .io_argOuts_18_valid(regs_io_argOuts_18_valid),
    .io_argOuts_18_bits(regs_io_argOuts_18_bits),
    .io_argOuts_19_valid(regs_io_argOuts_19_valid),
    .io_argOuts_19_bits(regs_io_argOuts_19_bits),
    .io_argOuts_20_valid(regs_io_argOuts_20_valid),
    .io_argOuts_20_bits(regs_io_argOuts_20_bits)
  );
  FringeCounter timeoutCtr ( // @[Fringe.scala 143:26:@53656.4]
    .clock(timeoutCtr_clock),
    .reset(timeoutCtr_reset),
    .io_enable(timeoutCtr_io_enable),
    .io_done(timeoutCtr_io_done)
  );
  Depulser depulser ( // @[Fringe.scala 153:24:@53674.4]
    .clock(depulser_clock),
    .reset(depulser_reset),
    .io_in(depulser_io_in),
    .io_rst(depulser_io_rst),
    .io_out(depulser_io_out)
  );
  assign _T_940 = regs_io_argIns_1; // @[:@53633.4 :@53634.4]
  assign curStatus_done = _T_940[0]; // @[Fringe.scala 133:45:@53635.4]
  assign curStatus_timeout = _T_940[1]; // @[Fringe.scala 133:45:@53637.4]
  assign curStatus_allocDealloc = _T_940[4:2]; // @[Fringe.scala 133:45:@53639.4]
  assign curStatus_sizeAddr = _T_940[63:5]; // @[Fringe.scala 133:45:@53641.4]
  assign _T_945 = regs_io_argIns_0[0]; // @[Fringe.scala 134:28:@53643.4]
  assign _T_949 = curStatus_done == 1'h0; // @[Fringe.scala 134:42:@53645.4]
  assign _T_950 = regs_io_argIns_0[1]; // @[Fringe.scala 135:27:@53647.4]
  assign _T_960 = ~ regs_io_argIns_0; // @[Fringe.scala 156:22:@53682.4]
  assign _T_968 = _T_967 ^ heap_io_host_0_req_valid; // @[package.scala 153:13:@53687.4]
  assign _T_969 = heap_io_host_0_req_valid & _T_968; // @[package.scala 153:8:@53688.4]
  assign _T_972 = _T_945 & depulser_io_out; // @[Fringe.scala 160:55:@53692.4]
  assign status_bits_done = depulser_io_out ? _T_972 : curStatus_done; // @[Fringe.scala 160:26:@53693.4]
  assign _T_975 = _T_945 & timeoutCtr_io_done; // @[Fringe.scala 161:58:@53696.4]
  assign status_bits_timeout = depulser_io_out ? _T_975 : curStatus_timeout; // @[Fringe.scala 161:29:@53697.4]
  assign _T_979 = heap_io_host_0_req_bits_allocDealloc ? 2'h1 : 2'h2; // @[Fringe.scala 162:57:@53699.4]
  assign _T_981 = heap_io_host_0_req_valid ? _T_979 : 2'h0; // @[Fringe.scala 162:34:@53700.4]
  assign _T_983 = heap_io_host_0_req_valid ? heap_io_host_0_req_bits_sizeAddr : 64'h0; // @[Fringe.scala 163:30:@53702.4]
  assign _T_984 = {status_bits_timeout,status_bits_done}; // @[Fringe.scala 171:37:@53705.4]
  assign status_bits_sizeAddr = _T_983[58:0]; // @[Fringe.scala 158:20:@53684.4 Fringe.scala 163:24:@53703.4]
  assign status_bits_allocDealloc = {{1'd0}, _T_981}; // @[Fringe.scala 158:20:@53684.4 Fringe.scala 162:28:@53701.4]
  assign _T_985 = {status_bits_sizeAddr,status_bits_allocDealloc}; // @[Fringe.scala 171:37:@53706.4]
  assign alloc = curStatus_allocDealloc == 3'h3; // @[Fringe.scala 202:38:@55048.4]
  assign dealloc = curStatus_allocDealloc == 3'h4; // @[Fringe.scala 203:40:@55049.4]
  assign _T_1489 = alloc | dealloc; // @[Fringe.scala 204:37:@55050.4]
  assign _T_1493 = _T_1492 ^ _T_1489; // @[package.scala 153:13:@55053.4]
  assign io_rdata = regs_io_rdata; // @[Fringe.scala 125:14:@53631.4]
  assign io_enable = _T_945 & _T_949; // @[Fringe.scala 136:13:@53651.4]
  assign io_reset = _T_950 | reset; // @[Fringe.scala 137:12:@53652.4]
  assign io_argIns_0 = regs_io_argIns_2; // @[Fringe.scala 151:51:@53673.4]
  assign io_heap_0_resp_valid = heap_io_accel_0_resp_valid; // @[Fringe.scala 108:17:@51527.4]
  assign io_heap_0_resp_bits_allocDealloc = heap_io_accel_0_resp_bits_allocDealloc; // @[Fringe.scala 108:17:@51526.4]
  assign io_heap_0_resp_bits_sizeAddr = heap_io_accel_0_resp_bits_sizeAddr; // @[Fringe.scala 108:17:@51525.4]
  assign heap_io_accel_0_req_valid = io_heap_0_req_valid; // @[Fringe.scala 108:17:@51530.4]
  assign heap_io_accel_0_req_bits_allocDealloc = io_heap_0_req_bits_allocDealloc; // @[Fringe.scala 108:17:@51529.4]
  assign heap_io_accel_0_req_bits_sizeAddr = io_heap_0_req_bits_sizeAddr; // @[Fringe.scala 108:17:@51528.4]
  assign heap_io_host_0_resp_valid = _T_1489 & _T_1493; // @[Fringe.scala 204:22:@55055.4]
  assign heap_io_host_0_resp_bits_allocDealloc = curStatus_allocDealloc == 3'h3; // @[Fringe.scala 205:34:@55056.4]
  assign heap_io_host_0_resp_bits_sizeAddr = {{5'd0}, curStatus_sizeAddr}; // @[Fringe.scala 206:30:@55057.4]
  assign regs_clock = clock; // @[:@51532.4]
  assign regs_reset = reset; // @[:@51533.4 Fringe.scala 139:14:@53655.4]
  assign regs_io_raddr = io_raddr; // @[Fringe.scala 118:17:@53627.4]
  assign regs_io_wen = io_wen; // @[Fringe.scala 120:15:@53629.4]
  assign regs_io_waddr = io_waddr; // @[Fringe.scala 119:17:@53628.4]
  assign regs_io_wdata = io_wdata; // @[Fringe.scala 121:17:@53630.4]
  assign regs_io_reset = _T_950 | reset; // @[Fringe.scala 138:17:@53653.4]
  assign regs_io_argOuts_0_valid = depulser_io_out | _T_969; // @[Fringe.scala 170:23:@53704.4]
  assign regs_io_argOuts_0_bits = {_T_985,_T_984}; // @[Fringe.scala 171:22:@53708.4]
  assign regs_io_argOuts_1_valid = io_argOuts_0_valid; // @[Fringe.scala 176:23:@53711.4]
  assign regs_io_argOuts_1_bits = io_argOuts_0_bits; // @[Fringe.scala 175:22:@53710.4]
  assign regs_io_argOuts_2_valid = io_argOuts_1_valid; // @[Fringe.scala 176:23:@53714.4]
  assign regs_io_argOuts_2_bits = io_argOuts_1_bits; // @[Fringe.scala 175:22:@53713.4]
  assign regs_io_argOuts_3_valid = io_argOuts_2_valid; // @[Fringe.scala 176:23:@53717.4]
  assign regs_io_argOuts_3_bits = io_argOuts_2_bits; // @[Fringe.scala 175:22:@53716.4]
  assign regs_io_argOuts_4_valid = io_argOuts_3_valid; // @[Fringe.scala 176:23:@53720.4]
  assign regs_io_argOuts_4_bits = io_argOuts_3_bits; // @[Fringe.scala 175:22:@53719.4]
  assign regs_io_argOuts_5_valid = io_argOuts_4_valid; // @[Fringe.scala 176:23:@53723.4]
  assign regs_io_argOuts_5_bits = io_argOuts_4_bits; // @[Fringe.scala 175:22:@53722.4]
  assign regs_io_argOuts_6_valid = io_argOuts_5_valid; // @[Fringe.scala 176:23:@53726.4]
  assign regs_io_argOuts_6_bits = io_argOuts_5_bits; // @[Fringe.scala 175:22:@53725.4]
  assign regs_io_argOuts_7_valid = io_argOuts_6_valid; // @[Fringe.scala 176:23:@53729.4]
  assign regs_io_argOuts_7_bits = io_argOuts_6_bits; // @[Fringe.scala 175:22:@53728.4]
  assign regs_io_argOuts_8_valid = io_argOuts_7_valid; // @[Fringe.scala 176:23:@53732.4]
  assign regs_io_argOuts_8_bits = io_argOuts_7_bits; // @[Fringe.scala 175:22:@53731.4]
  assign regs_io_argOuts_9_valid = io_argOuts_8_valid; // @[Fringe.scala 176:23:@53735.4]
  assign regs_io_argOuts_9_bits = io_argOuts_8_bits; // @[Fringe.scala 175:22:@53734.4]
  assign regs_io_argOuts_10_valid = io_argOuts_9_valid; // @[Fringe.scala 176:23:@53738.4]
  assign regs_io_argOuts_10_bits = io_argOuts_9_bits; // @[Fringe.scala 175:22:@53737.4]
  assign regs_io_argOuts_11_valid = io_argOuts_10_valid; // @[Fringe.scala 176:23:@53741.4]
  assign regs_io_argOuts_11_bits = io_argOuts_10_bits; // @[Fringe.scala 175:22:@53740.4]
  assign regs_io_argOuts_12_valid = io_argOuts_11_valid; // @[Fringe.scala 176:23:@53744.4]
  assign regs_io_argOuts_12_bits = io_argOuts_11_bits; // @[Fringe.scala 175:22:@53743.4]
  assign regs_io_argOuts_13_valid = io_argOuts_12_valid; // @[Fringe.scala 176:23:@53747.4]
  assign regs_io_argOuts_13_bits = io_argOuts_12_bits; // @[Fringe.scala 175:22:@53746.4]
  assign regs_io_argOuts_14_valid = io_argOuts_13_valid; // @[Fringe.scala 176:23:@53750.4]
  assign regs_io_argOuts_14_bits = io_argOuts_13_bits; // @[Fringe.scala 175:22:@53749.4]
  assign regs_io_argOuts_15_valid = io_argOuts_14_valid; // @[Fringe.scala 176:23:@53753.4]
  assign regs_io_argOuts_15_bits = io_argOuts_14_bits; // @[Fringe.scala 175:22:@53752.4]
  assign regs_io_argOuts_16_valid = io_argOuts_15_valid; // @[Fringe.scala 176:23:@53756.4]
  assign regs_io_argOuts_16_bits = io_argOuts_15_bits; // @[Fringe.scala 175:22:@53755.4]
  assign regs_io_argOuts_17_valid = io_argOuts_16_valid; // @[Fringe.scala 176:23:@53759.4]
  assign regs_io_argOuts_17_bits = io_argOuts_16_bits; // @[Fringe.scala 175:22:@53758.4]
  assign regs_io_argOuts_18_valid = io_argOuts_17_valid; // @[Fringe.scala 176:23:@53762.4]
  assign regs_io_argOuts_18_bits = io_argOuts_17_bits; // @[Fringe.scala 175:22:@53761.4]
  assign regs_io_argOuts_19_valid = io_argOuts_18_valid; // @[Fringe.scala 176:23:@53765.4]
  assign regs_io_argOuts_19_bits = io_argOuts_18_bits; // @[Fringe.scala 175:22:@53764.4]
  assign regs_io_argOuts_20_valid = io_argOuts_19_valid; // @[Fringe.scala 176:23:@53768.4]
  assign regs_io_argOuts_20_bits = io_argOuts_19_bits; // @[Fringe.scala 175:22:@53767.4]
  assign timeoutCtr_clock = clock; // @[:@53657.4]
  assign timeoutCtr_reset = reset; // @[:@53658.4]
  assign timeoutCtr_io_enable = _T_945 & _T_949; // @[Fringe.scala 149:24:@53672.4]
  assign depulser_clock = clock; // @[:@53675.4]
  assign depulser_reset = reset; // @[:@53676.4]
  assign depulser_io_in = io_done | timeoutCtr_io_done; // @[Fringe.scala 155:18:@53681.4]
  assign depulser_io_rst = _T_960[0]; // @[Fringe.scala 156:19:@53683.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_967 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1492 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_967 <= 1'h0;
    end else begin
      _T_967 <= heap_io_host_0_req_valid;
    end
    if (reset) begin
      _T_1492 <= 1'h0;
    end else begin
      _T_1492 <= _T_1489;
    end
  end
endmodule
module AXI4LiteToRFBridgeKCU1500( // @[:@55072.2]
  input         clock, // @[:@55073.4]
  input         reset, // @[:@55074.4]
  input  [31:0] io_S_AXI_AWADDR, // @[:@55075.4]
  input  [2:0]  io_S_AXI_AWPROT, // @[:@55075.4]
  input         io_S_AXI_AWVALID, // @[:@55075.4]
  output        io_S_AXI_AWREADY, // @[:@55075.4]
  input  [31:0] io_S_AXI_ARADDR, // @[:@55075.4]
  input  [2:0]  io_S_AXI_ARPROT, // @[:@55075.4]
  input         io_S_AXI_ARVALID, // @[:@55075.4]
  output        io_S_AXI_ARREADY, // @[:@55075.4]
  input  [31:0] io_S_AXI_WDATA, // @[:@55075.4]
  input  [3:0]  io_S_AXI_WSTRB, // @[:@55075.4]
  input         io_S_AXI_WVALID, // @[:@55075.4]
  output        io_S_AXI_WREADY, // @[:@55075.4]
  output [31:0] io_S_AXI_RDATA, // @[:@55075.4]
  output [1:0]  io_S_AXI_RRESP, // @[:@55075.4]
  output        io_S_AXI_RVALID, // @[:@55075.4]
  input         io_S_AXI_RREADY, // @[:@55075.4]
  output [1:0]  io_S_AXI_BRESP, // @[:@55075.4]
  output        io_S_AXI_BVALID, // @[:@55075.4]
  input         io_S_AXI_BREADY, // @[:@55075.4]
  output [31:0] io_raddr, // @[:@55075.4]
  output        io_wen, // @[:@55075.4]
  output [31:0] io_waddr, // @[:@55075.4]
  output [31:0] io_wdata, // @[:@55075.4]
  input  [31:0] io_rdata // @[:@55075.4]
);
  wire [31:0] d_rf_rdata; // @[AXI4LiteToRFBridge.scala 109:17:@55077.4]
  wire [31:0] d_rf_wdata; // @[AXI4LiteToRFBridge.scala 109:17:@55077.4]
  wire [31:0] d_rf_waddr; // @[AXI4LiteToRFBridge.scala 109:17:@55077.4]
  wire  d_rf_wen; // @[AXI4LiteToRFBridge.scala 109:17:@55077.4]
  wire [31:0] d_rf_raddr; // @[AXI4LiteToRFBridge.scala 109:17:@55077.4]
  wire  d_S_AXI_ARESETN; // @[AXI4LiteToRFBridge.scala 109:17:@55077.4]
  wire  d_S_AXI_ACLK; // @[AXI4LiteToRFBridge.scala 109:17:@55077.4]
  wire [31:0] d_S_AXI_AWADDR; // @[AXI4LiteToRFBridge.scala 109:17:@55077.4]
  wire [2:0] d_S_AXI_AWPROT; // @[AXI4LiteToRFBridge.scala 109:17:@55077.4]
  wire  d_S_AXI_AWVALID; // @[AXI4LiteToRFBridge.scala 109:17:@55077.4]
  wire  d_S_AXI_AWREADY; // @[AXI4LiteToRFBridge.scala 109:17:@55077.4]
  wire [31:0] d_S_AXI_ARADDR; // @[AXI4LiteToRFBridge.scala 109:17:@55077.4]
  wire [2:0] d_S_AXI_ARPROT; // @[AXI4LiteToRFBridge.scala 109:17:@55077.4]
  wire  d_S_AXI_ARVALID; // @[AXI4LiteToRFBridge.scala 109:17:@55077.4]
  wire  d_S_AXI_ARREADY; // @[AXI4LiteToRFBridge.scala 109:17:@55077.4]
  wire [31:0] d_S_AXI_WDATA; // @[AXI4LiteToRFBridge.scala 109:17:@55077.4]
  wire [3:0] d_S_AXI_WSTRB; // @[AXI4LiteToRFBridge.scala 109:17:@55077.4]
  wire  d_S_AXI_WVALID; // @[AXI4LiteToRFBridge.scala 109:17:@55077.4]
  wire  d_S_AXI_WREADY; // @[AXI4LiteToRFBridge.scala 109:17:@55077.4]
  wire [31:0] d_S_AXI_RDATA; // @[AXI4LiteToRFBridge.scala 109:17:@55077.4]
  wire [1:0] d_S_AXI_RRESP; // @[AXI4LiteToRFBridge.scala 109:17:@55077.4]
  wire  d_S_AXI_RVALID; // @[AXI4LiteToRFBridge.scala 109:17:@55077.4]
  wire  d_S_AXI_RREADY; // @[AXI4LiteToRFBridge.scala 109:17:@55077.4]
  wire [1:0] d_S_AXI_BRESP; // @[AXI4LiteToRFBridge.scala 109:17:@55077.4]
  wire  d_S_AXI_BVALID; // @[AXI4LiteToRFBridge.scala 109:17:@55077.4]
  wire  d_S_AXI_BREADY; // @[AXI4LiteToRFBridge.scala 109:17:@55077.4]
  AXI4LiteToRFBridgeVerilog d ( // @[AXI4LiteToRFBridge.scala 109:17:@55077.4]
    .rf_rdata(d_rf_rdata),
    .rf_wdata(d_rf_wdata),
    .rf_waddr(d_rf_waddr),
    .rf_wen(d_rf_wen),
    .rf_raddr(d_rf_raddr),
    .S_AXI_ARESETN(d_S_AXI_ARESETN),
    .S_AXI_ACLK(d_S_AXI_ACLK),
    .S_AXI_AWADDR(d_S_AXI_AWADDR),
    .S_AXI_AWPROT(d_S_AXI_AWPROT),
    .S_AXI_AWVALID(d_S_AXI_AWVALID),
    .S_AXI_AWREADY(d_S_AXI_AWREADY),
    .S_AXI_ARADDR(d_S_AXI_ARADDR),
    .S_AXI_ARPROT(d_S_AXI_ARPROT),
    .S_AXI_ARVALID(d_S_AXI_ARVALID),
    .S_AXI_ARREADY(d_S_AXI_ARREADY),
    .S_AXI_WDATA(d_S_AXI_WDATA),
    .S_AXI_WSTRB(d_S_AXI_WSTRB),
    .S_AXI_WVALID(d_S_AXI_WVALID),
    .S_AXI_WREADY(d_S_AXI_WREADY),
    .S_AXI_RDATA(d_S_AXI_RDATA),
    .S_AXI_RRESP(d_S_AXI_RRESP),
    .S_AXI_RVALID(d_S_AXI_RVALID),
    .S_AXI_RREADY(d_S_AXI_RREADY),
    .S_AXI_BRESP(d_S_AXI_BRESP),
    .S_AXI_BVALID(d_S_AXI_BVALID),
    .S_AXI_BREADY(d_S_AXI_BREADY)
  );
  assign io_S_AXI_AWREADY = d_S_AXI_AWREADY; // @[AXI4LiteToRFBridge.scala 111:14:@55101.4]
  assign io_S_AXI_ARREADY = d_S_AXI_ARREADY; // @[AXI4LiteToRFBridge.scala 111:14:@55097.4]
  assign io_S_AXI_WREADY = d_S_AXI_WREADY; // @[AXI4LiteToRFBridge.scala 111:14:@55093.4]
  assign io_S_AXI_RDATA = d_S_AXI_RDATA; // @[AXI4LiteToRFBridge.scala 111:14:@55092.4]
  assign io_S_AXI_RRESP = d_S_AXI_RRESP; // @[AXI4LiteToRFBridge.scala 111:14:@55091.4]
  assign io_S_AXI_RVALID = d_S_AXI_RVALID; // @[AXI4LiteToRFBridge.scala 111:14:@55090.4]
  assign io_S_AXI_BRESP = d_S_AXI_BRESP; // @[AXI4LiteToRFBridge.scala 111:14:@55088.4]
  assign io_S_AXI_BVALID = d_S_AXI_BVALID; // @[AXI4LiteToRFBridge.scala 111:14:@55087.4]
  assign io_raddr = d_rf_raddr; // @[AXI4LiteToRFBridge.scala 115:12:@55109.4]
  assign io_wen = d_rf_wen; // @[AXI4LiteToRFBridge.scala 118:12:@55112.4]
  assign io_waddr = d_rf_waddr; // @[AXI4LiteToRFBridge.scala 116:12:@55110.4]
  assign io_wdata = d_rf_wdata; // @[AXI4LiteToRFBridge.scala 117:12:@55111.4]
  assign d_rf_rdata = io_rdata; // @[AXI4LiteToRFBridge.scala 119:17:@55113.4]
  assign d_S_AXI_ARESETN = ~ reset; // @[AXI4LiteToRFBridge.scala 113:22:@55108.4]
  assign d_S_AXI_ACLK = clock; // @[AXI4LiteToRFBridge.scala 112:19:@55105.4]
  assign d_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[AXI4LiteToRFBridge.scala 111:14:@55104.4]
  assign d_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[AXI4LiteToRFBridge.scala 111:14:@55103.4]
  assign d_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[AXI4LiteToRFBridge.scala 111:14:@55102.4]
  assign d_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[AXI4LiteToRFBridge.scala 111:14:@55100.4]
  assign d_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[AXI4LiteToRFBridge.scala 111:14:@55099.4]
  assign d_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[AXI4LiteToRFBridge.scala 111:14:@55098.4]
  assign d_S_AXI_WDATA = io_S_AXI_WDATA; // @[AXI4LiteToRFBridge.scala 111:14:@55096.4]
  assign d_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[AXI4LiteToRFBridge.scala 111:14:@55095.4]
  assign d_S_AXI_WVALID = io_S_AXI_WVALID; // @[AXI4LiteToRFBridge.scala 111:14:@55094.4]
  assign d_S_AXI_RREADY = io_S_AXI_RREADY; // @[AXI4LiteToRFBridge.scala 111:14:@55089.4]
  assign d_S_AXI_BREADY = io_S_AXI_BREADY; // @[AXI4LiteToRFBridge.scala 111:14:@55086.4]
endmodule
module MAGToAXI4Bridge( // @[:@55115.2]
  output [7:0] io_M_AXI_AWLEN, // @[:@55118.4]
  output [7:0] io_M_AXI_ARLEN // @[:@55118.4]
);
  wire [32:0] _T_218; // @[MAGToAXI4Bridge.scala 27:29:@55275.4]
  wire [32:0] _T_219; // @[MAGToAXI4Bridge.scala 27:29:@55276.4]
  wire [31:0] _T_220; // @[MAGToAXI4Bridge.scala 27:29:@55277.4]
  assign _T_218 = 32'h0 - 32'h1; // @[MAGToAXI4Bridge.scala 27:29:@55275.4]
  assign _T_219 = $unsigned(_T_218); // @[MAGToAXI4Bridge.scala 27:29:@55276.4]
  assign _T_220 = _T_219[31:0]; // @[MAGToAXI4Bridge.scala 27:29:@55277.4]
  assign io_M_AXI_AWLEN = _T_220[7:0]; // @[MAGToAXI4Bridge.scala 41:21:@55295.4]
  assign io_M_AXI_ARLEN = _T_220[7:0]; // @[MAGToAXI4Bridge.scala 27:21:@55278.4]
endmodule
module FringeZynq( // @[:@55443.2]
  input         clock, // @[:@55444.4]
  input         reset, // @[:@55445.4]
  input  [31:0] io_S_AXI_AWADDR, // @[:@55446.4]
  input  [2:0]  io_S_AXI_AWPROT, // @[:@55446.4]
  input         io_S_AXI_AWVALID, // @[:@55446.4]
  output        io_S_AXI_AWREADY, // @[:@55446.4]
  input  [31:0] io_S_AXI_ARADDR, // @[:@55446.4]
  input  [2:0]  io_S_AXI_ARPROT, // @[:@55446.4]
  input         io_S_AXI_ARVALID, // @[:@55446.4]
  output        io_S_AXI_ARREADY, // @[:@55446.4]
  input  [31:0] io_S_AXI_WDATA, // @[:@55446.4]
  input  [3:0]  io_S_AXI_WSTRB, // @[:@55446.4]
  input         io_S_AXI_WVALID, // @[:@55446.4]
  output        io_S_AXI_WREADY, // @[:@55446.4]
  output [31:0] io_S_AXI_RDATA, // @[:@55446.4]
  output [1:0]  io_S_AXI_RRESP, // @[:@55446.4]
  output        io_S_AXI_RVALID, // @[:@55446.4]
  input         io_S_AXI_RREADY, // @[:@55446.4]
  output [1:0]  io_S_AXI_BRESP, // @[:@55446.4]
  output        io_S_AXI_BVALID, // @[:@55446.4]
  input         io_S_AXI_BREADY, // @[:@55446.4]
  output [7:0]  io_M_AXI_0_AWLEN, // @[:@55446.4]
  output [7:0]  io_M_AXI_0_ARLEN, // @[:@55446.4]
  output        io_enable, // @[:@55446.4]
  input         io_done, // @[:@55446.4]
  output        io_reset, // @[:@55446.4]
  output [63:0] io_argIns_0, // @[:@55446.4]
  input         io_argOuts_0_valid, // @[:@55446.4]
  input  [63:0] io_argOuts_0_bits, // @[:@55446.4]
  input         io_argOuts_1_valid, // @[:@55446.4]
  input  [63:0] io_argOuts_1_bits, // @[:@55446.4]
  input         io_argOuts_2_valid, // @[:@55446.4]
  input  [63:0] io_argOuts_2_bits, // @[:@55446.4]
  input         io_argOuts_3_valid, // @[:@55446.4]
  input  [63:0] io_argOuts_3_bits, // @[:@55446.4]
  input         io_argOuts_4_valid, // @[:@55446.4]
  input  [63:0] io_argOuts_4_bits, // @[:@55446.4]
  input         io_argOuts_5_valid, // @[:@55446.4]
  input  [63:0] io_argOuts_5_bits, // @[:@55446.4]
  input         io_argOuts_6_valid, // @[:@55446.4]
  input  [63:0] io_argOuts_6_bits, // @[:@55446.4]
  input         io_argOuts_7_valid, // @[:@55446.4]
  input  [63:0] io_argOuts_7_bits, // @[:@55446.4]
  input         io_argOuts_8_valid, // @[:@55446.4]
  input  [63:0] io_argOuts_8_bits, // @[:@55446.4]
  input         io_argOuts_9_valid, // @[:@55446.4]
  input  [63:0] io_argOuts_9_bits, // @[:@55446.4]
  input         io_argOuts_10_valid, // @[:@55446.4]
  input  [63:0] io_argOuts_10_bits, // @[:@55446.4]
  input         io_argOuts_11_valid, // @[:@55446.4]
  input  [63:0] io_argOuts_11_bits, // @[:@55446.4]
  input         io_argOuts_12_valid, // @[:@55446.4]
  input  [63:0] io_argOuts_12_bits, // @[:@55446.4]
  input         io_argOuts_13_valid, // @[:@55446.4]
  input  [63:0] io_argOuts_13_bits, // @[:@55446.4]
  input         io_argOuts_14_valid, // @[:@55446.4]
  input  [63:0] io_argOuts_14_bits, // @[:@55446.4]
  input         io_argOuts_15_valid, // @[:@55446.4]
  input  [63:0] io_argOuts_15_bits, // @[:@55446.4]
  input         io_argOuts_16_valid, // @[:@55446.4]
  input  [63:0] io_argOuts_16_bits, // @[:@55446.4]
  input         io_argOuts_17_valid, // @[:@55446.4]
  input  [63:0] io_argOuts_17_bits, // @[:@55446.4]
  input         io_argOuts_18_valid, // @[:@55446.4]
  input  [63:0] io_argOuts_18_bits, // @[:@55446.4]
  input         io_argOuts_19_valid, // @[:@55446.4]
  input  [63:0] io_argOuts_19_bits, // @[:@55446.4]
  input         io_heap_0_req_valid, // @[:@55446.4]
  input         io_heap_0_req_bits_allocDealloc, // @[:@55446.4]
  input  [63:0] io_heap_0_req_bits_sizeAddr, // @[:@55446.4]
  output        io_heap_0_resp_valid, // @[:@55446.4]
  output        io_heap_0_resp_bits_allocDealloc, // @[:@55446.4]
  output [63:0] io_heap_0_resp_bits_sizeAddr // @[:@55446.4]
);
  wire  fringeCommon_clock; // @[FringeZynq.scala 69:28:@55884.4]
  wire  fringeCommon_reset; // @[FringeZynq.scala 69:28:@55884.4]
  wire [31:0] fringeCommon_io_raddr; // @[FringeZynq.scala 69:28:@55884.4]
  wire  fringeCommon_io_wen; // @[FringeZynq.scala 69:28:@55884.4]
  wire [31:0] fringeCommon_io_waddr; // @[FringeZynq.scala 69:28:@55884.4]
  wire [63:0] fringeCommon_io_wdata; // @[FringeZynq.scala 69:28:@55884.4]
  wire [63:0] fringeCommon_io_rdata; // @[FringeZynq.scala 69:28:@55884.4]
  wire  fringeCommon_io_enable; // @[FringeZynq.scala 69:28:@55884.4]
  wire  fringeCommon_io_done; // @[FringeZynq.scala 69:28:@55884.4]
  wire  fringeCommon_io_reset; // @[FringeZynq.scala 69:28:@55884.4]
  wire [63:0] fringeCommon_io_argIns_0; // @[FringeZynq.scala 69:28:@55884.4]
  wire  fringeCommon_io_argOuts_0_valid; // @[FringeZynq.scala 69:28:@55884.4]
  wire [63:0] fringeCommon_io_argOuts_0_bits; // @[FringeZynq.scala 69:28:@55884.4]
  wire  fringeCommon_io_argOuts_1_valid; // @[FringeZynq.scala 69:28:@55884.4]
  wire [63:0] fringeCommon_io_argOuts_1_bits; // @[FringeZynq.scala 69:28:@55884.4]
  wire  fringeCommon_io_argOuts_2_valid; // @[FringeZynq.scala 69:28:@55884.4]
  wire [63:0] fringeCommon_io_argOuts_2_bits; // @[FringeZynq.scala 69:28:@55884.4]
  wire  fringeCommon_io_argOuts_3_valid; // @[FringeZynq.scala 69:28:@55884.4]
  wire [63:0] fringeCommon_io_argOuts_3_bits; // @[FringeZynq.scala 69:28:@55884.4]
  wire  fringeCommon_io_argOuts_4_valid; // @[FringeZynq.scala 69:28:@55884.4]
  wire [63:0] fringeCommon_io_argOuts_4_bits; // @[FringeZynq.scala 69:28:@55884.4]
  wire  fringeCommon_io_argOuts_5_valid; // @[FringeZynq.scala 69:28:@55884.4]
  wire [63:0] fringeCommon_io_argOuts_5_bits; // @[FringeZynq.scala 69:28:@55884.4]
  wire  fringeCommon_io_argOuts_6_valid; // @[FringeZynq.scala 69:28:@55884.4]
  wire [63:0] fringeCommon_io_argOuts_6_bits; // @[FringeZynq.scala 69:28:@55884.4]
  wire  fringeCommon_io_argOuts_7_valid; // @[FringeZynq.scala 69:28:@55884.4]
  wire [63:0] fringeCommon_io_argOuts_7_bits; // @[FringeZynq.scala 69:28:@55884.4]
  wire  fringeCommon_io_argOuts_8_valid; // @[FringeZynq.scala 69:28:@55884.4]
  wire [63:0] fringeCommon_io_argOuts_8_bits; // @[FringeZynq.scala 69:28:@55884.4]
  wire  fringeCommon_io_argOuts_9_valid; // @[FringeZynq.scala 69:28:@55884.4]
  wire [63:0] fringeCommon_io_argOuts_9_bits; // @[FringeZynq.scala 69:28:@55884.4]
  wire  fringeCommon_io_argOuts_10_valid; // @[FringeZynq.scala 69:28:@55884.4]
  wire [63:0] fringeCommon_io_argOuts_10_bits; // @[FringeZynq.scala 69:28:@55884.4]
  wire  fringeCommon_io_argOuts_11_valid; // @[FringeZynq.scala 69:28:@55884.4]
  wire [63:0] fringeCommon_io_argOuts_11_bits; // @[FringeZynq.scala 69:28:@55884.4]
  wire  fringeCommon_io_argOuts_12_valid; // @[FringeZynq.scala 69:28:@55884.4]
  wire [63:0] fringeCommon_io_argOuts_12_bits; // @[FringeZynq.scala 69:28:@55884.4]
  wire  fringeCommon_io_argOuts_13_valid; // @[FringeZynq.scala 69:28:@55884.4]
  wire [63:0] fringeCommon_io_argOuts_13_bits; // @[FringeZynq.scala 69:28:@55884.4]
  wire  fringeCommon_io_argOuts_14_valid; // @[FringeZynq.scala 69:28:@55884.4]
  wire [63:0] fringeCommon_io_argOuts_14_bits; // @[FringeZynq.scala 69:28:@55884.4]
  wire  fringeCommon_io_argOuts_15_valid; // @[FringeZynq.scala 69:28:@55884.4]
  wire [63:0] fringeCommon_io_argOuts_15_bits; // @[FringeZynq.scala 69:28:@55884.4]
  wire  fringeCommon_io_argOuts_16_valid; // @[FringeZynq.scala 69:28:@55884.4]
  wire [63:0] fringeCommon_io_argOuts_16_bits; // @[FringeZynq.scala 69:28:@55884.4]
  wire  fringeCommon_io_argOuts_17_valid; // @[FringeZynq.scala 69:28:@55884.4]
  wire [63:0] fringeCommon_io_argOuts_17_bits; // @[FringeZynq.scala 69:28:@55884.4]
  wire  fringeCommon_io_argOuts_18_valid; // @[FringeZynq.scala 69:28:@55884.4]
  wire [63:0] fringeCommon_io_argOuts_18_bits; // @[FringeZynq.scala 69:28:@55884.4]
  wire  fringeCommon_io_argOuts_19_valid; // @[FringeZynq.scala 69:28:@55884.4]
  wire [63:0] fringeCommon_io_argOuts_19_bits; // @[FringeZynq.scala 69:28:@55884.4]
  wire  fringeCommon_io_heap_0_req_valid; // @[FringeZynq.scala 69:28:@55884.4]
  wire  fringeCommon_io_heap_0_req_bits_allocDealloc; // @[FringeZynq.scala 69:28:@55884.4]
  wire [63:0] fringeCommon_io_heap_0_req_bits_sizeAddr; // @[FringeZynq.scala 69:28:@55884.4]
  wire  fringeCommon_io_heap_0_resp_valid; // @[FringeZynq.scala 69:28:@55884.4]
  wire  fringeCommon_io_heap_0_resp_bits_allocDealloc; // @[FringeZynq.scala 69:28:@55884.4]
  wire [63:0] fringeCommon_io_heap_0_resp_bits_sizeAddr; // @[FringeZynq.scala 69:28:@55884.4]
  wire  AXI4LiteToRFBridgeKCU1500_clock; // @[FringeZynq.scala 79:31:@56544.4]
  wire  AXI4LiteToRFBridgeKCU1500_reset; // @[FringeZynq.scala 79:31:@56544.4]
  wire [31:0] AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWADDR; // @[FringeZynq.scala 79:31:@56544.4]
  wire [2:0] AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWPROT; // @[FringeZynq.scala 79:31:@56544.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWVALID; // @[FringeZynq.scala 79:31:@56544.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWREADY; // @[FringeZynq.scala 79:31:@56544.4]
  wire [31:0] AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARADDR; // @[FringeZynq.scala 79:31:@56544.4]
  wire [2:0] AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARPROT; // @[FringeZynq.scala 79:31:@56544.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARVALID; // @[FringeZynq.scala 79:31:@56544.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARREADY; // @[FringeZynq.scala 79:31:@56544.4]
  wire [31:0] AXI4LiteToRFBridgeKCU1500_io_S_AXI_WDATA; // @[FringeZynq.scala 79:31:@56544.4]
  wire [3:0] AXI4LiteToRFBridgeKCU1500_io_S_AXI_WSTRB; // @[FringeZynq.scala 79:31:@56544.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_WVALID; // @[FringeZynq.scala 79:31:@56544.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_WREADY; // @[FringeZynq.scala 79:31:@56544.4]
  wire [31:0] AXI4LiteToRFBridgeKCU1500_io_S_AXI_RDATA; // @[FringeZynq.scala 79:31:@56544.4]
  wire [1:0] AXI4LiteToRFBridgeKCU1500_io_S_AXI_RRESP; // @[FringeZynq.scala 79:31:@56544.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_RVALID; // @[FringeZynq.scala 79:31:@56544.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_RREADY; // @[FringeZynq.scala 79:31:@56544.4]
  wire [1:0] AXI4LiteToRFBridgeKCU1500_io_S_AXI_BRESP; // @[FringeZynq.scala 79:31:@56544.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_BVALID; // @[FringeZynq.scala 79:31:@56544.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_BREADY; // @[FringeZynq.scala 79:31:@56544.4]
  wire [31:0] AXI4LiteToRFBridgeKCU1500_io_raddr; // @[FringeZynq.scala 79:31:@56544.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_wen; // @[FringeZynq.scala 79:31:@56544.4]
  wire [31:0] AXI4LiteToRFBridgeKCU1500_io_waddr; // @[FringeZynq.scala 79:31:@56544.4]
  wire [31:0] AXI4LiteToRFBridgeKCU1500_io_wdata; // @[FringeZynq.scala 79:31:@56544.4]
  wire [31:0] AXI4LiteToRFBridgeKCU1500_io_rdata; // @[FringeZynq.scala 79:31:@56544.4]
  wire [7:0] MAGToAXI4Bridge_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@56767.4]
  wire [7:0] MAGToAXI4Bridge_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@56767.4]
  Fringe fringeCommon ( // @[FringeZynq.scala 69:28:@55884.4]
    .clock(fringeCommon_clock),
    .reset(fringeCommon_reset),
    .io_raddr(fringeCommon_io_raddr),
    .io_wen(fringeCommon_io_wen),
    .io_waddr(fringeCommon_io_waddr),
    .io_wdata(fringeCommon_io_wdata),
    .io_rdata(fringeCommon_io_rdata),
    .io_enable(fringeCommon_io_enable),
    .io_done(fringeCommon_io_done),
    .io_reset(fringeCommon_io_reset),
    .io_argIns_0(fringeCommon_io_argIns_0),
    .io_argOuts_0_valid(fringeCommon_io_argOuts_0_valid),
    .io_argOuts_0_bits(fringeCommon_io_argOuts_0_bits),
    .io_argOuts_1_valid(fringeCommon_io_argOuts_1_valid),
    .io_argOuts_1_bits(fringeCommon_io_argOuts_1_bits),
    .io_argOuts_2_valid(fringeCommon_io_argOuts_2_valid),
    .io_argOuts_2_bits(fringeCommon_io_argOuts_2_bits),
    .io_argOuts_3_valid(fringeCommon_io_argOuts_3_valid),
    .io_argOuts_3_bits(fringeCommon_io_argOuts_3_bits),
    .io_argOuts_4_valid(fringeCommon_io_argOuts_4_valid),
    .io_argOuts_4_bits(fringeCommon_io_argOuts_4_bits),
    .io_argOuts_5_valid(fringeCommon_io_argOuts_5_valid),
    .io_argOuts_5_bits(fringeCommon_io_argOuts_5_bits),
    .io_argOuts_6_valid(fringeCommon_io_argOuts_6_valid),
    .io_argOuts_6_bits(fringeCommon_io_argOuts_6_bits),
    .io_argOuts_7_valid(fringeCommon_io_argOuts_7_valid),
    .io_argOuts_7_bits(fringeCommon_io_argOuts_7_bits),
    .io_argOuts_8_valid(fringeCommon_io_argOuts_8_valid),
    .io_argOuts_8_bits(fringeCommon_io_argOuts_8_bits),
    .io_argOuts_9_valid(fringeCommon_io_argOuts_9_valid),
    .io_argOuts_9_bits(fringeCommon_io_argOuts_9_bits),
    .io_argOuts_10_valid(fringeCommon_io_argOuts_10_valid),
    .io_argOuts_10_bits(fringeCommon_io_argOuts_10_bits),
    .io_argOuts_11_valid(fringeCommon_io_argOuts_11_valid),
    .io_argOuts_11_bits(fringeCommon_io_argOuts_11_bits),
    .io_argOuts_12_valid(fringeCommon_io_argOuts_12_valid),
    .io_argOuts_12_bits(fringeCommon_io_argOuts_12_bits),
    .io_argOuts_13_valid(fringeCommon_io_argOuts_13_valid),
    .io_argOuts_13_bits(fringeCommon_io_argOuts_13_bits),
    .io_argOuts_14_valid(fringeCommon_io_argOuts_14_valid),
    .io_argOuts_14_bits(fringeCommon_io_argOuts_14_bits),
    .io_argOuts_15_valid(fringeCommon_io_argOuts_15_valid),
    .io_argOuts_15_bits(fringeCommon_io_argOuts_15_bits),
    .io_argOuts_16_valid(fringeCommon_io_argOuts_16_valid),
    .io_argOuts_16_bits(fringeCommon_io_argOuts_16_bits),
    .io_argOuts_17_valid(fringeCommon_io_argOuts_17_valid),
    .io_argOuts_17_bits(fringeCommon_io_argOuts_17_bits),
    .io_argOuts_18_valid(fringeCommon_io_argOuts_18_valid),
    .io_argOuts_18_bits(fringeCommon_io_argOuts_18_bits),
    .io_argOuts_19_valid(fringeCommon_io_argOuts_19_valid),
    .io_argOuts_19_bits(fringeCommon_io_argOuts_19_bits),
    .io_heap_0_req_valid(fringeCommon_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(fringeCommon_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(fringeCommon_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(fringeCommon_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(fringeCommon_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(fringeCommon_io_heap_0_resp_bits_sizeAddr)
  );
  AXI4LiteToRFBridgeKCU1500 AXI4LiteToRFBridgeKCU1500 ( // @[FringeZynq.scala 79:31:@56544.4]
    .clock(AXI4LiteToRFBridgeKCU1500_clock),
    .reset(AXI4LiteToRFBridgeKCU1500_reset),
    .io_S_AXI_AWADDR(AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWADDR),
    .io_S_AXI_AWPROT(AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWPROT),
    .io_S_AXI_AWVALID(AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWVALID),
    .io_S_AXI_AWREADY(AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWREADY),
    .io_S_AXI_ARADDR(AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARADDR),
    .io_S_AXI_ARPROT(AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARPROT),
    .io_S_AXI_ARVALID(AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARVALID),
    .io_S_AXI_ARREADY(AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARREADY),
    .io_S_AXI_WDATA(AXI4LiteToRFBridgeKCU1500_io_S_AXI_WDATA),
    .io_S_AXI_WSTRB(AXI4LiteToRFBridgeKCU1500_io_S_AXI_WSTRB),
    .io_S_AXI_WVALID(AXI4LiteToRFBridgeKCU1500_io_S_AXI_WVALID),
    .io_S_AXI_WREADY(AXI4LiteToRFBridgeKCU1500_io_S_AXI_WREADY),
    .io_S_AXI_RDATA(AXI4LiteToRFBridgeKCU1500_io_S_AXI_RDATA),
    .io_S_AXI_RRESP(AXI4LiteToRFBridgeKCU1500_io_S_AXI_RRESP),
    .io_S_AXI_RVALID(AXI4LiteToRFBridgeKCU1500_io_S_AXI_RVALID),
    .io_S_AXI_RREADY(AXI4LiteToRFBridgeKCU1500_io_S_AXI_RREADY),
    .io_S_AXI_BRESP(AXI4LiteToRFBridgeKCU1500_io_S_AXI_BRESP),
    .io_S_AXI_BVALID(AXI4LiteToRFBridgeKCU1500_io_S_AXI_BVALID),
    .io_S_AXI_BREADY(AXI4LiteToRFBridgeKCU1500_io_S_AXI_BREADY),
    .io_raddr(AXI4LiteToRFBridgeKCU1500_io_raddr),
    .io_wen(AXI4LiteToRFBridgeKCU1500_io_wen),
    .io_waddr(AXI4LiteToRFBridgeKCU1500_io_waddr),
    .io_wdata(AXI4LiteToRFBridgeKCU1500_io_wdata),
    .io_rdata(AXI4LiteToRFBridgeKCU1500_io_rdata)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge ( // @[FringeZynq.scala 131:27:@56767.4]
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_io_M_AXI_AWLEN),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_io_M_AXI_ARLEN)
  );
  assign io_S_AXI_AWREADY = AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWREADY; // @[FringeZynq.scala 80:28:@56562.4]
  assign io_S_AXI_ARREADY = AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARREADY; // @[FringeZynq.scala 80:28:@56558.4]
  assign io_S_AXI_WREADY = AXI4LiteToRFBridgeKCU1500_io_S_AXI_WREADY; // @[FringeZynq.scala 80:28:@56554.4]
  assign io_S_AXI_RDATA = AXI4LiteToRFBridgeKCU1500_io_S_AXI_RDATA; // @[FringeZynq.scala 80:28:@56553.4]
  assign io_S_AXI_RRESP = AXI4LiteToRFBridgeKCU1500_io_S_AXI_RRESP; // @[FringeZynq.scala 80:28:@56552.4]
  assign io_S_AXI_RVALID = AXI4LiteToRFBridgeKCU1500_io_S_AXI_RVALID; // @[FringeZynq.scala 80:28:@56551.4]
  assign io_S_AXI_BRESP = AXI4LiteToRFBridgeKCU1500_io_S_AXI_BRESP; // @[FringeZynq.scala 80:28:@56549.4]
  assign io_S_AXI_BVALID = AXI4LiteToRFBridgeKCU1500_io_S_AXI_BVALID; // @[FringeZynq.scala 80:28:@56548.4]
  assign io_M_AXI_0_AWLEN = MAGToAXI4Bridge_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@56919.4]
  assign io_M_AXI_0_ARLEN = MAGToAXI4Bridge_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@56907.4]
  assign io_enable = fringeCommon_io_enable; // @[FringeZynq.scala 115:13:@56574.4]
  assign io_reset = fringeCommon_io_reset; // @[FringeZynq.scala 119:12:@56578.4]
  assign io_argIns_0 = fringeCommon_io_argIns_0; // @[FringeZynq.scala 121:13:@56579.4]
  assign io_heap_0_resp_valid = fringeCommon_io_heap_0_resp_valid; // @[FringeZynq.scala 127:11:@56763.4]
  assign io_heap_0_resp_bits_allocDealloc = fringeCommon_io_heap_0_resp_bits_allocDealloc; // @[FringeZynq.scala 127:11:@56762.4]
  assign io_heap_0_resp_bits_sizeAddr = fringeCommon_io_heap_0_resp_bits_sizeAddr; // @[FringeZynq.scala 127:11:@56761.4]
  assign fringeCommon_clock = clock; // @[:@55885.4]
  assign fringeCommon_reset = reset; // @[:@55886.4 FringeZynq.scala 82:24:@56567.4 FringeZynq.scala 117:22:@56577.4]
  assign fringeCommon_io_raddr = AXI4LiteToRFBridgeKCU1500_io_raddr; // @[FringeZynq.scala 83:27:@56568.4]
  assign fringeCommon_io_wen = AXI4LiteToRFBridgeKCU1500_io_wen; // @[FringeZynq.scala 84:27:@56569.4]
  assign fringeCommon_io_waddr = AXI4LiteToRFBridgeKCU1500_io_waddr; // @[FringeZynq.scala 85:27:@56570.4]
  assign fringeCommon_io_wdata = {{32'd0}, AXI4LiteToRFBridgeKCU1500_io_wdata}; // @[FringeZynq.scala 86:27:@56571.4]
  assign fringeCommon_io_done = io_done; // @[FringeZynq.scala 116:24:@56575.4]
  assign fringeCommon_io_argOuts_0_valid = io_argOuts_0_valid; // @[FringeZynq.scala 122:27:@56581.4]
  assign fringeCommon_io_argOuts_0_bits = io_argOuts_0_bits; // @[FringeZynq.scala 122:27:@56580.4]
  assign fringeCommon_io_argOuts_1_valid = io_argOuts_1_valid; // @[FringeZynq.scala 122:27:@56584.4]
  assign fringeCommon_io_argOuts_1_bits = io_argOuts_1_bits; // @[FringeZynq.scala 122:27:@56583.4]
  assign fringeCommon_io_argOuts_2_valid = io_argOuts_2_valid; // @[FringeZynq.scala 122:27:@56587.4]
  assign fringeCommon_io_argOuts_2_bits = io_argOuts_2_bits; // @[FringeZynq.scala 122:27:@56586.4]
  assign fringeCommon_io_argOuts_3_valid = io_argOuts_3_valid; // @[FringeZynq.scala 122:27:@56590.4]
  assign fringeCommon_io_argOuts_3_bits = io_argOuts_3_bits; // @[FringeZynq.scala 122:27:@56589.4]
  assign fringeCommon_io_argOuts_4_valid = io_argOuts_4_valid; // @[FringeZynq.scala 122:27:@56593.4]
  assign fringeCommon_io_argOuts_4_bits = io_argOuts_4_bits; // @[FringeZynq.scala 122:27:@56592.4]
  assign fringeCommon_io_argOuts_5_valid = io_argOuts_5_valid; // @[FringeZynq.scala 122:27:@56596.4]
  assign fringeCommon_io_argOuts_5_bits = io_argOuts_5_bits; // @[FringeZynq.scala 122:27:@56595.4]
  assign fringeCommon_io_argOuts_6_valid = io_argOuts_6_valid; // @[FringeZynq.scala 122:27:@56599.4]
  assign fringeCommon_io_argOuts_6_bits = io_argOuts_6_bits; // @[FringeZynq.scala 122:27:@56598.4]
  assign fringeCommon_io_argOuts_7_valid = io_argOuts_7_valid; // @[FringeZynq.scala 122:27:@56602.4]
  assign fringeCommon_io_argOuts_7_bits = io_argOuts_7_bits; // @[FringeZynq.scala 122:27:@56601.4]
  assign fringeCommon_io_argOuts_8_valid = io_argOuts_8_valid; // @[FringeZynq.scala 122:27:@56605.4]
  assign fringeCommon_io_argOuts_8_bits = io_argOuts_8_bits; // @[FringeZynq.scala 122:27:@56604.4]
  assign fringeCommon_io_argOuts_9_valid = io_argOuts_9_valid; // @[FringeZynq.scala 122:27:@56608.4]
  assign fringeCommon_io_argOuts_9_bits = io_argOuts_9_bits; // @[FringeZynq.scala 122:27:@56607.4]
  assign fringeCommon_io_argOuts_10_valid = io_argOuts_10_valid; // @[FringeZynq.scala 122:27:@56611.4]
  assign fringeCommon_io_argOuts_10_bits = io_argOuts_10_bits; // @[FringeZynq.scala 122:27:@56610.4]
  assign fringeCommon_io_argOuts_11_valid = io_argOuts_11_valid; // @[FringeZynq.scala 122:27:@56614.4]
  assign fringeCommon_io_argOuts_11_bits = io_argOuts_11_bits; // @[FringeZynq.scala 122:27:@56613.4]
  assign fringeCommon_io_argOuts_12_valid = io_argOuts_12_valid; // @[FringeZynq.scala 122:27:@56617.4]
  assign fringeCommon_io_argOuts_12_bits = io_argOuts_12_bits; // @[FringeZynq.scala 122:27:@56616.4]
  assign fringeCommon_io_argOuts_13_valid = io_argOuts_13_valid; // @[FringeZynq.scala 122:27:@56620.4]
  assign fringeCommon_io_argOuts_13_bits = io_argOuts_13_bits; // @[FringeZynq.scala 122:27:@56619.4]
  assign fringeCommon_io_argOuts_14_valid = io_argOuts_14_valid; // @[FringeZynq.scala 122:27:@56623.4]
  assign fringeCommon_io_argOuts_14_bits = io_argOuts_14_bits; // @[FringeZynq.scala 122:27:@56622.4]
  assign fringeCommon_io_argOuts_15_valid = io_argOuts_15_valid; // @[FringeZynq.scala 122:27:@56626.4]
  assign fringeCommon_io_argOuts_15_bits = io_argOuts_15_bits; // @[FringeZynq.scala 122:27:@56625.4]
  assign fringeCommon_io_argOuts_16_valid = io_argOuts_16_valid; // @[FringeZynq.scala 122:27:@56629.4]
  assign fringeCommon_io_argOuts_16_bits = io_argOuts_16_bits; // @[FringeZynq.scala 122:27:@56628.4]
  assign fringeCommon_io_argOuts_17_valid = io_argOuts_17_valid; // @[FringeZynq.scala 122:27:@56632.4]
  assign fringeCommon_io_argOuts_17_bits = io_argOuts_17_bits; // @[FringeZynq.scala 122:27:@56631.4]
  assign fringeCommon_io_argOuts_18_valid = io_argOuts_18_valid; // @[FringeZynq.scala 122:27:@56635.4]
  assign fringeCommon_io_argOuts_18_bits = io_argOuts_18_bits; // @[FringeZynq.scala 122:27:@56634.4]
  assign fringeCommon_io_argOuts_19_valid = io_argOuts_19_valid; // @[FringeZynq.scala 122:27:@56638.4]
  assign fringeCommon_io_argOuts_19_bits = io_argOuts_19_bits; // @[FringeZynq.scala 122:27:@56637.4]
  assign fringeCommon_io_heap_0_req_valid = io_heap_0_req_valid; // @[FringeZynq.scala 127:11:@56766.4]
  assign fringeCommon_io_heap_0_req_bits_allocDealloc = io_heap_0_req_bits_allocDealloc; // @[FringeZynq.scala 127:11:@56765.4]
  assign fringeCommon_io_heap_0_req_bits_sizeAddr = io_heap_0_req_bits_sizeAddr; // @[FringeZynq.scala 127:11:@56764.4]
  assign AXI4LiteToRFBridgeKCU1500_clock = clock; // @[:@56545.4]
  assign AXI4LiteToRFBridgeKCU1500_reset = reset; // @[:@56546.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[FringeZynq.scala 80:28:@56565.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[FringeZynq.scala 80:28:@56564.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[FringeZynq.scala 80:28:@56563.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[FringeZynq.scala 80:28:@56561.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[FringeZynq.scala 80:28:@56560.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[FringeZynq.scala 80:28:@56559.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_WDATA = io_S_AXI_WDATA; // @[FringeZynq.scala 80:28:@56557.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[FringeZynq.scala 80:28:@56556.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_WVALID = io_S_AXI_WVALID; // @[FringeZynq.scala 80:28:@56555.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_RREADY = io_S_AXI_RREADY; // @[FringeZynq.scala 80:28:@56550.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_BREADY = io_S_AXI_BREADY; // @[FringeZynq.scala 80:28:@56547.4]
  assign AXI4LiteToRFBridgeKCU1500_io_rdata = fringeCommon_io_rdata[31:0]; // @[FringeZynq.scala 87:28:@56572.4]
endmodule
module SpatialIP( // @[:@56926.2]
  input          clock, // @[:@56927.4]
  input          reset, // @[:@56928.4]
  input          io_raddr, // @[:@56929.4]
  input          io_wen, // @[:@56929.4]
  input          io_waddr, // @[:@56929.4]
  input          io_wdata, // @[:@56929.4]
  output         io_rdata, // @[:@56929.4]
  input  [31:0]  io_S_AXI_AWADDR, // @[:@56929.4]
  input  [2:0]   io_S_AXI_AWPROT, // @[:@56929.4]
  input          io_S_AXI_AWVALID, // @[:@56929.4]
  output         io_S_AXI_AWREADY, // @[:@56929.4]
  input  [31:0]  io_S_AXI_ARADDR, // @[:@56929.4]
  input  [2:0]   io_S_AXI_ARPROT, // @[:@56929.4]
  input          io_S_AXI_ARVALID, // @[:@56929.4]
  output         io_S_AXI_ARREADY, // @[:@56929.4]
  input  [31:0]  io_S_AXI_WDATA, // @[:@56929.4]
  input  [3:0]   io_S_AXI_WSTRB, // @[:@56929.4]
  input          io_S_AXI_WVALID, // @[:@56929.4]
  output         io_S_AXI_WREADY, // @[:@56929.4]
  output [31:0]  io_S_AXI_RDATA, // @[:@56929.4]
  output [1:0]   io_S_AXI_RRESP, // @[:@56929.4]
  output         io_S_AXI_RVALID, // @[:@56929.4]
  input          io_S_AXI_RREADY, // @[:@56929.4]
  output [1:0]   io_S_AXI_BRESP, // @[:@56929.4]
  output         io_S_AXI_BVALID, // @[:@56929.4]
  input          io_S_AXI_BREADY, // @[:@56929.4]
  output [3:0]   io_M_AXI_0_AWID, // @[:@56929.4]
  output [3:0]   io_M_AXI_0_AWUSER, // @[:@56929.4]
  output [31:0]  io_M_AXI_0_AWADDR, // @[:@56929.4]
  output [7:0]   io_M_AXI_0_AWLEN, // @[:@56929.4]
  output [2:0]   io_M_AXI_0_AWSIZE, // @[:@56929.4]
  output [1:0]   io_M_AXI_0_AWBURST, // @[:@56929.4]
  output         io_M_AXI_0_AWLOCK, // @[:@56929.4]
  output [3:0]   io_M_AXI_0_AWCACHE, // @[:@56929.4]
  output [2:0]   io_M_AXI_0_AWPROT, // @[:@56929.4]
  output [3:0]   io_M_AXI_0_AWQOS, // @[:@56929.4]
  output         io_M_AXI_0_AWVALID, // @[:@56929.4]
  input          io_M_AXI_0_AWREADY, // @[:@56929.4]
  output [3:0]   io_M_AXI_0_ARID, // @[:@56929.4]
  output [3:0]   io_M_AXI_0_ARUSER, // @[:@56929.4]
  output [31:0]  io_M_AXI_0_ARADDR, // @[:@56929.4]
  output [7:0]   io_M_AXI_0_ARLEN, // @[:@56929.4]
  output [2:0]   io_M_AXI_0_ARSIZE, // @[:@56929.4]
  output [1:0]   io_M_AXI_0_ARBURST, // @[:@56929.4]
  output         io_M_AXI_0_ARLOCK, // @[:@56929.4]
  output [3:0]   io_M_AXI_0_ARCACHE, // @[:@56929.4]
  output [2:0]   io_M_AXI_0_ARPROT, // @[:@56929.4]
  output [3:0]   io_M_AXI_0_ARQOS, // @[:@56929.4]
  output         io_M_AXI_0_ARVALID, // @[:@56929.4]
  input          io_M_AXI_0_ARREADY, // @[:@56929.4]
  output [511:0] io_M_AXI_0_WDATA, // @[:@56929.4]
  output [63:0]  io_M_AXI_0_WSTRB, // @[:@56929.4]
  output         io_M_AXI_0_WLAST, // @[:@56929.4]
  output         io_M_AXI_0_WVALID, // @[:@56929.4]
  input          io_M_AXI_0_WREADY, // @[:@56929.4]
  input  [3:0]   io_M_AXI_0_RID, // @[:@56929.4]
  input  [31:0]  io_M_AXI_0_RUSER, // @[:@56929.4]
  input  [511:0] io_M_AXI_0_RDATA, // @[:@56929.4]
  input  [1:0]   io_M_AXI_0_RRESP, // @[:@56929.4]
  input          io_M_AXI_0_RLAST, // @[:@56929.4]
  input          io_M_AXI_0_RVALID, // @[:@56929.4]
  output         io_M_AXI_0_RREADY, // @[:@56929.4]
  input  [3:0]   io_M_AXI_0_BID, // @[:@56929.4]
  input  [3:0]   io_M_AXI_0_BUSER, // @[:@56929.4]
  input  [1:0]   io_M_AXI_0_BRESP, // @[:@56929.4]
  input          io_M_AXI_0_BVALID, // @[:@56929.4]
  output         io_M_AXI_0_BREADY, // @[:@56929.4]
  input          io_AXIS_IN_TVALID, // @[:@56929.4]
  output         io_AXIS_IN_TREADY, // @[:@56929.4]
  input  [63:0]  io_AXIS_IN_TDATA, // @[:@56929.4]
  input  [7:0]   io_AXIS_IN_TSTRB, // @[:@56929.4]
  input  [7:0]   io_AXIS_IN_TKEEP, // @[:@56929.4]
  input          io_AXIS_IN_TLAST, // @[:@56929.4]
  input  [7:0]   io_AXIS_IN_TID, // @[:@56929.4]
  input  [7:0]   io_AXIS_IN_TDEST, // @[:@56929.4]
  input  [63:0]  io_AXIS_IN_TUSER, // @[:@56929.4]
  output         io_AXIS_OUT_TVALID, // @[:@56929.4]
  input          io_AXIS_OUT_TREADY, // @[:@56929.4]
  output [63:0]  io_AXIS_OUT_TDATA, // @[:@56929.4]
  output [7:0]   io_AXIS_OUT_TSTRB, // @[:@56929.4]
  output [7:0]   io_AXIS_OUT_TKEEP, // @[:@56929.4]
  output         io_AXIS_OUT_TLAST, // @[:@56929.4]
  output [7:0]   io_AXIS_OUT_TID, // @[:@56929.4]
  output [7:0]   io_AXIS_OUT_TDEST, // @[:@56929.4]
  output [63:0]  io_AXIS_OUT_TUSER // @[:@56929.4]
);
  wire  accel_clock; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_reset; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_enable; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_done; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_reset; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_memStreams_loads_0_cmd_ready; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_memStreams_loads_0_cmd_valid; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_memStreams_loads_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_loads_0_cmd_bits_size; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_memStreams_loads_0_data_ready; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_memStreams_loads_0_data_valid; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_0; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_1; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_2; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_3; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_4; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_5; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_6; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_7; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_8; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_9; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_10; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_11; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_12; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_13; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_14; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_15; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_memStreams_stores_0_cmd_ready; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_memStreams_stores_0_cmd_valid; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_memStreams_stores_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_stores_0_cmd_bits_size; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_memStreams_stores_0_data_ready; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_memStreams_stores_0_data_valid; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_0; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_1; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_2; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_3; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_4; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_5; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_6; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_7; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_8; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_9; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_10; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_11; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_12; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_13; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_14; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_15; // @[Instantiator.scala 53:44:@56931.4]
  wire [15:0] accel_io_memStreams_stores_0_data_bits_wstrb; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_memStreams_stores_0_wresp_ready; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_memStreams_stores_0_wresp_valid; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_memStreams_stores_0_wresp_bits; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_memStreams_gathers_0_cmd_ready; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_memStreams_gathers_0_cmd_valid; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_0; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_1; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_2; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_3; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_4; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_5; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_6; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_7; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_8; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_9; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_10; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_11; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_12; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_13; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_14; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_15; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_memStreams_gathers_0_data_ready; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_memStreams_gathers_0_data_valid; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_0; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_1; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_2; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_3; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_4; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_5; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_6; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_7; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_8; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_9; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_10; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_11; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_12; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_13; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_14; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_15; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_memStreams_scatters_0_cmd_ready; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_memStreams_scatters_0_cmd_valid; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_0; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_1; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_2; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_3; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_4; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_5; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_6; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_7; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_8; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_9; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_10; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_11; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_12; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_13; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_14; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_15; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_memStreams_scatters_0_wresp_ready; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_memStreams_scatters_0_wresp_valid; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_memStreams_scatters_0_wresp_bits; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_axiStreamsIn_0_TVALID; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_axiStreamsIn_0_TREADY; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_axiStreamsIn_0_TDATA; // @[Instantiator.scala 53:44:@56931.4]
  wire [7:0] accel_io_axiStreamsIn_0_TSTRB; // @[Instantiator.scala 53:44:@56931.4]
  wire [7:0] accel_io_axiStreamsIn_0_TKEEP; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_axiStreamsIn_0_TLAST; // @[Instantiator.scala 53:44:@56931.4]
  wire [7:0] accel_io_axiStreamsIn_0_TID; // @[Instantiator.scala 53:44:@56931.4]
  wire [7:0] accel_io_axiStreamsIn_0_TDEST; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_axiStreamsIn_0_TUSER; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_axiStreamsOut_0_TVALID; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_axiStreamsOut_0_TREADY; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_axiStreamsOut_0_TDATA; // @[Instantiator.scala 53:44:@56931.4]
  wire [7:0] accel_io_axiStreamsOut_0_TSTRB; // @[Instantiator.scala 53:44:@56931.4]
  wire [7:0] accel_io_axiStreamsOut_0_TKEEP; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_axiStreamsOut_0_TLAST; // @[Instantiator.scala 53:44:@56931.4]
  wire [7:0] accel_io_axiStreamsOut_0_TID; // @[Instantiator.scala 53:44:@56931.4]
  wire [7:0] accel_io_axiStreamsOut_0_TDEST; // @[Instantiator.scala 53:44:@56931.4]
  wire [31:0] accel_io_axiStreamsOut_0_TUSER; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_heap_0_req_valid; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_heap_0_req_bits_allocDealloc; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_heap_0_req_bits_sizeAddr; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_heap_0_resp_valid; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_heap_0_resp_bits_allocDealloc; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_heap_0_resp_bits_sizeAddr; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_argIns_0; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_argOuts_0_port_ready; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_argOuts_0_port_valid; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_argOuts_0_port_bits; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_argOuts_0_echo; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_argOuts_1_port_ready; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_argOuts_1_port_valid; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_argOuts_1_port_bits; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_argOuts_1_echo; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_argOuts_2_port_ready; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_argOuts_2_port_valid; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_argOuts_2_port_bits; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_argOuts_2_echo; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_argOuts_3_port_ready; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_argOuts_3_port_valid; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_argOuts_3_port_bits; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_argOuts_3_echo; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_argOuts_4_port_ready; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_argOuts_4_port_valid; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_argOuts_4_port_bits; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_argOuts_4_echo; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_argOuts_5_port_ready; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_argOuts_5_port_valid; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_argOuts_5_port_bits; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_argOuts_5_echo; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_argOuts_6_port_ready; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_argOuts_6_port_valid; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_argOuts_6_port_bits; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_argOuts_6_echo; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_argOuts_7_port_ready; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_argOuts_7_port_valid; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_argOuts_7_port_bits; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_argOuts_7_echo; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_argOuts_8_port_ready; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_argOuts_8_port_valid; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_argOuts_8_port_bits; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_argOuts_8_echo; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_argOuts_9_port_ready; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_argOuts_9_port_valid; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_argOuts_9_port_bits; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_argOuts_9_echo; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_argOuts_10_port_ready; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_argOuts_10_port_valid; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_argOuts_10_port_bits; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_argOuts_10_echo; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_argOuts_11_port_ready; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_argOuts_11_port_valid; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_argOuts_11_port_bits; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_argOuts_11_echo; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_argOuts_12_port_ready; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_argOuts_12_port_valid; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_argOuts_12_port_bits; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_argOuts_12_echo; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_argOuts_13_port_ready; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_argOuts_13_port_valid; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_argOuts_13_port_bits; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_argOuts_13_echo; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_argOuts_14_port_ready; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_argOuts_14_port_valid; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_argOuts_14_port_bits; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_argOuts_14_echo; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_argOuts_15_port_ready; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_argOuts_15_port_valid; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_argOuts_15_port_bits; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_argOuts_15_echo; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_argOuts_16_port_ready; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_argOuts_16_port_valid; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_argOuts_16_port_bits; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_argOuts_16_echo; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_argOuts_17_port_ready; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_argOuts_17_port_valid; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_argOuts_17_port_bits; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_argOuts_17_echo; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_argOuts_18_port_ready; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_argOuts_18_port_valid; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_argOuts_18_port_bits; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_argOuts_18_echo; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_argOuts_19_port_ready; // @[Instantiator.scala 53:44:@56931.4]
  wire  accel_io_argOuts_19_port_valid; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_argOuts_19_port_bits; // @[Instantiator.scala 53:44:@56931.4]
  wire [63:0] accel_io_argOuts_19_echo; // @[Instantiator.scala 53:44:@56931.4]
  wire  FringeZynq_clock; // @[KCU1500.scala 21:24:@57163.4]
  wire  FringeZynq_reset; // @[KCU1500.scala 21:24:@57163.4]
  wire [31:0] FringeZynq_io_S_AXI_AWADDR; // @[KCU1500.scala 21:24:@57163.4]
  wire [2:0] FringeZynq_io_S_AXI_AWPROT; // @[KCU1500.scala 21:24:@57163.4]
  wire  FringeZynq_io_S_AXI_AWVALID; // @[KCU1500.scala 21:24:@57163.4]
  wire  FringeZynq_io_S_AXI_AWREADY; // @[KCU1500.scala 21:24:@57163.4]
  wire [31:0] FringeZynq_io_S_AXI_ARADDR; // @[KCU1500.scala 21:24:@57163.4]
  wire [2:0] FringeZynq_io_S_AXI_ARPROT; // @[KCU1500.scala 21:24:@57163.4]
  wire  FringeZynq_io_S_AXI_ARVALID; // @[KCU1500.scala 21:24:@57163.4]
  wire  FringeZynq_io_S_AXI_ARREADY; // @[KCU1500.scala 21:24:@57163.4]
  wire [31:0] FringeZynq_io_S_AXI_WDATA; // @[KCU1500.scala 21:24:@57163.4]
  wire [3:0] FringeZynq_io_S_AXI_WSTRB; // @[KCU1500.scala 21:24:@57163.4]
  wire  FringeZynq_io_S_AXI_WVALID; // @[KCU1500.scala 21:24:@57163.4]
  wire  FringeZynq_io_S_AXI_WREADY; // @[KCU1500.scala 21:24:@57163.4]
  wire [31:0] FringeZynq_io_S_AXI_RDATA; // @[KCU1500.scala 21:24:@57163.4]
  wire [1:0] FringeZynq_io_S_AXI_RRESP; // @[KCU1500.scala 21:24:@57163.4]
  wire  FringeZynq_io_S_AXI_RVALID; // @[KCU1500.scala 21:24:@57163.4]
  wire  FringeZynq_io_S_AXI_RREADY; // @[KCU1500.scala 21:24:@57163.4]
  wire [1:0] FringeZynq_io_S_AXI_BRESP; // @[KCU1500.scala 21:24:@57163.4]
  wire  FringeZynq_io_S_AXI_BVALID; // @[KCU1500.scala 21:24:@57163.4]
  wire  FringeZynq_io_S_AXI_BREADY; // @[KCU1500.scala 21:24:@57163.4]
  wire [7:0] FringeZynq_io_M_AXI_0_AWLEN; // @[KCU1500.scala 21:24:@57163.4]
  wire [7:0] FringeZynq_io_M_AXI_0_ARLEN; // @[KCU1500.scala 21:24:@57163.4]
  wire  FringeZynq_io_enable; // @[KCU1500.scala 21:24:@57163.4]
  wire  FringeZynq_io_done; // @[KCU1500.scala 21:24:@57163.4]
  wire  FringeZynq_io_reset; // @[KCU1500.scala 21:24:@57163.4]
  wire [63:0] FringeZynq_io_argIns_0; // @[KCU1500.scala 21:24:@57163.4]
  wire  FringeZynq_io_argOuts_0_valid; // @[KCU1500.scala 21:24:@57163.4]
  wire [63:0] FringeZynq_io_argOuts_0_bits; // @[KCU1500.scala 21:24:@57163.4]
  wire  FringeZynq_io_argOuts_1_valid; // @[KCU1500.scala 21:24:@57163.4]
  wire [63:0] FringeZynq_io_argOuts_1_bits; // @[KCU1500.scala 21:24:@57163.4]
  wire  FringeZynq_io_argOuts_2_valid; // @[KCU1500.scala 21:24:@57163.4]
  wire [63:0] FringeZynq_io_argOuts_2_bits; // @[KCU1500.scala 21:24:@57163.4]
  wire  FringeZynq_io_argOuts_3_valid; // @[KCU1500.scala 21:24:@57163.4]
  wire [63:0] FringeZynq_io_argOuts_3_bits; // @[KCU1500.scala 21:24:@57163.4]
  wire  FringeZynq_io_argOuts_4_valid; // @[KCU1500.scala 21:24:@57163.4]
  wire [63:0] FringeZynq_io_argOuts_4_bits; // @[KCU1500.scala 21:24:@57163.4]
  wire  FringeZynq_io_argOuts_5_valid; // @[KCU1500.scala 21:24:@57163.4]
  wire [63:0] FringeZynq_io_argOuts_5_bits; // @[KCU1500.scala 21:24:@57163.4]
  wire  FringeZynq_io_argOuts_6_valid; // @[KCU1500.scala 21:24:@57163.4]
  wire [63:0] FringeZynq_io_argOuts_6_bits; // @[KCU1500.scala 21:24:@57163.4]
  wire  FringeZynq_io_argOuts_7_valid; // @[KCU1500.scala 21:24:@57163.4]
  wire [63:0] FringeZynq_io_argOuts_7_bits; // @[KCU1500.scala 21:24:@57163.4]
  wire  FringeZynq_io_argOuts_8_valid; // @[KCU1500.scala 21:24:@57163.4]
  wire [63:0] FringeZynq_io_argOuts_8_bits; // @[KCU1500.scala 21:24:@57163.4]
  wire  FringeZynq_io_argOuts_9_valid; // @[KCU1500.scala 21:24:@57163.4]
  wire [63:0] FringeZynq_io_argOuts_9_bits; // @[KCU1500.scala 21:24:@57163.4]
  wire  FringeZynq_io_argOuts_10_valid; // @[KCU1500.scala 21:24:@57163.4]
  wire [63:0] FringeZynq_io_argOuts_10_bits; // @[KCU1500.scala 21:24:@57163.4]
  wire  FringeZynq_io_argOuts_11_valid; // @[KCU1500.scala 21:24:@57163.4]
  wire [63:0] FringeZynq_io_argOuts_11_bits; // @[KCU1500.scala 21:24:@57163.4]
  wire  FringeZynq_io_argOuts_12_valid; // @[KCU1500.scala 21:24:@57163.4]
  wire [63:0] FringeZynq_io_argOuts_12_bits; // @[KCU1500.scala 21:24:@57163.4]
  wire  FringeZynq_io_argOuts_13_valid; // @[KCU1500.scala 21:24:@57163.4]
  wire [63:0] FringeZynq_io_argOuts_13_bits; // @[KCU1500.scala 21:24:@57163.4]
  wire  FringeZynq_io_argOuts_14_valid; // @[KCU1500.scala 21:24:@57163.4]
  wire [63:0] FringeZynq_io_argOuts_14_bits; // @[KCU1500.scala 21:24:@57163.4]
  wire  FringeZynq_io_argOuts_15_valid; // @[KCU1500.scala 21:24:@57163.4]
  wire [63:0] FringeZynq_io_argOuts_15_bits; // @[KCU1500.scala 21:24:@57163.4]
  wire  FringeZynq_io_argOuts_16_valid; // @[KCU1500.scala 21:24:@57163.4]
  wire [63:0] FringeZynq_io_argOuts_16_bits; // @[KCU1500.scala 21:24:@57163.4]
  wire  FringeZynq_io_argOuts_17_valid; // @[KCU1500.scala 21:24:@57163.4]
  wire [63:0] FringeZynq_io_argOuts_17_bits; // @[KCU1500.scala 21:24:@57163.4]
  wire  FringeZynq_io_argOuts_18_valid; // @[KCU1500.scala 21:24:@57163.4]
  wire [63:0] FringeZynq_io_argOuts_18_bits; // @[KCU1500.scala 21:24:@57163.4]
  wire  FringeZynq_io_argOuts_19_valid; // @[KCU1500.scala 21:24:@57163.4]
  wire [63:0] FringeZynq_io_argOuts_19_bits; // @[KCU1500.scala 21:24:@57163.4]
  wire  FringeZynq_io_heap_0_req_valid; // @[KCU1500.scala 21:24:@57163.4]
  wire  FringeZynq_io_heap_0_req_bits_allocDealloc; // @[KCU1500.scala 21:24:@57163.4]
  wire [63:0] FringeZynq_io_heap_0_req_bits_sizeAddr; // @[KCU1500.scala 21:24:@57163.4]
  wire  FringeZynq_io_heap_0_resp_valid; // @[KCU1500.scala 21:24:@57163.4]
  wire  FringeZynq_io_heap_0_resp_bits_allocDealloc; // @[KCU1500.scala 21:24:@57163.4]
  wire [63:0] FringeZynq_io_heap_0_resp_bits_sizeAddr; // @[KCU1500.scala 21:24:@57163.4]
  AccelUnit accel ( // @[Instantiator.scala 53:44:@56931.4]
    .clock(accel_clock),
    .reset(accel_reset),
    .io_enable(accel_io_enable),
    .io_done(accel_io_done),
    .io_reset(accel_io_reset),
    .io_memStreams_loads_0_cmd_ready(accel_io_memStreams_loads_0_cmd_ready),
    .io_memStreams_loads_0_cmd_valid(accel_io_memStreams_loads_0_cmd_valid),
    .io_memStreams_loads_0_cmd_bits_addr(accel_io_memStreams_loads_0_cmd_bits_addr),
    .io_memStreams_loads_0_cmd_bits_size(accel_io_memStreams_loads_0_cmd_bits_size),
    .io_memStreams_loads_0_data_ready(accel_io_memStreams_loads_0_data_ready),
    .io_memStreams_loads_0_data_valid(accel_io_memStreams_loads_0_data_valid),
    .io_memStreams_loads_0_data_bits_rdata_0(accel_io_memStreams_loads_0_data_bits_rdata_0),
    .io_memStreams_loads_0_data_bits_rdata_1(accel_io_memStreams_loads_0_data_bits_rdata_1),
    .io_memStreams_loads_0_data_bits_rdata_2(accel_io_memStreams_loads_0_data_bits_rdata_2),
    .io_memStreams_loads_0_data_bits_rdata_3(accel_io_memStreams_loads_0_data_bits_rdata_3),
    .io_memStreams_loads_0_data_bits_rdata_4(accel_io_memStreams_loads_0_data_bits_rdata_4),
    .io_memStreams_loads_0_data_bits_rdata_5(accel_io_memStreams_loads_0_data_bits_rdata_5),
    .io_memStreams_loads_0_data_bits_rdata_6(accel_io_memStreams_loads_0_data_bits_rdata_6),
    .io_memStreams_loads_0_data_bits_rdata_7(accel_io_memStreams_loads_0_data_bits_rdata_7),
    .io_memStreams_loads_0_data_bits_rdata_8(accel_io_memStreams_loads_0_data_bits_rdata_8),
    .io_memStreams_loads_0_data_bits_rdata_9(accel_io_memStreams_loads_0_data_bits_rdata_9),
    .io_memStreams_loads_0_data_bits_rdata_10(accel_io_memStreams_loads_0_data_bits_rdata_10),
    .io_memStreams_loads_0_data_bits_rdata_11(accel_io_memStreams_loads_0_data_bits_rdata_11),
    .io_memStreams_loads_0_data_bits_rdata_12(accel_io_memStreams_loads_0_data_bits_rdata_12),
    .io_memStreams_loads_0_data_bits_rdata_13(accel_io_memStreams_loads_0_data_bits_rdata_13),
    .io_memStreams_loads_0_data_bits_rdata_14(accel_io_memStreams_loads_0_data_bits_rdata_14),
    .io_memStreams_loads_0_data_bits_rdata_15(accel_io_memStreams_loads_0_data_bits_rdata_15),
    .io_memStreams_stores_0_cmd_ready(accel_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(accel_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(accel_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(accel_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(accel_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(accel_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(accel_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wdata_1(accel_io_memStreams_stores_0_data_bits_wdata_1),
    .io_memStreams_stores_0_data_bits_wdata_2(accel_io_memStreams_stores_0_data_bits_wdata_2),
    .io_memStreams_stores_0_data_bits_wdata_3(accel_io_memStreams_stores_0_data_bits_wdata_3),
    .io_memStreams_stores_0_data_bits_wdata_4(accel_io_memStreams_stores_0_data_bits_wdata_4),
    .io_memStreams_stores_0_data_bits_wdata_5(accel_io_memStreams_stores_0_data_bits_wdata_5),
    .io_memStreams_stores_0_data_bits_wdata_6(accel_io_memStreams_stores_0_data_bits_wdata_6),
    .io_memStreams_stores_0_data_bits_wdata_7(accel_io_memStreams_stores_0_data_bits_wdata_7),
    .io_memStreams_stores_0_data_bits_wdata_8(accel_io_memStreams_stores_0_data_bits_wdata_8),
    .io_memStreams_stores_0_data_bits_wdata_9(accel_io_memStreams_stores_0_data_bits_wdata_9),
    .io_memStreams_stores_0_data_bits_wdata_10(accel_io_memStreams_stores_0_data_bits_wdata_10),
    .io_memStreams_stores_0_data_bits_wdata_11(accel_io_memStreams_stores_0_data_bits_wdata_11),
    .io_memStreams_stores_0_data_bits_wdata_12(accel_io_memStreams_stores_0_data_bits_wdata_12),
    .io_memStreams_stores_0_data_bits_wdata_13(accel_io_memStreams_stores_0_data_bits_wdata_13),
    .io_memStreams_stores_0_data_bits_wdata_14(accel_io_memStreams_stores_0_data_bits_wdata_14),
    .io_memStreams_stores_0_data_bits_wdata_15(accel_io_memStreams_stores_0_data_bits_wdata_15),
    .io_memStreams_stores_0_data_bits_wstrb(accel_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(accel_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(accel_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(accel_io_memStreams_stores_0_wresp_bits),
    .io_memStreams_gathers_0_cmd_ready(accel_io_memStreams_gathers_0_cmd_ready),
    .io_memStreams_gathers_0_cmd_valid(accel_io_memStreams_gathers_0_cmd_valid),
    .io_memStreams_gathers_0_cmd_bits_addr_0(accel_io_memStreams_gathers_0_cmd_bits_addr_0),
    .io_memStreams_gathers_0_cmd_bits_addr_1(accel_io_memStreams_gathers_0_cmd_bits_addr_1),
    .io_memStreams_gathers_0_cmd_bits_addr_2(accel_io_memStreams_gathers_0_cmd_bits_addr_2),
    .io_memStreams_gathers_0_cmd_bits_addr_3(accel_io_memStreams_gathers_0_cmd_bits_addr_3),
    .io_memStreams_gathers_0_cmd_bits_addr_4(accel_io_memStreams_gathers_0_cmd_bits_addr_4),
    .io_memStreams_gathers_0_cmd_bits_addr_5(accel_io_memStreams_gathers_0_cmd_bits_addr_5),
    .io_memStreams_gathers_0_cmd_bits_addr_6(accel_io_memStreams_gathers_0_cmd_bits_addr_6),
    .io_memStreams_gathers_0_cmd_bits_addr_7(accel_io_memStreams_gathers_0_cmd_bits_addr_7),
    .io_memStreams_gathers_0_cmd_bits_addr_8(accel_io_memStreams_gathers_0_cmd_bits_addr_8),
    .io_memStreams_gathers_0_cmd_bits_addr_9(accel_io_memStreams_gathers_0_cmd_bits_addr_9),
    .io_memStreams_gathers_0_cmd_bits_addr_10(accel_io_memStreams_gathers_0_cmd_bits_addr_10),
    .io_memStreams_gathers_0_cmd_bits_addr_11(accel_io_memStreams_gathers_0_cmd_bits_addr_11),
    .io_memStreams_gathers_0_cmd_bits_addr_12(accel_io_memStreams_gathers_0_cmd_bits_addr_12),
    .io_memStreams_gathers_0_cmd_bits_addr_13(accel_io_memStreams_gathers_0_cmd_bits_addr_13),
    .io_memStreams_gathers_0_cmd_bits_addr_14(accel_io_memStreams_gathers_0_cmd_bits_addr_14),
    .io_memStreams_gathers_0_cmd_bits_addr_15(accel_io_memStreams_gathers_0_cmd_bits_addr_15),
    .io_memStreams_gathers_0_data_ready(accel_io_memStreams_gathers_0_data_ready),
    .io_memStreams_gathers_0_data_valid(accel_io_memStreams_gathers_0_data_valid),
    .io_memStreams_gathers_0_data_bits_0(accel_io_memStreams_gathers_0_data_bits_0),
    .io_memStreams_gathers_0_data_bits_1(accel_io_memStreams_gathers_0_data_bits_1),
    .io_memStreams_gathers_0_data_bits_2(accel_io_memStreams_gathers_0_data_bits_2),
    .io_memStreams_gathers_0_data_bits_3(accel_io_memStreams_gathers_0_data_bits_3),
    .io_memStreams_gathers_0_data_bits_4(accel_io_memStreams_gathers_0_data_bits_4),
    .io_memStreams_gathers_0_data_bits_5(accel_io_memStreams_gathers_0_data_bits_5),
    .io_memStreams_gathers_0_data_bits_6(accel_io_memStreams_gathers_0_data_bits_6),
    .io_memStreams_gathers_0_data_bits_7(accel_io_memStreams_gathers_0_data_bits_7),
    .io_memStreams_gathers_0_data_bits_8(accel_io_memStreams_gathers_0_data_bits_8),
    .io_memStreams_gathers_0_data_bits_9(accel_io_memStreams_gathers_0_data_bits_9),
    .io_memStreams_gathers_0_data_bits_10(accel_io_memStreams_gathers_0_data_bits_10),
    .io_memStreams_gathers_0_data_bits_11(accel_io_memStreams_gathers_0_data_bits_11),
    .io_memStreams_gathers_0_data_bits_12(accel_io_memStreams_gathers_0_data_bits_12),
    .io_memStreams_gathers_0_data_bits_13(accel_io_memStreams_gathers_0_data_bits_13),
    .io_memStreams_gathers_0_data_bits_14(accel_io_memStreams_gathers_0_data_bits_14),
    .io_memStreams_gathers_0_data_bits_15(accel_io_memStreams_gathers_0_data_bits_15),
    .io_memStreams_scatters_0_cmd_ready(accel_io_memStreams_scatters_0_cmd_ready),
    .io_memStreams_scatters_0_cmd_valid(accel_io_memStreams_scatters_0_cmd_valid),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_0(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_1(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_2(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_3(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_4(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_5(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_6(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_7(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_8(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_9(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_10(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_11(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_12(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_13(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_14(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_15(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15),
    .io_memStreams_scatters_0_cmd_bits_wdata_0(accel_io_memStreams_scatters_0_cmd_bits_wdata_0),
    .io_memStreams_scatters_0_cmd_bits_wdata_1(accel_io_memStreams_scatters_0_cmd_bits_wdata_1),
    .io_memStreams_scatters_0_cmd_bits_wdata_2(accel_io_memStreams_scatters_0_cmd_bits_wdata_2),
    .io_memStreams_scatters_0_cmd_bits_wdata_3(accel_io_memStreams_scatters_0_cmd_bits_wdata_3),
    .io_memStreams_scatters_0_cmd_bits_wdata_4(accel_io_memStreams_scatters_0_cmd_bits_wdata_4),
    .io_memStreams_scatters_0_cmd_bits_wdata_5(accel_io_memStreams_scatters_0_cmd_bits_wdata_5),
    .io_memStreams_scatters_0_cmd_bits_wdata_6(accel_io_memStreams_scatters_0_cmd_bits_wdata_6),
    .io_memStreams_scatters_0_cmd_bits_wdata_7(accel_io_memStreams_scatters_0_cmd_bits_wdata_7),
    .io_memStreams_scatters_0_cmd_bits_wdata_8(accel_io_memStreams_scatters_0_cmd_bits_wdata_8),
    .io_memStreams_scatters_0_cmd_bits_wdata_9(accel_io_memStreams_scatters_0_cmd_bits_wdata_9),
    .io_memStreams_scatters_0_cmd_bits_wdata_10(accel_io_memStreams_scatters_0_cmd_bits_wdata_10),
    .io_memStreams_scatters_0_cmd_bits_wdata_11(accel_io_memStreams_scatters_0_cmd_bits_wdata_11),
    .io_memStreams_scatters_0_cmd_bits_wdata_12(accel_io_memStreams_scatters_0_cmd_bits_wdata_12),
    .io_memStreams_scatters_0_cmd_bits_wdata_13(accel_io_memStreams_scatters_0_cmd_bits_wdata_13),
    .io_memStreams_scatters_0_cmd_bits_wdata_14(accel_io_memStreams_scatters_0_cmd_bits_wdata_14),
    .io_memStreams_scatters_0_cmd_bits_wdata_15(accel_io_memStreams_scatters_0_cmd_bits_wdata_15),
    .io_memStreams_scatters_0_wresp_ready(accel_io_memStreams_scatters_0_wresp_ready),
    .io_memStreams_scatters_0_wresp_valid(accel_io_memStreams_scatters_0_wresp_valid),
    .io_memStreams_scatters_0_wresp_bits(accel_io_memStreams_scatters_0_wresp_bits),
    .io_axiStreamsIn_0_TVALID(accel_io_axiStreamsIn_0_TVALID),
    .io_axiStreamsIn_0_TREADY(accel_io_axiStreamsIn_0_TREADY),
    .io_axiStreamsIn_0_TDATA(accel_io_axiStreamsIn_0_TDATA),
    .io_axiStreamsIn_0_TSTRB(accel_io_axiStreamsIn_0_TSTRB),
    .io_axiStreamsIn_0_TKEEP(accel_io_axiStreamsIn_0_TKEEP),
    .io_axiStreamsIn_0_TLAST(accel_io_axiStreamsIn_0_TLAST),
    .io_axiStreamsIn_0_TID(accel_io_axiStreamsIn_0_TID),
    .io_axiStreamsIn_0_TDEST(accel_io_axiStreamsIn_0_TDEST),
    .io_axiStreamsIn_0_TUSER(accel_io_axiStreamsIn_0_TUSER),
    .io_axiStreamsOut_0_TVALID(accel_io_axiStreamsOut_0_TVALID),
    .io_axiStreamsOut_0_TREADY(accel_io_axiStreamsOut_0_TREADY),
    .io_axiStreamsOut_0_TDATA(accel_io_axiStreamsOut_0_TDATA),
    .io_axiStreamsOut_0_TSTRB(accel_io_axiStreamsOut_0_TSTRB),
    .io_axiStreamsOut_0_TKEEP(accel_io_axiStreamsOut_0_TKEEP),
    .io_axiStreamsOut_0_TLAST(accel_io_axiStreamsOut_0_TLAST),
    .io_axiStreamsOut_0_TID(accel_io_axiStreamsOut_0_TID),
    .io_axiStreamsOut_0_TDEST(accel_io_axiStreamsOut_0_TDEST),
    .io_axiStreamsOut_0_TUSER(accel_io_axiStreamsOut_0_TUSER),
    .io_heap_0_req_valid(accel_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(accel_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(accel_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(accel_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(accel_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(accel_io_heap_0_resp_bits_sizeAddr),
    .io_argIns_0(accel_io_argIns_0),
    .io_argOuts_0_port_ready(accel_io_argOuts_0_port_ready),
    .io_argOuts_0_port_valid(accel_io_argOuts_0_port_valid),
    .io_argOuts_0_port_bits(accel_io_argOuts_0_port_bits),
    .io_argOuts_0_echo(accel_io_argOuts_0_echo),
    .io_argOuts_1_port_ready(accel_io_argOuts_1_port_ready),
    .io_argOuts_1_port_valid(accel_io_argOuts_1_port_valid),
    .io_argOuts_1_port_bits(accel_io_argOuts_1_port_bits),
    .io_argOuts_1_echo(accel_io_argOuts_1_echo),
    .io_argOuts_2_port_ready(accel_io_argOuts_2_port_ready),
    .io_argOuts_2_port_valid(accel_io_argOuts_2_port_valid),
    .io_argOuts_2_port_bits(accel_io_argOuts_2_port_bits),
    .io_argOuts_2_echo(accel_io_argOuts_2_echo),
    .io_argOuts_3_port_ready(accel_io_argOuts_3_port_ready),
    .io_argOuts_3_port_valid(accel_io_argOuts_3_port_valid),
    .io_argOuts_3_port_bits(accel_io_argOuts_3_port_bits),
    .io_argOuts_3_echo(accel_io_argOuts_3_echo),
    .io_argOuts_4_port_ready(accel_io_argOuts_4_port_ready),
    .io_argOuts_4_port_valid(accel_io_argOuts_4_port_valid),
    .io_argOuts_4_port_bits(accel_io_argOuts_4_port_bits),
    .io_argOuts_4_echo(accel_io_argOuts_4_echo),
    .io_argOuts_5_port_ready(accel_io_argOuts_5_port_ready),
    .io_argOuts_5_port_valid(accel_io_argOuts_5_port_valid),
    .io_argOuts_5_port_bits(accel_io_argOuts_5_port_bits),
    .io_argOuts_5_echo(accel_io_argOuts_5_echo),
    .io_argOuts_6_port_ready(accel_io_argOuts_6_port_ready),
    .io_argOuts_6_port_valid(accel_io_argOuts_6_port_valid),
    .io_argOuts_6_port_bits(accel_io_argOuts_6_port_bits),
    .io_argOuts_6_echo(accel_io_argOuts_6_echo),
    .io_argOuts_7_port_ready(accel_io_argOuts_7_port_ready),
    .io_argOuts_7_port_valid(accel_io_argOuts_7_port_valid),
    .io_argOuts_7_port_bits(accel_io_argOuts_7_port_bits),
    .io_argOuts_7_echo(accel_io_argOuts_7_echo),
    .io_argOuts_8_port_ready(accel_io_argOuts_8_port_ready),
    .io_argOuts_8_port_valid(accel_io_argOuts_8_port_valid),
    .io_argOuts_8_port_bits(accel_io_argOuts_8_port_bits),
    .io_argOuts_8_echo(accel_io_argOuts_8_echo),
    .io_argOuts_9_port_ready(accel_io_argOuts_9_port_ready),
    .io_argOuts_9_port_valid(accel_io_argOuts_9_port_valid),
    .io_argOuts_9_port_bits(accel_io_argOuts_9_port_bits),
    .io_argOuts_9_echo(accel_io_argOuts_9_echo),
    .io_argOuts_10_port_ready(accel_io_argOuts_10_port_ready),
    .io_argOuts_10_port_valid(accel_io_argOuts_10_port_valid),
    .io_argOuts_10_port_bits(accel_io_argOuts_10_port_bits),
    .io_argOuts_10_echo(accel_io_argOuts_10_echo),
    .io_argOuts_11_port_ready(accel_io_argOuts_11_port_ready),
    .io_argOuts_11_port_valid(accel_io_argOuts_11_port_valid),
    .io_argOuts_11_port_bits(accel_io_argOuts_11_port_bits),
    .io_argOuts_11_echo(accel_io_argOuts_11_echo),
    .io_argOuts_12_port_ready(accel_io_argOuts_12_port_ready),
    .io_argOuts_12_port_valid(accel_io_argOuts_12_port_valid),
    .io_argOuts_12_port_bits(accel_io_argOuts_12_port_bits),
    .io_argOuts_12_echo(accel_io_argOuts_12_echo),
    .io_argOuts_13_port_ready(accel_io_argOuts_13_port_ready),
    .io_argOuts_13_port_valid(accel_io_argOuts_13_port_valid),
    .io_argOuts_13_port_bits(accel_io_argOuts_13_port_bits),
    .io_argOuts_13_echo(accel_io_argOuts_13_echo),
    .io_argOuts_14_port_ready(accel_io_argOuts_14_port_ready),
    .io_argOuts_14_port_valid(accel_io_argOuts_14_port_valid),
    .io_argOuts_14_port_bits(accel_io_argOuts_14_port_bits),
    .io_argOuts_14_echo(accel_io_argOuts_14_echo),
    .io_argOuts_15_port_ready(accel_io_argOuts_15_port_ready),
    .io_argOuts_15_port_valid(accel_io_argOuts_15_port_valid),
    .io_argOuts_15_port_bits(accel_io_argOuts_15_port_bits),
    .io_argOuts_15_echo(accel_io_argOuts_15_echo),
    .io_argOuts_16_port_ready(accel_io_argOuts_16_port_ready),
    .io_argOuts_16_port_valid(accel_io_argOuts_16_port_valid),
    .io_argOuts_16_port_bits(accel_io_argOuts_16_port_bits),
    .io_argOuts_16_echo(accel_io_argOuts_16_echo),
    .io_argOuts_17_port_ready(accel_io_argOuts_17_port_ready),
    .io_argOuts_17_port_valid(accel_io_argOuts_17_port_valid),
    .io_argOuts_17_port_bits(accel_io_argOuts_17_port_bits),
    .io_argOuts_17_echo(accel_io_argOuts_17_echo),
    .io_argOuts_18_port_ready(accel_io_argOuts_18_port_ready),
    .io_argOuts_18_port_valid(accel_io_argOuts_18_port_valid),
    .io_argOuts_18_port_bits(accel_io_argOuts_18_port_bits),
    .io_argOuts_18_echo(accel_io_argOuts_18_echo),
    .io_argOuts_19_port_ready(accel_io_argOuts_19_port_ready),
    .io_argOuts_19_port_valid(accel_io_argOuts_19_port_valid),
    .io_argOuts_19_port_bits(accel_io_argOuts_19_port_bits),
    .io_argOuts_19_echo(accel_io_argOuts_19_echo)
  );
  FringeZynq FringeZynq ( // @[KCU1500.scala 21:24:@57163.4]
    .clock(FringeZynq_clock),
    .reset(FringeZynq_reset),
    .io_S_AXI_AWADDR(FringeZynq_io_S_AXI_AWADDR),
    .io_S_AXI_AWPROT(FringeZynq_io_S_AXI_AWPROT),
    .io_S_AXI_AWVALID(FringeZynq_io_S_AXI_AWVALID),
    .io_S_AXI_AWREADY(FringeZynq_io_S_AXI_AWREADY),
    .io_S_AXI_ARADDR(FringeZynq_io_S_AXI_ARADDR),
    .io_S_AXI_ARPROT(FringeZynq_io_S_AXI_ARPROT),
    .io_S_AXI_ARVALID(FringeZynq_io_S_AXI_ARVALID),
    .io_S_AXI_ARREADY(FringeZynq_io_S_AXI_ARREADY),
    .io_S_AXI_WDATA(FringeZynq_io_S_AXI_WDATA),
    .io_S_AXI_WSTRB(FringeZynq_io_S_AXI_WSTRB),
    .io_S_AXI_WVALID(FringeZynq_io_S_AXI_WVALID),
    .io_S_AXI_WREADY(FringeZynq_io_S_AXI_WREADY),
    .io_S_AXI_RDATA(FringeZynq_io_S_AXI_RDATA),
    .io_S_AXI_RRESP(FringeZynq_io_S_AXI_RRESP),
    .io_S_AXI_RVALID(FringeZynq_io_S_AXI_RVALID),
    .io_S_AXI_RREADY(FringeZynq_io_S_AXI_RREADY),
    .io_S_AXI_BRESP(FringeZynq_io_S_AXI_BRESP),
    .io_S_AXI_BVALID(FringeZynq_io_S_AXI_BVALID),
    .io_S_AXI_BREADY(FringeZynq_io_S_AXI_BREADY),
    .io_M_AXI_0_AWLEN(FringeZynq_io_M_AXI_0_AWLEN),
    .io_M_AXI_0_ARLEN(FringeZynq_io_M_AXI_0_ARLEN),
    .io_enable(FringeZynq_io_enable),
    .io_done(FringeZynq_io_done),
    .io_reset(FringeZynq_io_reset),
    .io_argIns_0(FringeZynq_io_argIns_0),
    .io_argOuts_0_valid(FringeZynq_io_argOuts_0_valid),
    .io_argOuts_0_bits(FringeZynq_io_argOuts_0_bits),
    .io_argOuts_1_valid(FringeZynq_io_argOuts_1_valid),
    .io_argOuts_1_bits(FringeZynq_io_argOuts_1_bits),
    .io_argOuts_2_valid(FringeZynq_io_argOuts_2_valid),
    .io_argOuts_2_bits(FringeZynq_io_argOuts_2_bits),
    .io_argOuts_3_valid(FringeZynq_io_argOuts_3_valid),
    .io_argOuts_3_bits(FringeZynq_io_argOuts_3_bits),
    .io_argOuts_4_valid(FringeZynq_io_argOuts_4_valid),
    .io_argOuts_4_bits(FringeZynq_io_argOuts_4_bits),
    .io_argOuts_5_valid(FringeZynq_io_argOuts_5_valid),
    .io_argOuts_5_bits(FringeZynq_io_argOuts_5_bits),
    .io_argOuts_6_valid(FringeZynq_io_argOuts_6_valid),
    .io_argOuts_6_bits(FringeZynq_io_argOuts_6_bits),
    .io_argOuts_7_valid(FringeZynq_io_argOuts_7_valid),
    .io_argOuts_7_bits(FringeZynq_io_argOuts_7_bits),
    .io_argOuts_8_valid(FringeZynq_io_argOuts_8_valid),
    .io_argOuts_8_bits(FringeZynq_io_argOuts_8_bits),
    .io_argOuts_9_valid(FringeZynq_io_argOuts_9_valid),
    .io_argOuts_9_bits(FringeZynq_io_argOuts_9_bits),
    .io_argOuts_10_valid(FringeZynq_io_argOuts_10_valid),
    .io_argOuts_10_bits(FringeZynq_io_argOuts_10_bits),
    .io_argOuts_11_valid(FringeZynq_io_argOuts_11_valid),
    .io_argOuts_11_bits(FringeZynq_io_argOuts_11_bits),
    .io_argOuts_12_valid(FringeZynq_io_argOuts_12_valid),
    .io_argOuts_12_bits(FringeZynq_io_argOuts_12_bits),
    .io_argOuts_13_valid(FringeZynq_io_argOuts_13_valid),
    .io_argOuts_13_bits(FringeZynq_io_argOuts_13_bits),
    .io_argOuts_14_valid(FringeZynq_io_argOuts_14_valid),
    .io_argOuts_14_bits(FringeZynq_io_argOuts_14_bits),
    .io_argOuts_15_valid(FringeZynq_io_argOuts_15_valid),
    .io_argOuts_15_bits(FringeZynq_io_argOuts_15_bits),
    .io_argOuts_16_valid(FringeZynq_io_argOuts_16_valid),
    .io_argOuts_16_bits(FringeZynq_io_argOuts_16_bits),
    .io_argOuts_17_valid(FringeZynq_io_argOuts_17_valid),
    .io_argOuts_17_bits(FringeZynq_io_argOuts_17_bits),
    .io_argOuts_18_valid(FringeZynq_io_argOuts_18_valid),
    .io_argOuts_18_bits(FringeZynq_io_argOuts_18_bits),
    .io_argOuts_19_valid(FringeZynq_io_argOuts_19_valid),
    .io_argOuts_19_bits(FringeZynq_io_argOuts_19_bits),
    .io_heap_0_req_valid(FringeZynq_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(FringeZynq_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(FringeZynq_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(FringeZynq_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(FringeZynq_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(FringeZynq_io_heap_0_resp_bits_sizeAddr)
  );
  assign io_rdata = 1'h0;
  assign io_S_AXI_AWREADY = FringeZynq_io_S_AXI_AWREADY; // @[KCU1500.scala 24:21:@57181.4]
  assign io_S_AXI_ARREADY = FringeZynq_io_S_AXI_ARREADY; // @[KCU1500.scala 24:21:@57177.4]
  assign io_S_AXI_WREADY = FringeZynq_io_S_AXI_WREADY; // @[KCU1500.scala 24:21:@57173.4]
  assign io_S_AXI_RDATA = FringeZynq_io_S_AXI_RDATA; // @[KCU1500.scala 24:21:@57172.4]
  assign io_S_AXI_RRESP = FringeZynq_io_S_AXI_RRESP; // @[KCU1500.scala 24:21:@57171.4]
  assign io_S_AXI_RVALID = FringeZynq_io_S_AXI_RVALID; // @[KCU1500.scala 24:21:@57170.4]
  assign io_S_AXI_BRESP = FringeZynq_io_S_AXI_BRESP; // @[KCU1500.scala 24:21:@57168.4]
  assign io_S_AXI_BVALID = FringeZynq_io_S_AXI_BVALID; // @[KCU1500.scala 24:21:@57167.4]
  assign io_M_AXI_0_AWID = 4'h0; // @[KCU1500.scala 31:14:@57243.4]
  assign io_M_AXI_0_AWUSER = 4'h0; // @[KCU1500.scala 31:14:@57242.4]
  assign io_M_AXI_0_AWADDR = 32'h0; // @[KCU1500.scala 31:14:@57241.4]
  assign io_M_AXI_0_AWLEN = FringeZynq_io_M_AXI_0_AWLEN; // @[KCU1500.scala 31:14:@57240.4]
  assign io_M_AXI_0_AWSIZE = 3'h6; // @[KCU1500.scala 31:14:@57239.4]
  assign io_M_AXI_0_AWBURST = 2'h1; // @[KCU1500.scala 31:14:@57238.4]
  assign io_M_AXI_0_AWLOCK = 1'h0; // @[KCU1500.scala 31:14:@57237.4]
  assign io_M_AXI_0_AWCACHE = 4'h3; // @[KCU1500.scala 31:14:@57236.4]
  assign io_M_AXI_0_AWPROT = 3'h0; // @[KCU1500.scala 31:14:@57235.4]
  assign io_M_AXI_0_AWQOS = 4'h0; // @[KCU1500.scala 31:14:@57234.4]
  assign io_M_AXI_0_AWVALID = 1'h0; // @[KCU1500.scala 31:14:@57233.4]
  assign io_M_AXI_0_ARID = 4'h0; // @[KCU1500.scala 31:14:@57231.4]
  assign io_M_AXI_0_ARUSER = 4'h0; // @[KCU1500.scala 31:14:@57230.4]
  assign io_M_AXI_0_ARADDR = 32'h0; // @[KCU1500.scala 31:14:@57229.4]
  assign io_M_AXI_0_ARLEN = FringeZynq_io_M_AXI_0_ARLEN; // @[KCU1500.scala 31:14:@57228.4]
  assign io_M_AXI_0_ARSIZE = 3'h6; // @[KCU1500.scala 31:14:@57227.4]
  assign io_M_AXI_0_ARBURST = 2'h1; // @[KCU1500.scala 31:14:@57226.4]
  assign io_M_AXI_0_ARLOCK = 1'h0; // @[KCU1500.scala 31:14:@57225.4]
  assign io_M_AXI_0_ARCACHE = 4'h3; // @[KCU1500.scala 31:14:@57224.4]
  assign io_M_AXI_0_ARPROT = 3'h0; // @[KCU1500.scala 31:14:@57223.4]
  assign io_M_AXI_0_ARQOS = 4'h0; // @[KCU1500.scala 31:14:@57222.4]
  assign io_M_AXI_0_ARVALID = 1'h0; // @[KCU1500.scala 31:14:@57221.4]
  assign io_M_AXI_0_WDATA = 512'h0; // @[KCU1500.scala 31:14:@57219.4]
  assign io_M_AXI_0_WSTRB = 64'h0; // @[KCU1500.scala 31:14:@57218.4]
  assign io_M_AXI_0_WLAST = 1'h0; // @[KCU1500.scala 31:14:@57217.4]
  assign io_M_AXI_0_WVALID = 1'h0; // @[KCU1500.scala 31:14:@57216.4]
  assign io_M_AXI_0_RREADY = 1'h0; // @[KCU1500.scala 31:14:@57208.4]
  assign io_M_AXI_0_BREADY = 1'h0; // @[KCU1500.scala 31:14:@57203.4]
  assign io_AXIS_IN_TREADY = accel_io_axiStreamsIn_0_TREADY; // @[KCU1500.scala 27:16:@57192.4]
  assign io_AXIS_OUT_TVALID = accel_io_axiStreamsOut_0_TVALID; // @[KCU1500.scala 28:17:@57202.4]
  assign io_AXIS_OUT_TDATA = accel_io_axiStreamsOut_0_TDATA; // @[KCU1500.scala 28:17:@57200.4]
  assign io_AXIS_OUT_TSTRB = accel_io_axiStreamsOut_0_TSTRB; // @[KCU1500.scala 28:17:@57199.4]
  assign io_AXIS_OUT_TKEEP = accel_io_axiStreamsOut_0_TKEEP; // @[KCU1500.scala 28:17:@57198.4]
  assign io_AXIS_OUT_TLAST = accel_io_axiStreamsOut_0_TLAST; // @[KCU1500.scala 28:17:@57197.4]
  assign io_AXIS_OUT_TID = accel_io_axiStreamsOut_0_TID; // @[KCU1500.scala 28:17:@57196.4]
  assign io_AXIS_OUT_TDEST = accel_io_axiStreamsOut_0_TDEST; // @[KCU1500.scala 28:17:@57195.4]
  assign io_AXIS_OUT_TUSER = {{32'd0}, accel_io_axiStreamsOut_0_TUSER}; // @[KCU1500.scala 28:17:@57194.4]
  assign accel_clock = clock; // @[:@56932.4]
  assign accel_reset = FringeZynq_io_reset; // @[:@56933.4 KCU1500.scala 61:17:@57602.4]
  assign accel_io_enable = FringeZynq_io_enable; // @[KCU1500.scala 58:21:@57598.4]
  assign accel_io_reset = 1'h0;
  assign accel_io_memStreams_loads_0_cmd_ready = 1'h0; // @[KCU1500.scala 56:26:@57591.4]
  assign accel_io_memStreams_loads_0_data_valid = 1'h0; // @[KCU1500.scala 56:26:@57586.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_0 = 32'h0; // @[KCU1500.scala 56:26:@57570.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_1 = 32'h0; // @[KCU1500.scala 56:26:@57571.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_2 = 32'h0; // @[KCU1500.scala 56:26:@57572.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_3 = 32'h0; // @[KCU1500.scala 56:26:@57573.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_4 = 32'h0; // @[KCU1500.scala 56:26:@57574.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_5 = 32'h0; // @[KCU1500.scala 56:26:@57575.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_6 = 32'h0; // @[KCU1500.scala 56:26:@57576.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_7 = 32'h0; // @[KCU1500.scala 56:26:@57577.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_8 = 32'h0; // @[KCU1500.scala 56:26:@57578.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_9 = 32'h0; // @[KCU1500.scala 56:26:@57579.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_10 = 32'h0; // @[KCU1500.scala 56:26:@57580.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_11 = 32'h0; // @[KCU1500.scala 56:26:@57581.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_12 = 32'h0; // @[KCU1500.scala 56:26:@57582.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_13 = 32'h0; // @[KCU1500.scala 56:26:@57583.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_14 = 32'h0; // @[KCU1500.scala 56:26:@57584.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_15 = 32'h0; // @[KCU1500.scala 56:26:@57585.4]
  assign accel_io_memStreams_stores_0_cmd_ready = 1'h0; // @[KCU1500.scala 56:26:@57569.4]
  assign accel_io_memStreams_stores_0_data_ready = 1'h0; // @[KCU1500.scala 56:26:@57565.4]
  assign accel_io_memStreams_stores_0_wresp_valid = 1'h0; // @[KCU1500.scala 56:26:@57545.4]
  assign accel_io_memStreams_stores_0_wresp_bits = 1'h0; // @[KCU1500.scala 56:26:@57544.4]
  assign accel_io_memStreams_gathers_0_cmd_ready = 1'h0; // @[KCU1500.scala 56:26:@57543.4]
  assign accel_io_memStreams_gathers_0_data_valid = 1'h0; // @[KCU1500.scala 56:26:@57524.4]
  assign accel_io_memStreams_gathers_0_data_bits_0 = 32'h0; // @[KCU1500.scala 56:26:@57508.4]
  assign accel_io_memStreams_gathers_0_data_bits_1 = 32'h0; // @[KCU1500.scala 56:26:@57509.4]
  assign accel_io_memStreams_gathers_0_data_bits_2 = 32'h0; // @[KCU1500.scala 56:26:@57510.4]
  assign accel_io_memStreams_gathers_0_data_bits_3 = 32'h0; // @[KCU1500.scala 56:26:@57511.4]
  assign accel_io_memStreams_gathers_0_data_bits_4 = 32'h0; // @[KCU1500.scala 56:26:@57512.4]
  assign accel_io_memStreams_gathers_0_data_bits_5 = 32'h0; // @[KCU1500.scala 56:26:@57513.4]
  assign accel_io_memStreams_gathers_0_data_bits_6 = 32'h0; // @[KCU1500.scala 56:26:@57514.4]
  assign accel_io_memStreams_gathers_0_data_bits_7 = 32'h0; // @[KCU1500.scala 56:26:@57515.4]
  assign accel_io_memStreams_gathers_0_data_bits_8 = 32'h0; // @[KCU1500.scala 56:26:@57516.4]
  assign accel_io_memStreams_gathers_0_data_bits_9 = 32'h0; // @[KCU1500.scala 56:26:@57517.4]
  assign accel_io_memStreams_gathers_0_data_bits_10 = 32'h0; // @[KCU1500.scala 56:26:@57518.4]
  assign accel_io_memStreams_gathers_0_data_bits_11 = 32'h0; // @[KCU1500.scala 56:26:@57519.4]
  assign accel_io_memStreams_gathers_0_data_bits_12 = 32'h0; // @[KCU1500.scala 56:26:@57520.4]
  assign accel_io_memStreams_gathers_0_data_bits_13 = 32'h0; // @[KCU1500.scala 56:26:@57521.4]
  assign accel_io_memStreams_gathers_0_data_bits_14 = 32'h0; // @[KCU1500.scala 56:26:@57522.4]
  assign accel_io_memStreams_gathers_0_data_bits_15 = 32'h0; // @[KCU1500.scala 56:26:@57523.4]
  assign accel_io_memStreams_scatters_0_cmd_ready = 1'h0; // @[KCU1500.scala 56:26:@57507.4]
  assign accel_io_memStreams_scatters_0_wresp_valid = 1'h0; // @[KCU1500.scala 56:26:@57472.4]
  assign accel_io_memStreams_scatters_0_wresp_bits = 1'h0; // @[KCU1500.scala 56:26:@57471.4]
  assign accel_io_axiStreamsIn_0_TVALID = io_AXIS_IN_TVALID; // @[KCU1500.scala 27:16:@57193.4]
  assign accel_io_axiStreamsIn_0_TDATA = io_AXIS_IN_TDATA; // @[KCU1500.scala 27:16:@57191.4]
  assign accel_io_axiStreamsIn_0_TSTRB = io_AXIS_IN_TSTRB; // @[KCU1500.scala 27:16:@57190.4]
  assign accel_io_axiStreamsIn_0_TKEEP = io_AXIS_IN_TKEEP; // @[KCU1500.scala 27:16:@57189.4]
  assign accel_io_axiStreamsIn_0_TLAST = io_AXIS_IN_TLAST; // @[KCU1500.scala 27:16:@57188.4]
  assign accel_io_axiStreamsIn_0_TID = io_AXIS_IN_TID; // @[KCU1500.scala 27:16:@57187.4]
  assign accel_io_axiStreamsIn_0_TDEST = io_AXIS_IN_TDEST; // @[KCU1500.scala 27:16:@57186.4]
  assign accel_io_axiStreamsIn_0_TUSER = io_AXIS_IN_TUSER[31:0]; // @[KCU1500.scala 27:16:@57185.4]
  assign accel_io_axiStreamsOut_0_TREADY = io_AXIS_OUT_TREADY; // @[KCU1500.scala 28:17:@57201.4]
  assign accel_io_heap_0_resp_valid = FringeZynq_io_heap_0_resp_valid; // @[KCU1500.scala 57:20:@57594.4]
  assign accel_io_heap_0_resp_bits_allocDealloc = FringeZynq_io_heap_0_resp_bits_allocDealloc; // @[KCU1500.scala 57:20:@57593.4]
  assign accel_io_heap_0_resp_bits_sizeAddr = FringeZynq_io_heap_0_resp_bits_sizeAddr; // @[KCU1500.scala 57:20:@57592.4]
  assign accel_io_argIns_0 = FringeZynq_io_argIns_0; // @[KCU1500.scala 41:21:@57409.4]
  assign accel_io_argOuts_0_port_ready = 1'h0;
  assign accel_io_argOuts_0_echo = 64'h0; // @[KCU1500.scala 47:24:@57450.4]
  assign accel_io_argOuts_1_port_ready = 1'h0;
  assign accel_io_argOuts_1_echo = 64'h0; // @[KCU1500.scala 47:24:@57451.4]
  assign accel_io_argOuts_2_port_ready = 1'h0;
  assign accel_io_argOuts_2_echo = 64'h0; // @[KCU1500.scala 47:24:@57452.4]
  assign accel_io_argOuts_3_port_ready = 1'h0;
  assign accel_io_argOuts_3_echo = 64'h0; // @[KCU1500.scala 47:24:@57453.4]
  assign accel_io_argOuts_4_port_ready = 1'h0;
  assign accel_io_argOuts_4_echo = 64'h0; // @[KCU1500.scala 47:24:@57454.4]
  assign accel_io_argOuts_5_port_ready = 1'h0;
  assign accel_io_argOuts_5_echo = 64'h0; // @[KCU1500.scala 47:24:@57455.4]
  assign accel_io_argOuts_6_port_ready = 1'h0;
  assign accel_io_argOuts_6_echo = 64'h0; // @[KCU1500.scala 47:24:@57456.4]
  assign accel_io_argOuts_7_port_ready = 1'h0;
  assign accel_io_argOuts_7_echo = 64'h0; // @[KCU1500.scala 47:24:@57457.4]
  assign accel_io_argOuts_8_port_ready = 1'h0;
  assign accel_io_argOuts_8_echo = 64'h0; // @[KCU1500.scala 47:24:@57458.4]
  assign accel_io_argOuts_9_port_ready = 1'h0;
  assign accel_io_argOuts_9_echo = 64'h0; // @[KCU1500.scala 47:24:@57459.4]
  assign accel_io_argOuts_10_port_ready = 1'h0;
  assign accel_io_argOuts_10_echo = 64'h0; // @[KCU1500.scala 47:24:@57460.4]
  assign accel_io_argOuts_11_port_ready = 1'h0;
  assign accel_io_argOuts_11_echo = 64'h0; // @[KCU1500.scala 47:24:@57461.4]
  assign accel_io_argOuts_12_port_ready = 1'h0;
  assign accel_io_argOuts_12_echo = 64'h0; // @[KCU1500.scala 47:24:@57462.4]
  assign accel_io_argOuts_13_port_ready = 1'h0;
  assign accel_io_argOuts_13_echo = 64'h0; // @[KCU1500.scala 47:24:@57463.4]
  assign accel_io_argOuts_14_port_ready = 1'h0;
  assign accel_io_argOuts_14_echo = 64'h0; // @[KCU1500.scala 47:24:@57464.4]
  assign accel_io_argOuts_15_port_ready = 1'h0;
  assign accel_io_argOuts_15_echo = 64'h0; // @[KCU1500.scala 47:24:@57465.4]
  assign accel_io_argOuts_16_port_ready = 1'h0;
  assign accel_io_argOuts_16_echo = 64'h0; // @[KCU1500.scala 47:24:@57466.4]
  assign accel_io_argOuts_17_port_ready = 1'h0;
  assign accel_io_argOuts_17_echo = 64'h0; // @[KCU1500.scala 47:24:@57467.4]
  assign accel_io_argOuts_18_port_ready = 1'h0;
  assign accel_io_argOuts_18_echo = 64'h0; // @[KCU1500.scala 47:24:@57468.4]
  assign accel_io_argOuts_19_port_ready = 1'h0;
  assign accel_io_argOuts_19_echo = 64'h0; // @[KCU1500.scala 47:24:@57469.4]
  assign FringeZynq_clock = clock; // @[:@57164.4]
  assign FringeZynq_reset = reset; // @[:@57165.4 KCU1500.scala 60:18:@57601.4]
  assign FringeZynq_io_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[KCU1500.scala 24:21:@57184.4]
  assign FringeZynq_io_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[KCU1500.scala 24:21:@57183.4]
  assign FringeZynq_io_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[KCU1500.scala 24:21:@57182.4]
  assign FringeZynq_io_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[KCU1500.scala 24:21:@57180.4]
  assign FringeZynq_io_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[KCU1500.scala 24:21:@57179.4]
  assign FringeZynq_io_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[KCU1500.scala 24:21:@57178.4]
  assign FringeZynq_io_S_AXI_WDATA = io_S_AXI_WDATA; // @[KCU1500.scala 24:21:@57176.4]
  assign FringeZynq_io_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[KCU1500.scala 24:21:@57175.4]
  assign FringeZynq_io_S_AXI_WVALID = io_S_AXI_WVALID; // @[KCU1500.scala 24:21:@57174.4]
  assign FringeZynq_io_S_AXI_RREADY = io_S_AXI_RREADY; // @[KCU1500.scala 24:21:@57169.4]
  assign FringeZynq_io_S_AXI_BREADY = io_S_AXI_BREADY; // @[KCU1500.scala 24:21:@57166.4]
  assign FringeZynq_io_done = accel_io_done; // @[KCU1500.scala 59:20:@57599.4]
  assign FringeZynq_io_argOuts_0_valid = accel_io_argOuts_0_port_valid; // @[KCU1500.scala 44:26:@57411.4]
  assign FringeZynq_io_argOuts_0_bits = accel_io_argOuts_0_port_bits; // @[KCU1500.scala 43:25:@57410.4]
  assign FringeZynq_io_argOuts_1_valid = accel_io_argOuts_1_port_valid; // @[KCU1500.scala 44:26:@57413.4]
  assign FringeZynq_io_argOuts_1_bits = accel_io_argOuts_1_port_bits; // @[KCU1500.scala 43:25:@57412.4]
  assign FringeZynq_io_argOuts_2_valid = accel_io_argOuts_2_port_valid; // @[KCU1500.scala 44:26:@57415.4]
  assign FringeZynq_io_argOuts_2_bits = accel_io_argOuts_2_port_bits; // @[KCU1500.scala 43:25:@57414.4]
  assign FringeZynq_io_argOuts_3_valid = accel_io_argOuts_3_port_valid; // @[KCU1500.scala 44:26:@57417.4]
  assign FringeZynq_io_argOuts_3_bits = accel_io_argOuts_3_port_bits; // @[KCU1500.scala 43:25:@57416.4]
  assign FringeZynq_io_argOuts_4_valid = accel_io_argOuts_4_port_valid; // @[KCU1500.scala 44:26:@57419.4]
  assign FringeZynq_io_argOuts_4_bits = accel_io_argOuts_4_port_bits; // @[KCU1500.scala 43:25:@57418.4]
  assign FringeZynq_io_argOuts_5_valid = accel_io_argOuts_5_port_valid; // @[KCU1500.scala 44:26:@57421.4]
  assign FringeZynq_io_argOuts_5_bits = accel_io_argOuts_5_port_bits; // @[KCU1500.scala 43:25:@57420.4]
  assign FringeZynq_io_argOuts_6_valid = accel_io_argOuts_6_port_valid; // @[KCU1500.scala 44:26:@57423.4]
  assign FringeZynq_io_argOuts_6_bits = accel_io_argOuts_6_port_bits; // @[KCU1500.scala 43:25:@57422.4]
  assign FringeZynq_io_argOuts_7_valid = accel_io_argOuts_7_port_valid; // @[KCU1500.scala 44:26:@57425.4]
  assign FringeZynq_io_argOuts_7_bits = accel_io_argOuts_7_port_bits; // @[KCU1500.scala 43:25:@57424.4]
  assign FringeZynq_io_argOuts_8_valid = accel_io_argOuts_8_port_valid; // @[KCU1500.scala 44:26:@57427.4]
  assign FringeZynq_io_argOuts_8_bits = accel_io_argOuts_8_port_bits; // @[KCU1500.scala 43:25:@57426.4]
  assign FringeZynq_io_argOuts_9_valid = accel_io_argOuts_9_port_valid; // @[KCU1500.scala 44:26:@57429.4]
  assign FringeZynq_io_argOuts_9_bits = accel_io_argOuts_9_port_bits; // @[KCU1500.scala 43:25:@57428.4]
  assign FringeZynq_io_argOuts_10_valid = accel_io_argOuts_10_port_valid; // @[KCU1500.scala 44:26:@57431.4]
  assign FringeZynq_io_argOuts_10_bits = accel_io_argOuts_10_port_bits; // @[KCU1500.scala 43:25:@57430.4]
  assign FringeZynq_io_argOuts_11_valid = accel_io_argOuts_11_port_valid; // @[KCU1500.scala 44:26:@57433.4]
  assign FringeZynq_io_argOuts_11_bits = accel_io_argOuts_11_port_bits; // @[KCU1500.scala 43:25:@57432.4]
  assign FringeZynq_io_argOuts_12_valid = accel_io_argOuts_12_port_valid; // @[KCU1500.scala 44:26:@57435.4]
  assign FringeZynq_io_argOuts_12_bits = accel_io_argOuts_12_port_bits; // @[KCU1500.scala 43:25:@57434.4]
  assign FringeZynq_io_argOuts_13_valid = accel_io_argOuts_13_port_valid; // @[KCU1500.scala 44:26:@57437.4]
  assign FringeZynq_io_argOuts_13_bits = accel_io_argOuts_13_port_bits; // @[KCU1500.scala 43:25:@57436.4]
  assign FringeZynq_io_argOuts_14_valid = accel_io_argOuts_14_port_valid; // @[KCU1500.scala 44:26:@57439.4]
  assign FringeZynq_io_argOuts_14_bits = accel_io_argOuts_14_port_bits; // @[KCU1500.scala 43:25:@57438.4]
  assign FringeZynq_io_argOuts_15_valid = accel_io_argOuts_15_port_valid; // @[KCU1500.scala 44:26:@57441.4]
  assign FringeZynq_io_argOuts_15_bits = accel_io_argOuts_15_port_bits; // @[KCU1500.scala 43:25:@57440.4]
  assign FringeZynq_io_argOuts_16_valid = accel_io_argOuts_16_port_valid; // @[KCU1500.scala 44:26:@57443.4]
  assign FringeZynq_io_argOuts_16_bits = accel_io_argOuts_16_port_bits; // @[KCU1500.scala 43:25:@57442.4]
  assign FringeZynq_io_argOuts_17_valid = accel_io_argOuts_17_port_valid; // @[KCU1500.scala 44:26:@57445.4]
  assign FringeZynq_io_argOuts_17_bits = accel_io_argOuts_17_port_bits; // @[KCU1500.scala 43:25:@57444.4]
  assign FringeZynq_io_argOuts_18_valid = accel_io_argOuts_18_port_valid; // @[KCU1500.scala 44:26:@57447.4]
  assign FringeZynq_io_argOuts_18_bits = accel_io_argOuts_18_port_bits; // @[KCU1500.scala 43:25:@57446.4]
  assign FringeZynq_io_argOuts_19_valid = accel_io_argOuts_19_port_valid; // @[KCU1500.scala 44:26:@57449.4]
  assign FringeZynq_io_argOuts_19_bits = accel_io_argOuts_19_port_bits; // @[KCU1500.scala 43:25:@57448.4]
  assign FringeZynq_io_heap_0_req_valid = accel_io_heap_0_req_valid; // @[KCU1500.scala 57:20:@57597.4]
  assign FringeZynq_io_heap_0_req_bits_allocDealloc = accel_io_heap_0_req_bits_allocDealloc; // @[KCU1500.scala 57:20:@57596.4]
  assign FringeZynq_io_heap_0_req_bits_sizeAddr = accel_io_heap_0_req_bits_sizeAddr; // @[KCU1500.scala 57:20:@57595.4]
endmodule
module SRAMVerilogAWS
#(
    parameter WORDS = 1024,
    parameter AWIDTH = 10,
    parameter DWIDTH = 32)
(
    input clk,
    input [AWIDTH-1:0] raddr,
    input [AWIDTH-1:0] waddr,
    input raddrEn,
    input waddrEn,
    input wen,
    input [DWIDTH-1:0] wdata,
    input backpressure,
    output reg [DWIDTH-1:0] rdata
);

    reg [DWIDTH-1:0] mem [0:WORDS-1];

    always @(posedge clk) begin
      if (wen) mem[waddr] <= wdata;
      if (backpressure) rdata <= mem[raddr];
    end

endmodule
