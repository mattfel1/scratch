module FF( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  output [31:0] io_rPort_0_output_0, // @[:@6.4]
  input  [31:0] io_wPort_0_data_0, // @[:@6.4]
  input         io_wPort_0_reset, // @[:@6.4]
  input         io_wPort_0_en_0 // @[:@6.4]
);
  reg [31:0] ff; // @[MemPrimitives.scala 173:19:@21.4]
  reg [31:0] _RAND_0;
  wire [31:0] _T_68; // @[MemPrimitives.scala 177:32:@23.4]
  wire [31:0] _T_69; // @[MemPrimitives.scala 177:12:@24.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 177:32:@23.4]
  assign _T_69 = io_wPort_0_reset ? 32'h0 : _T_68; // @[MemPrimitives.scala 177:12:@24.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 178:34:@26.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 32'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 32'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SRFF( // @[:@28.2]
  input   clock, // @[:@29.4]
  input   reset, // @[:@30.4]
  input   io_input_set, // @[:@31.4]
  input   io_input_reset, // @[:@31.4]
  input   io_input_asyn_reset, // @[:@31.4]
  output  io_output // @[:@31.4]
);
  reg  _T_15; // @[SRFF.scala 20:21:@33.4]
  reg [31:0] _RAND_0;
  wire  _T_19; // @[SRFF.scala 21:74:@34.4]
  wire  _T_20; // @[SRFF.scala 21:48:@35.4]
  wire  _T_21; // @[SRFF.scala 21:14:@36.4]
  assign _T_19 = io_input_reset ? 1'h0 : _T_15; // @[SRFF.scala 21:74:@34.4]
  assign _T_20 = io_input_set ? 1'h1 : _T_19; // @[SRFF.scala 21:48:@35.4]
  assign _T_21 = io_input_asyn_reset ? 1'h0 : _T_20; // @[SRFF.scala 21:14:@36.4]
  assign io_output = io_input_asyn_reset ? 1'h0 : _T_15; // @[SRFF.scala 22:15:@39.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_15 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_15 <= 1'h0;
    end else begin
      if (io_input_asyn_reset) begin
        _T_15 <= 1'h0;
      end else begin
        if (io_input_set) begin
          _T_15 <= 1'h1;
        end else begin
          if (io_input_reset) begin
            _T_15 <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module SingleCounter( // @[:@41.2]
  input   clock, // @[:@42.4]
  input   reset, // @[:@43.4]
  input   io_input_reset, // @[:@44.4]
  output  io_output_done // @[:@44.4]
);
  wire  bases_0_clock; // @[Counter.scala 253:53:@57.4]
  wire  bases_0_reset; // @[Counter.scala 253:53:@57.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 253:53:@57.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 253:53:@57.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 253:53:@57.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 253:53:@57.4]
  wire  SRFF_clock; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_reset; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_input_set; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_output; // @[Counter.scala 255:22:@73.4]
  wire [31:0] _T_48; // @[Counter.scala 279:52:@101.4]
  wire [32:0] _T_50; // @[Counter.scala 283:33:@102.4]
  wire [31:0] _T_51; // @[Counter.scala 283:33:@103.4]
  wire [31:0] _T_52; // @[Counter.scala 283:33:@104.4]
  wire  _T_57; // @[Counter.scala 285:18:@106.4]
  wire [31:0] _T_68; // @[Counter.scala 291:115:@114.4]
  wire [31:0] _T_71; // @[Counter.scala 291:152:@117.4]
  wire [31:0] _T_72; // @[Counter.scala 291:74:@118.4]
  FF bases_0 ( // @[Counter.scala 253:53:@57.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 255:22:@73.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 279:52:@101.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@102.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@103.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 283:33:@104.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh2); // @[Counter.scala 285:18:@106.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 291:115:@114.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 291:152:@117.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 291:74:@118.4]
  assign io_output_done = $signed(_T_52) >= $signed(32'sh2); // @[Counter.scala 325:20:@127.4]
  assign bases_0_clock = clock; // @[:@58.4]
  assign bases_0_reset = reset; // @[:@59.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 291:31:@120.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 273:27:@99.4]
  assign bases_0_io_wPort_0_en_0 = 1'h1; // @[Counter.scala 276:29:@100.4]
  assign SRFF_clock = clock; // @[:@74.4]
  assign SRFF_reset = reset; // @[:@75.4]
  assign SRFF_io_input_set = io_input_reset == 1'h0; // @[Counter.scala 256:23:@78.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 257:25:@80.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 258:30:@81.4]
endmodule
module RetimeWrapper( // @[:@144.2]
  input   clock, // @[:@145.4]
  input   reset, // @[:@146.4]
  input   io_flow, // @[:@147.4]
  input   io_in, // @[:@147.4]
  output  io_out // @[:@147.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@149.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@149.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@162.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@161.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@160.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@159.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@158.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@156.4]
endmodule
module RootController_sm( // @[:@351.2]
  input   clock, // @[:@352.4]
  input   reset, // @[:@353.4]
  input   io_enable, // @[:@354.4]
  output  io_done, // @[:@354.4]
  input   io_rst, // @[:@354.4]
  input   io_ctrDone, // @[:@354.4]
  output  io_ctrInc, // @[:@354.4]
  input   io_doneIn_0, // @[:@354.4]
  input   io_doneIn_1, // @[:@354.4]
  output  io_enableOut_0, // @[:@354.4]
  output  io_enableOut_1, // @[:@354.4]
  output  io_childAck_0, // @[:@354.4]
  output  io_childAck_1 // @[:@354.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@357.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@357.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@357.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@357.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@357.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@357.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@360.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@360.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@360.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@360.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@360.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@360.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@363.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@363.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@363.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@363.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@363.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@363.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@366.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@366.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@366.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@366.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@366.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@366.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@395.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@395.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@395.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@395.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@395.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@395.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@398.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@398.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@398.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@398.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@398.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@398.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@427.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@427.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@427.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@427.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@427.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@523.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@523.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@523.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@523.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@523.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@540.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@540.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@540.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@540.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@540.4]
  wire  allDone; // @[Controllers.scala 80:47:@369.4]
  wire  _T_77; // @[Controllers.scala 81:26:@370.4]
  wire  finished; // @[Controllers.scala 81:37:@371.4]
  wire  synchronize; // @[package.scala 96:25:@432.4 package.scala 96:25:@433.4]
  wire  _T_144; // @[Controllers.scala 128:33:@441.4]
  wire  _T_146; // @[Controllers.scala 128:54:@442.4]
  wire  _T_147; // @[Controllers.scala 128:52:@443.4]
  wire  _T_148; // @[Controllers.scala 128:66:@444.4]
  wire  _T_150; // @[Controllers.scala 128:98:@446.4]
  wire  _T_151; // @[Controllers.scala 128:96:@447.4]
  wire  _T_153; // @[Controllers.scala 128:123:@448.4]
  wire  _T_155; // @[Controllers.scala 129:48:@451.4]
  wire  _T_160; // @[Controllers.scala 130:52:@456.4]
  wire  _T_161; // @[Controllers.scala 130:50:@457.4]
  wire  _T_169; // @[Controllers.scala 130:129:@463.4]
  wire  _T_172; // @[Controllers.scala 131:45:@466.4]
  wire  _T_175; // @[Controllers.scala 135:80:@470.4]
  wire  _T_176; // @[Controllers.scala 135:78:@471.4]
  wire  _T_178; // @[Controllers.scala 135:105:@472.4]
  wire  _T_179; // @[Controllers.scala 135:103:@473.4]
  wire  _T_180; // @[Controllers.scala 135:119:@474.4]
  wire  _T_182; // @[Controllers.scala 135:51:@476.4]
  wire  _T_205; // @[Controllers.scala 213:68:@501.4]
  wire  _T_207; // @[Controllers.scala 213:90:@503.4]
  wire  _T_209; // @[Controllers.scala 213:132:@505.4]
  wire  _T_210; // @[Controllers.scala 213:130:@506.4]
  wire  _T_211; // @[Controllers.scala 213:156:@507.4]
  wire  _T_213; // @[Controllers.scala 213:68:@510.4]
  wire  _T_215; // @[Controllers.scala 213:90:@512.4]
  wire  _T_222; // @[package.scala 100:49:@518.4]
  reg  _T_225; // @[package.scala 48:56:@519.4]
  reg [31:0] _RAND_0;
  reg  _T_239; // @[package.scala 48:56:@537.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@357.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@360.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@363.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@366.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@395.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@398.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@427.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@523.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@540.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  assign allDone = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@369.4]
  assign _T_77 = allDone | io_done; // @[Controllers.scala 81:26:@370.4]
  assign finished = _T_77 | done_1_io_input_set; // @[Controllers.scala 81:37:@371.4]
  assign synchronize = RetimeWrapper_io_out; // @[package.scala 96:25:@432.4 package.scala 96:25:@433.4]
  assign _T_144 = done_0_io_output == 1'h0; // @[Controllers.scala 128:33:@441.4]
  assign _T_146 = io_ctrDone == 1'h0; // @[Controllers.scala 128:54:@442.4]
  assign _T_147 = _T_144 & _T_146; // @[Controllers.scala 128:52:@443.4]
  assign _T_148 = _T_147 & io_enable; // @[Controllers.scala 128:66:@444.4]
  assign _T_150 = ~ iterDone_0_io_output; // @[Controllers.scala 128:98:@446.4]
  assign _T_151 = _T_148 & _T_150; // @[Controllers.scala 128:96:@447.4]
  assign _T_153 = io_doneIn_0 == 1'h0; // @[Controllers.scala 128:123:@448.4]
  assign _T_155 = io_doneIn_0 | io_rst; // @[Controllers.scala 129:48:@451.4]
  assign _T_160 = synchronize == 1'h0; // @[Controllers.scala 130:52:@456.4]
  assign _T_161 = io_doneIn_0 & _T_160; // @[Controllers.scala 130:50:@457.4]
  assign _T_169 = finished == 1'h0; // @[Controllers.scala 130:129:@463.4]
  assign _T_172 = io_rst == 1'h0; // @[Controllers.scala 131:45:@466.4]
  assign _T_175 = ~ iterDone_1_io_output; // @[Controllers.scala 135:80:@470.4]
  assign _T_176 = iterDone_0_io_output & _T_175; // @[Controllers.scala 135:78:@471.4]
  assign _T_178 = io_doneIn_1 == 1'h0; // @[Controllers.scala 135:105:@472.4]
  assign _T_179 = _T_176 & _T_178; // @[Controllers.scala 135:103:@473.4]
  assign _T_180 = _T_179 & io_enable; // @[Controllers.scala 135:119:@474.4]
  assign _T_182 = io_doneIn_0 | _T_180; // @[Controllers.scala 135:51:@476.4]
  assign _T_205 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@501.4]
  assign _T_207 = _T_205 & _T_150; // @[Controllers.scala 213:90:@503.4]
  assign _T_209 = ~ allDone; // @[Controllers.scala 213:132:@505.4]
  assign _T_210 = _T_207 & _T_209; // @[Controllers.scala 213:130:@506.4]
  assign _T_211 = ~ io_ctrDone; // @[Controllers.scala 213:156:@507.4]
  assign _T_213 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@510.4]
  assign _T_215 = _T_213 & _T_175; // @[Controllers.scala 213:90:@512.4]
  assign _T_222 = allDone == 1'h0; // @[package.scala 100:49:@518.4]
  assign io_done = RetimeWrapper_2_io_out; // @[Controllers.scala 245:13:@547.4]
  assign io_ctrInc = io_doneIn_1; // @[Controllers.scala 122:17:@426.4]
  assign io_enableOut_0 = _T_210 & _T_211; // @[Controllers.scala 213:55:@509.4]
  assign io_enableOut_1 = _T_215 & _T_209; // @[Controllers.scala 213:55:@517.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@498.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@500.4]
  assign active_0_clock = clock; // @[:@358.4]
  assign active_0_reset = reset; // @[:@359.4]
  assign active_0_io_input_set = _T_151 & _T_153; // @[Controllers.scala 128:30:@450.4]
  assign active_0_io_input_reset = _T_155 | allDone; // @[Controllers.scala 129:32:@455.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@372.4]
  assign active_1_clock = clock; // @[:@361.4]
  assign active_1_reset = reset; // @[:@362.4]
  assign active_1_io_input_set = _T_182 & _T_160; // @[Controllers.scala 135:32:@479.4]
  assign active_1_io_input_reset = io_doneIn_1 | io_rst; // @[Controllers.scala 136:34:@483.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@373.4]
  assign done_0_clock = clock; // @[:@364.4]
  assign done_0_reset = reset; // @[:@365.4]
  assign done_0_io_input_set = io_ctrDone & _T_172; // @[Controllers.scala 131:28:@469.4]
  assign done_0_io_input_reset = io_rst | allDone; // @[Controllers.scala 86:33:@384.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@374.4]
  assign done_1_clock = clock; // @[:@367.4]
  assign done_1_reset = reset; // @[:@368.4]
  assign done_1_io_input_set = io_ctrDone & _T_172; // @[Controllers.scala 138:30:@496.4]
  assign done_1_io_input_reset = io_rst | allDone; // @[Controllers.scala 86:33:@393.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@375.4]
  assign iterDone_0_clock = clock; // @[:@396.4]
  assign iterDone_0_reset = reset; // @[:@397.4]
  assign iterDone_0_io_input_set = _T_161 & _T_169; // @[Controllers.scala 130:32:@465.4]
  assign iterDone_0_io_input_reset = synchronize | io_rst; // @[Controllers.scala 92:37:@411.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@401.4]
  assign iterDone_1_clock = clock; // @[:@399.4]
  assign iterDone_1_reset = reset; // @[:@400.4]
  assign iterDone_1_io_input_set = io_doneIn_1 & _T_160; // @[Controllers.scala 137:34:@492.4]
  assign iterDone_1_io_input_reset = synchronize | io_rst; // @[Controllers.scala 92:37:@420.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@402.4]
  assign RetimeWrapper_clock = clock; // @[:@428.4]
  assign RetimeWrapper_reset = reset; // @[:@429.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@431.4]
  assign RetimeWrapper_io_in = io_doneIn_1; // @[package.scala 94:16:@430.4]
  assign RetimeWrapper_1_clock = clock; // @[:@524.4]
  assign RetimeWrapper_1_reset = reset; // @[:@525.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@527.4]
  assign RetimeWrapper_1_io_in = allDone & _T_225; // @[package.scala 94:16:@526.4]
  assign RetimeWrapper_2_clock = clock; // @[:@541.4]
  assign RetimeWrapper_2_reset = reset; // @[:@542.4]
  assign RetimeWrapper_2_io_flow = io_enable; // @[package.scala 95:18:@544.4]
  assign RetimeWrapper_2_io_in = allDone & _T_239; // @[package.scala 94:16:@543.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_225 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_239 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_225 <= 1'h0;
    end else begin
      _T_225 <= _T_222;
    end
    if (reset) begin
      _T_239 <= 1'h0;
    end else begin
      _T_239 <= _T_222;
    end
  end
endmodule
module InstrumentationCounter( // @[:@597.2]
  input         clock, // @[:@598.4]
  input         reset, // @[:@599.4]
  input         io_enable, // @[:@600.4]
  output [63:0] io_count // @[:@600.4]
);
  reg [63:0] ff; // @[Counter.scala 214:19:@602.4]
  reg [63:0] _RAND_0;
  wire [64:0] _T_12; // @[Counter.scala 215:27:@603.4]
  wire [63:0] _T_13; // @[Counter.scala 215:27:@604.4]
  wire [63:0] _T_14; // @[Counter.scala 215:12:@605.4]
  assign _T_12 = ff + 64'h1; // @[Counter.scala 215:27:@603.4]
  assign _T_13 = ff + 64'h1; // @[Counter.scala 215:27:@604.4]
  assign _T_14 = io_enable ? _T_13 : ff; // @[Counter.scala 215:12:@605.4]
  assign io_count = ff; // @[Counter.scala 216:12:@607.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  ff = _RAND_0[63:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 64'h0;
    end else begin
      if (io_enable) begin
        ff <= _T_13;
      end
    end
  end
endmodule
module SRAM( // @[:@637.2]
  input         clock, // @[:@638.4]
  input         reset, // @[:@639.4]
  input  [2:0]  io_raddr, // @[:@640.4]
  input         io_wen, // @[:@640.4]
  input  [2:0]  io_waddr, // @[:@640.4]
  input  [63:0] io_wdata, // @[:@640.4]
  output [63:0] io_rdata, // @[:@640.4]
  input         io_backpressure // @[:@640.4]
);
  wire [63:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 124:30:@642.4]
  wire [63:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 124:30:@642.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 124:30:@642.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 124:30:@642.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 124:30:@642.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 124:30:@642.4]
  wire [2:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 124:30:@642.4]
  wire [2:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 124:30:@642.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 124:30:@642.4]
  wire  _T_19; // @[SRAM.scala 137:49:@660.4]
  wire  _T_20; // @[SRAM.scala 137:37:@661.4]
  reg  _T_23; // @[SRAM.scala 137:29:@662.4]
  reg [31:0] _RAND_0;
  reg [63:0] _T_26; // @[SRAM.scala 138:29:@664.4]
  reg [63:0] _RAND_1;
  SRAMVerilogAWS #(.DWIDTH(64), .WORDS(8), .AWIDTH(3)) SRAMVerilogAWS ( // @[SRAM.scala 124:30:@642.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_19 = io_raddr == io_waddr; // @[SRAM.scala 137:49:@660.4]
  assign _T_20 = io_wen & _T_19; // @[SRAM.scala 137:37:@661.4]
  assign io_rdata = _T_23 ? _T_26 : SRAMVerilogAWS_rdata; // @[SRAM.scala 139:16:@669.4]
  assign SRAMVerilogAWS_wdata = io_wdata; // @[SRAM.scala 130:20:@656.4]
  assign SRAMVerilogAWS_backpressure = io_backpressure; // @[SRAM.scala 131:27:@657.4]
  assign SRAMVerilogAWS_wen = io_wen; // @[SRAM.scala 128:18:@654.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 133:22:@659.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 132:22:@658.4]
  assign SRAMVerilogAWS_waddr = io_waddr; // @[SRAM.scala 129:20:@655.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 127:20:@653.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 126:18:@652.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_23 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {2{`RANDOM}};
  _T_26 = _RAND_1[63:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_23 <= 1'h0;
    end else begin
      _T_23 <= _T_20;
    end
    if (reset) begin
      _T_26 <= 64'h0;
    end else begin
      _T_26 <= io_wdata;
    end
  end
endmodule
module RetimeWrapper_5( // @[:@683.2]
  input        clock, // @[:@684.4]
  input        reset, // @[:@685.4]
  input        io_flow, // @[:@686.4]
  input  [3:0] io_in, // @[:@686.4]
  output [3:0] io_out // @[:@686.4]
);
  wire [3:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@688.4]
  wire [3:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@688.4]
  wire [3:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@688.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@688.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@688.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@688.4]
  RetimeShiftRegister #(.WIDTH(4), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@688.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@701.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@700.4]
  assign sr_init = 4'h0; // @[RetimeShiftRegister.scala 19:16:@699.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@698.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@697.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@695.4]
endmodule
module Mem1D( // @[:@703.2]
  input         clock, // @[:@704.4]
  input         reset, // @[:@705.4]
  input  [3:0]  io_r_ofs_0, // @[:@706.4]
  input         io_r_backpressure, // @[:@706.4]
  input  [3:0]  io_w_ofs_0, // @[:@706.4]
  input  [63:0] io_w_data_0, // @[:@706.4]
  input         io_w_en_0, // @[:@706.4]
  output [63:0] io_output // @[:@706.4]
);
  wire  SRAM_clock; // @[MemPrimitives.scala 567:21:@710.4]
  wire  SRAM_reset; // @[MemPrimitives.scala 567:21:@710.4]
  wire [2:0] SRAM_io_raddr; // @[MemPrimitives.scala 567:21:@710.4]
  wire  SRAM_io_wen; // @[MemPrimitives.scala 567:21:@710.4]
  wire [2:0] SRAM_io_waddr; // @[MemPrimitives.scala 567:21:@710.4]
  wire [63:0] SRAM_io_wdata; // @[MemPrimitives.scala 567:21:@710.4]
  wire [63:0] SRAM_io_rdata; // @[MemPrimitives.scala 567:21:@710.4]
  wire  SRAM_io_backpressure; // @[MemPrimitives.scala 567:21:@710.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@713.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@713.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@713.4]
  wire [3:0] RetimeWrapper_io_in; // @[package.scala 93:22:@713.4]
  wire [3:0] RetimeWrapper_io_out; // @[package.scala 93:22:@713.4]
  wire  wInBound; // @[MemPrimitives.scala 554:32:@708.4]
  wire [3:0] _T_126; // @[package.scala 96:25:@718.4 package.scala 96:25:@719.4]
  SRAM SRAM ( // @[MemPrimitives.scala 567:21:@710.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata(SRAM_io_wdata),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  RetimeWrapper_5 RetimeWrapper ( // @[package.scala 93:22:@713.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign wInBound = io_w_ofs_0 <= 4'h8; // @[MemPrimitives.scala 554:32:@708.4]
  assign _T_126 = RetimeWrapper_io_out; // @[package.scala 96:25:@718.4 package.scala 96:25:@719.4]
  assign io_output = SRAM_io_rdata; // @[MemPrimitives.scala 574:17:@726.4]
  assign SRAM_clock = clock; // @[:@711.4]
  assign SRAM_reset = reset; // @[:@712.4]
  assign SRAM_io_raddr = _T_126[2:0]; // @[MemPrimitives.scala 568:37:@720.4]
  assign SRAM_io_wen = io_w_en_0 & wInBound; // @[MemPrimitives.scala 571:22:@723.4]
  assign SRAM_io_waddr = io_w_ofs_0[2:0]; // @[MemPrimitives.scala 570:22:@721.4]
  assign SRAM_io_wdata = io_w_data_0; // @[MemPrimitives.scala 572:22:@724.4]
  assign SRAM_io_backpressure = io_r_backpressure; // @[MemPrimitives.scala 573:30:@725.4]
  assign RetimeWrapper_clock = clock; // @[:@714.4]
  assign RetimeWrapper_reset = reset; // @[:@715.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@717.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@716.4]
endmodule
module StickySelects( // @[:@728.2]
  input   io_ins_0, // @[:@731.4]
  output  io_outs_0 // @[:@731.4]
);
  assign io_outs_0 = io_ins_0; // @[StickySelects.scala 12:26:@733.4]
endmodule
module RetimeWrapper_6( // @[:@747.2]
  input   clock, // @[:@748.4]
  input   reset, // @[:@749.4]
  input   io_flow, // @[:@750.4]
  input   io_in, // @[:@750.4]
  output  io_out // @[:@750.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@752.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@752.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@752.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@752.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@752.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@752.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@752.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@765.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@764.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@763.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@762.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@761.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@759.4]
endmodule
module x84_a_0( // @[:@767.2]
  input         clock, // @[:@768.4]
  input         reset, // @[:@769.4]
  input  [3:0]  io_rPort_0_ofs_0, // @[:@770.4]
  input         io_rPort_0_en_0, // @[:@770.4]
  input         io_rPort_0_backpressure, // @[:@770.4]
  output [63:0] io_rPort_0_output_0, // @[:@770.4]
  input  [3:0]  io_wPort_0_ofs_0, // @[:@770.4]
  input  [63:0] io_wPort_0_data_0, // @[:@770.4]
  input         io_wPort_0_en_0 // @[:@770.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@785.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@785.4]
  wire [3:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@785.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@785.4]
  wire [3:0] Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@785.4]
  wire [63:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@785.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@785.4]
  wire [63:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@785.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 121:29:@811.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 121:29:@811.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@825.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@825.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@825.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@825.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@825.4]
  wire [68:0] _T_70; // @[Cat.scala 30:58:@803.4]
  wire  _T_76; // @[MemPrimitives.scala 123:41:@815.4]
  wire [5:0] _T_78; // @[Cat.scala 30:58:@817.4]
  Mem1D Mem1D ( // @[MemPrimitives.scala 64:21:@785.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  StickySelects StickySelects ( // @[MemPrimitives.scala 121:29:@811.4]
    .io_ins_0(StickySelects_io_ins_0),
    .io_outs_0(StickySelects_io_outs_0)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@825.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_70 = {io_wPort_0_en_0,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@803.4]
  assign _T_76 = StickySelects_io_outs_0; // @[MemPrimitives.scala 123:41:@815.4]
  assign _T_78 = {_T_76,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@817.4]
  assign io_rPort_0_output_0 = Mem1D_io_output; // @[MemPrimitives.scala 148:13:@832.4]
  assign Mem1D_clock = clock; // @[:@786.4]
  assign Mem1D_reset = reset; // @[:@787.4]
  assign Mem1D_io_r_ofs_0 = _T_78[3:0]; // @[MemPrimitives.scala 127:28:@821.4]
  assign Mem1D_io_r_backpressure = _T_78[4]; // @[MemPrimitives.scala 128:32:@822.4]
  assign Mem1D_io_w_ofs_0 = _T_70[3:0]; // @[MemPrimitives.scala 94:28:@807.4]
  assign Mem1D_io_w_data_0 = _T_70[67:4]; // @[MemPrimitives.scala 95:29:@808.4]
  assign Mem1D_io_w_en_0 = _T_70[68]; // @[MemPrimitives.scala 96:27:@809.4]
  assign StickySelects_io_ins_0 = io_rPort_0_en_0; // @[MemPrimitives.scala 122:60:@814.4]
  assign RetimeWrapper_clock = clock; // @[:@826.4]
  assign RetimeWrapper_reset = reset; // @[:@827.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@829.4]
  assign RetimeWrapper_io_in = io_rPort_0_en_0; // @[package.scala 94:16:@828.4]
endmodule
module SingleCounter_1( // @[:@872.2]
  input         clock, // @[:@873.4]
  input         reset, // @[:@874.4]
  input         io_input_reset, // @[:@875.4]
  input         io_input_enable, // @[:@875.4]
  output [31:0] io_output_count_0, // @[:@875.4]
  output        io_output_oobs_0, // @[:@875.4]
  output        io_output_done // @[:@875.4]
);
  wire  bases_0_clock; // @[Counter.scala 253:53:@888.4]
  wire  bases_0_reset; // @[Counter.scala 253:53:@888.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 253:53:@888.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 253:53:@888.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 253:53:@888.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 253:53:@888.4]
  wire  SRFF_clock; // @[Counter.scala 255:22:@904.4]
  wire  SRFF_reset; // @[Counter.scala 255:22:@904.4]
  wire  SRFF_io_input_set; // @[Counter.scala 255:22:@904.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 255:22:@904.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 255:22:@904.4]
  wire  SRFF_io_output; // @[Counter.scala 255:22:@904.4]
  wire  _T_36; // @[Counter.scala 256:45:@907.4]
  wire [31:0] _T_48; // @[Counter.scala 279:52:@932.4]
  wire [32:0] _T_50; // @[Counter.scala 283:33:@933.4]
  wire [31:0] _T_51; // @[Counter.scala 283:33:@934.4]
  wire [31:0] _T_52; // @[Counter.scala 283:33:@935.4]
  wire  _T_57; // @[Counter.scala 285:18:@937.4]
  wire [31:0] _T_68; // @[Counter.scala 291:115:@945.4]
  wire [31:0] _T_71; // @[Counter.scala 291:152:@948.4]
  wire [31:0] _T_72; // @[Counter.scala 291:74:@949.4]
  wire  _T_75; // @[Counter.scala 314:102:@953.4]
  wire  _T_77; // @[Counter.scala 314:130:@954.4]
  FF bases_0 ( // @[Counter.scala 253:53:@888.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 255:22:@904.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 256:45:@907.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 279:52:@932.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh4); // @[Counter.scala 283:33:@933.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh4); // @[Counter.scala 283:33:@934.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 283:33:@935.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh20); // @[Counter.scala 285:18:@937.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 291:115:@945.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 291:152:@948.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 291:74:@949.4]
  assign _T_75 = $signed(_T_48) < $signed(32'sh0); // @[Counter.scala 314:102:@953.4]
  assign _T_77 = $signed(_T_48) >= $signed(32'sh20); // @[Counter.scala 314:130:@954.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 296:28:@952.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 314:60:@956.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 325:20:@958.4]
  assign bases_0_clock = clock; // @[:@889.4]
  assign bases_0_reset = reset; // @[:@890.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 291:31:@951.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 273:27:@930.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 276:29:@931.4]
  assign SRFF_clock = clock; // @[:@905.4]
  assign SRFF_reset = reset; // @[:@906.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 256:23:@909.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 257:25:@911.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 258:30:@912.4]
endmodule
module x86_ctrchain( // @[:@963.2]
  input         clock, // @[:@964.4]
  input         reset, // @[:@965.4]
  input         io_input_reset, // @[:@966.4]
  input         io_input_enable, // @[:@966.4]
  output [31:0] io_output_counts_0, // @[:@966.4]
  output        io_output_oobs_0, // @[:@966.4]
  output        io_output_done // @[:@966.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 505:46:@968.4]
  wire  ctrs_0_reset; // @[Counter.scala 505:46:@968.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 505:46:@968.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 505:46:@968.4]
  wire [31:0] ctrs_0_io_output_count_0; // @[Counter.scala 505:46:@968.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 505:46:@968.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 505:46:@968.4]
  reg  wasDone; // @[Counter.scala 534:24:@977.4]
  reg [31:0] _RAND_0;
  wire  _T_45; // @[Counter.scala 538:69:@983.4]
  wire  _T_47; // @[Counter.scala 538:80:@984.4]
  reg  doneLatch; // @[Counter.scala 542:26:@989.4]
  reg [31:0] _RAND_1;
  wire  _T_54; // @[Counter.scala 543:48:@990.4]
  wire  _T_55; // @[Counter.scala 543:19:@991.4]
  SingleCounter_1 ctrs_0 ( // @[Counter.scala 505:46:@968.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done)
  );
  assign _T_45 = io_input_enable & ctrs_0_io_output_done; // @[Counter.scala 538:69:@983.4]
  assign _T_47 = wasDone == 1'h0; // @[Counter.scala 538:80:@984.4]
  assign _T_54 = ctrs_0_io_output_done ? 1'h1 : doneLatch; // @[Counter.scala 543:48:@990.4]
  assign _T_55 = io_input_reset ? 1'h0 : _T_54; // @[Counter.scala 543:19:@991.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 549:32:@993.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 550:30:@995.4]
  assign io_output_done = _T_45 & _T_47; // @[Counter.scala 538:18:@986.4]
  assign ctrs_0_clock = clock; // @[:@969.4]
  assign ctrs_0_reset = reset; // @[:@970.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 512:24:@974.4]
  assign ctrs_0_io_input_enable = io_input_enable; // @[Counter.scala 516:33:@975.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= ctrs_0_io_output_done;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (ctrs_0_io_output_done) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module x102_inr_Foreach_sm( // @[:@1183.2]
  input   clock, // @[:@1184.4]
  input   reset, // @[:@1185.4]
  input   io_enable, // @[:@1186.4]
  output  io_done, // @[:@1186.4]
  output  io_doneLatch, // @[:@1186.4]
  input   io_ctrDone, // @[:@1186.4]
  output  io_datapathEn, // @[:@1186.4]
  output  io_ctrInc, // @[:@1186.4]
  output  io_ctrRst, // @[:@1186.4]
  input   io_parentAck, // @[:@1186.4]
  input   io_backpressure, // @[:@1186.4]
  input   io_break // @[:@1186.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@1188.4]
  wire  active_reset; // @[Controllers.scala 261:22:@1188.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@1188.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@1188.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@1188.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@1188.4]
  wire  done_clock; // @[Controllers.scala 262:20:@1191.4]
  wire  done_reset; // @[Controllers.scala 262:20:@1191.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@1191.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@1191.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@1191.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@1191.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@1225.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@1225.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@1225.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@1225.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@1225.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@1247.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@1247.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@1247.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@1247.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@1247.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@1259.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@1259.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@1259.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@1259.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@1259.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@1267.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@1267.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@1267.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@1267.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@1267.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@1283.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@1283.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@1283.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@1283.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@1283.4]
  wire  _T_80; // @[Controllers.scala 264:48:@1196.4]
  wire  _T_81; // @[Controllers.scala 264:46:@1197.4]
  wire  _T_82; // @[Controllers.scala 264:62:@1198.4]
  wire  _T_83; // @[Controllers.scala 264:60:@1199.4]
  wire  _T_100; // @[package.scala 100:49:@1216.4]
  reg  _T_103; // @[package.scala 48:56:@1217.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@1230.4 package.scala 96:25:@1231.4]
  wire  _T_110; // @[package.scala 100:49:@1232.4]
  reg  _T_113; // @[package.scala 48:56:@1233.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@1235.4]
  wire  _T_118; // @[Controllers.scala 283:41:@1240.4]
  wire  _T_119; // @[Controllers.scala 283:59:@1241.4]
  wire  _T_121; // @[Controllers.scala 284:37:@1244.4]
  wire  _T_124; // @[package.scala 96:25:@1252.4 package.scala 96:25:@1253.4]
  wire  _T_126; // @[package.scala 100:49:@1254.4]
  reg  _T_129; // @[package.scala 48:56:@1255.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@1277.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@1279.4]
  reg  _T_153; // @[package.scala 48:56:@1280.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@1288.4 package.scala 96:25:@1289.4]
  wire  _T_158; // @[Controllers.scala 292:61:@1290.4]
  wire  _T_159; // @[Controllers.scala 292:24:@1291.4]
  SRFF active ( // @[Controllers.scala 261:22:@1188.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@1191.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@1225.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@1247.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@1259.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@1267.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@1283.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@1196.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@1197.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@1198.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@1199.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@1216.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@1230.4 package.scala 96:25:@1231.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@1232.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@1235.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@1240.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@1241.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@1244.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@1252.4 package.scala 96:25:@1253.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@1254.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@1279.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@1288.4 package.scala 96:25:@1289.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@1290.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@1291.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@1258.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@1293.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@1243.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@1246.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@1238.4]
  assign active_clock = clock; // @[:@1189.4]
  assign active_reset = reset; // @[:@1190.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@1201.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@1205.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@1206.4]
  assign done_clock = clock; // @[:@1192.4]
  assign done_reset = reset; // @[:@1193.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@1221.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@1214.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@1215.4]
  assign RetimeWrapper_clock = clock; // @[:@1226.4]
  assign RetimeWrapper_reset = reset; // @[:@1227.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@1229.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@1228.4]
  assign RetimeWrapper_1_clock = clock; // @[:@1248.4]
  assign RetimeWrapper_1_reset = reset; // @[:@1249.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@1251.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@1250.4]
  assign RetimeWrapper_2_clock = clock; // @[:@1260.4]
  assign RetimeWrapper_2_reset = reset; // @[:@1261.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@1263.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@1262.4]
  assign RetimeWrapper_3_clock = clock; // @[:@1268.4]
  assign RetimeWrapper_3_reset = reset; // @[:@1269.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@1271.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@1270.4]
  assign RetimeWrapper_4_clock = clock; // @[:@1284.4]
  assign RetimeWrapper_4_reset = reset; // @[:@1285.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@1287.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@1286.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module fix2fixBox( // @[:@1423.2]
  input  [31:0] io_a, // @[:@1426.4]
  output [31:0] io_b // @[:@1426.4]
);
  assign io_b = io_a; // @[Converter.scala 95:38:@1436.4]
endmodule
module _( // @[:@1438.2]
  input  [31:0] io_b, // @[:@1441.4]
  output [31:0] io_result // @[:@1441.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@1446.4]
  wire [31:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@1446.4]
  fix2fixBox fix2fixBox ( // @[BigIPZynq.scala 219:30:@1446.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 706:17:@1454.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@1449.4]
endmodule
module fix2fixBox_1( // @[:@1456.2]
  input  [31:0] io_a, // @[:@1459.4]
  output [7:0]  io_b // @[:@1459.4]
);
  assign io_b = io_a[7:0]; // @[Converter.scala 95:38:@1469.4]
endmodule
module x90( // @[:@1471.2]
  input  [31:0] io_b, // @[:@1474.4]
  output [7:0]  io_result // @[:@1474.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@1479.4]
  wire [7:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@1479.4]
  fix2fixBox_1 fix2fixBox ( // @[BigIPZynq.scala 219:30:@1479.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 706:17:@1487.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@1482.4]
endmodule
module fix2fixBox_2( // @[:@1489.2]
  input  [31:0] io_a, // @[:@1492.4]
  output [32:0] io_b // @[:@1492.4]
);
  wire  _T_20; // @[implicits.scala 69:16:@1499.4]
  assign _T_20 = io_a[31]; // @[implicits.scala 69:16:@1499.4]
  assign io_b = {_T_20,io_a}; // @[Converter.scala 95:38:@1504.4]
endmodule
module __1( // @[:@1506.2]
  input  [31:0] io_b, // @[:@1509.4]
  output [32:0] io_result // @[:@1509.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@1514.4]
  wire [32:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@1514.4]
  fix2fixBox_2 fix2fixBox ( // @[BigIPZynq.scala 219:30:@1514.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 706:17:@1522.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@1517.4]
endmodule
module RetimeWrapper_15( // @[:@1571.2]
  input         clock, // @[:@1572.4]
  input         reset, // @[:@1573.4]
  input         io_flow, // @[:@1574.4]
  input  [31:0] io_in, // @[:@1574.4]
  output [31:0] io_out // @[:@1574.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@1576.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@1576.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@1576.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@1576.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@1576.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@1576.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@1576.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@1589.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@1588.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@1587.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@1586.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@1585.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@1583.4]
endmodule
module fix2fixBox_4( // @[:@1591.2]
  input         clock, // @[:@1592.4]
  input         reset, // @[:@1593.4]
  input  [32:0] io_a, // @[:@1594.4]
  input         io_flow, // @[:@1594.4]
  output [31:0] io_b // @[:@1594.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@1604.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@1604.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@1604.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@1604.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@1604.4]
  RetimeWrapper_15 RetimeWrapper ( // @[package.scala 93:22:@1604.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@1611.4]
  assign RetimeWrapper_clock = clock; // @[:@1605.4]
  assign RetimeWrapper_reset = reset; // @[:@1606.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@1608.4]
  assign RetimeWrapper_io_in = io_a[31:0]; // @[package.scala 94:16:@1607.4]
endmodule
module x91_sum( // @[:@1613.2]
  input         clock, // @[:@1614.4]
  input         reset, // @[:@1615.4]
  input  [31:0] io_a, // @[:@1616.4]
  input  [31:0] io_b, // @[:@1616.4]
  output [31:0] io_result // @[:@1616.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@1624.4]
  wire [32:0] __io_result; // @[Math.scala 709:24:@1624.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@1631.4]
  wire [32:0] __1_io_result; // @[Math.scala 709:24:@1631.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@1649.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@1649.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@1649.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@1649.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@1649.4]
  wire [32:0] a_upcast_number; // @[Math.scala 712:22:@1629.4 Math.scala 713:14:@1630.4]
  wire [32:0] b_upcast_number; // @[Math.scala 712:22:@1636.4 Math.scala 713:14:@1637.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@1638.4]
  __1 _ ( // @[Math.scala 709:24:@1624.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __1 __1 ( // @[Math.scala 709:24:@1631.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_4 fix2fixBox ( // @[Math.scala 141:30:@1649.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@1629.4 Math.scala 713:14:@1630.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@1636.4 Math.scala 713:14:@1637.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@1638.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@1657.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@1627.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@1634.4]
  assign fix2fixBox_clock = clock; // @[:@1650.4]
  assign fix2fixBox_reset = reset; // @[:@1651.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@1652.4]
  assign fix2fixBox_io_flow = 1'h1; // @[Math.scala 145:26:@1655.4]
endmodule
module RetimeWrapper_18( // @[:@2110.2]
  input        clock, // @[:@2111.4]
  input        reset, // @[:@2112.4]
  input  [7:0] io_in, // @[:@2113.4]
  output [7:0] io_out // @[:@2113.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@2115.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@2115.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@2115.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@2115.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@2115.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@2115.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@2115.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@2128.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@2127.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@2126.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@2125.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@2124.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@2122.4]
endmodule
module x102_inr_Foreach_kernelx102_inr_Foreach_concrete1( // @[:@2226.2]
  input         clock, // @[:@2227.4]
  input         reset, // @[:@2228.4]
  output [3:0]  io_in_x84_a_0_wPort_0_ofs_0, // @[:@2229.4]
  output [63:0] io_in_x84_a_0_wPort_0_data_0, // @[:@2229.4]
  output        io_in_x84_a_0_wPort_0_en_0, // @[:@2229.4]
  output [63:0] io_in_instrctrs_1_cycs, // @[:@2229.4]
  output [63:0] io_in_instrctrs_1_iters, // @[:@2229.4]
  input         io_sigsIn_done, // @[:@2229.4]
  input         io_sigsIn_datapathEn, // @[:@2229.4]
  input         io_sigsIn_baseEn, // @[:@2229.4]
  input         io_sigsIn_break, // @[:@2229.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@2229.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@2229.4]
  input         io_rr // @[:@2229.4]
);
  wire  cycles_clock; // @[sm_x102_inr_Foreach.scala 58:26:@2268.4]
  wire  cycles_reset; // @[sm_x102_inr_Foreach.scala 58:26:@2268.4]
  wire  cycles_io_enable; // @[sm_x102_inr_Foreach.scala 58:26:@2268.4]
  wire [63:0] cycles_io_count; // @[sm_x102_inr_Foreach.scala 58:26:@2268.4]
  wire  iters_clock; // @[sm_x102_inr_Foreach.scala 59:25:@2271.4]
  wire  iters_reset; // @[sm_x102_inr_Foreach.scala 59:25:@2271.4]
  wire  iters_io_enable; // @[sm_x102_inr_Foreach.scala 59:25:@2271.4]
  wire [63:0] iters_io_count; // @[sm_x102_inr_Foreach.scala 59:25:@2271.4]
  wire [31:0] __io_b; // @[Math.scala 709:24:@2288.4]
  wire [31:0] __io_result; // @[Math.scala 709:24:@2288.4]
  wire [31:0] x90_1_io_b; // @[Math.scala 709:24:@2307.4]
  wire [7:0] x90_1_io_result; // @[Math.scala 709:24:@2307.4]
  wire  x91_sum_1_clock; // @[Math.scala 150:24:@2318.4]
  wire  x91_sum_1_reset; // @[Math.scala 150:24:@2318.4]
  wire [31:0] x91_sum_1_io_a; // @[Math.scala 150:24:@2318.4]
  wire [31:0] x91_sum_1_io_b; // @[Math.scala 150:24:@2318.4]
  wire [31:0] x91_sum_1_io_result; // @[Math.scala 150:24:@2318.4]
  wire [31:0] x92_1_io_b; // @[Math.scala 709:24:@2328.4]
  wire [7:0] x92_1_io_result; // @[Math.scala 709:24:@2328.4]
  wire  x93_sum_1_clock; // @[Math.scala 150:24:@2339.4]
  wire  x93_sum_1_reset; // @[Math.scala 150:24:@2339.4]
  wire [31:0] x93_sum_1_io_a; // @[Math.scala 150:24:@2339.4]
  wire [31:0] x93_sum_1_io_b; // @[Math.scala 150:24:@2339.4]
  wire [31:0] x93_sum_1_io_result; // @[Math.scala 150:24:@2339.4]
  wire [31:0] x94_1_io_b; // @[Math.scala 709:24:@2349.4]
  wire [7:0] x94_1_io_result; // @[Math.scala 709:24:@2349.4]
  wire  x95_sum_1_clock; // @[Math.scala 150:24:@2360.4]
  wire  x95_sum_1_reset; // @[Math.scala 150:24:@2360.4]
  wire [31:0] x95_sum_1_io_a; // @[Math.scala 150:24:@2360.4]
  wire [31:0] x95_sum_1_io_b; // @[Math.scala 150:24:@2360.4]
  wire [31:0] x95_sum_1_io_result; // @[Math.scala 150:24:@2360.4]
  wire [31:0] x96_1_io_b; // @[Math.scala 709:24:@2370.4]
  wire [7:0] x96_1_io_result; // @[Math.scala 709:24:@2370.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@2379.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@2379.4]
  wire [7:0] RetimeWrapper_io_in; // @[package.scala 93:22:@2379.4]
  wire [7:0] RetimeWrapper_io_out; // @[package.scala 93:22:@2379.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@2414.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@2414.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@2414.4]
  wire [31:0] RetimeWrapper_1_io_in; // @[package.scala 93:22:@2414.4]
  wire [31:0] RetimeWrapper_1_io_out; // @[package.scala 93:22:@2414.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@2423.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@2423.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@2423.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@2423.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@2423.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@2436.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@2436.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@2436.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@2436.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@2436.4]
  wire  _T_250; // @[package.scala 100:49:@2275.4]
  reg  _T_253; // @[package.scala 48:56:@2276.4]
  reg [31:0] _RAND_0;
  wire [31:0] b87_number; // @[Math.scala 712:22:@2293.4 Math.scala 713:14:@2294.4]
  wire  _T_268; // @[FixedPoint.scala 50:25:@2299.4]
  wire [1:0] _T_272; // @[Bitwise.scala 72:12:@2301.4]
  wire [29:0] _T_273; // @[FixedPoint.scala 18:52:@2302.4]
  wire [7:0] x92_number; // @[Math.scala 712:22:@2333.4 Math.scala 713:14:@2334.4]
  wire [7:0] x151_x90_D1_number; // @[package.scala 96:25:@2384.4 package.scala 96:25:@2385.4]
  wire [7:0] x96_number; // @[Math.scala 712:22:@2375.4 Math.scala 713:14:@2376.4]
  wire [7:0] x94_number; // @[Math.scala 712:22:@2354.4 Math.scala 713:14:@2355.4]
  wire [31:0] _T_350; // @[Cat.scala 30:58:@2407.4]
  wire  _T_365; // @[sm_x102_inr_Foreach.scala 94:95:@2433.4]
  wire  _T_369; // @[package.scala 96:25:@2441.4 package.scala 96:25:@2442.4]
  wire  _T_371; // @[implicits.scala 55:10:@2443.4]
  wire  _T_372; // @[sm_x102_inr_Foreach.scala 94:112:@2444.4]
  wire  _T_374; // @[sm_x102_inr_Foreach.scala 94:199:@2446.4]
  wire  x153_b88_D1; // @[package.scala 96:25:@2428.4 package.scala 96:25:@2429.4]
  wire [31:0] x152_x89_D1_number; // @[package.scala 96:25:@2419.4 package.scala 96:25:@2420.4]
  InstrumentationCounter cycles ( // @[sm_x102_inr_Foreach.scala 58:26:@2268.4]
    .clock(cycles_clock),
    .reset(cycles_reset),
    .io_enable(cycles_io_enable),
    .io_count(cycles_io_count)
  );
  InstrumentationCounter iters ( // @[sm_x102_inr_Foreach.scala 59:25:@2271.4]
    .clock(iters_clock),
    .reset(iters_reset),
    .io_enable(iters_io_enable),
    .io_count(iters_io_count)
  );
  _ _ ( // @[Math.scala 709:24:@2288.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  x90 x90_1 ( // @[Math.scala 709:24:@2307.4]
    .io_b(x90_1_io_b),
    .io_result(x90_1_io_result)
  );
  x91_sum x91_sum_1 ( // @[Math.scala 150:24:@2318.4]
    .clock(x91_sum_1_clock),
    .reset(x91_sum_1_reset),
    .io_a(x91_sum_1_io_a),
    .io_b(x91_sum_1_io_b),
    .io_result(x91_sum_1_io_result)
  );
  x90 x92_1 ( // @[Math.scala 709:24:@2328.4]
    .io_b(x92_1_io_b),
    .io_result(x92_1_io_result)
  );
  x91_sum x93_sum_1 ( // @[Math.scala 150:24:@2339.4]
    .clock(x93_sum_1_clock),
    .reset(x93_sum_1_reset),
    .io_a(x93_sum_1_io_a),
    .io_b(x93_sum_1_io_b),
    .io_result(x93_sum_1_io_result)
  );
  x90 x94_1 ( // @[Math.scala 709:24:@2349.4]
    .io_b(x94_1_io_b),
    .io_result(x94_1_io_result)
  );
  x91_sum x95_sum_1 ( // @[Math.scala 150:24:@2360.4]
    .clock(x95_sum_1_clock),
    .reset(x95_sum_1_reset),
    .io_a(x95_sum_1_io_a),
    .io_b(x95_sum_1_io_b),
    .io_result(x95_sum_1_io_result)
  );
  x90 x96_1 ( // @[Math.scala 709:24:@2370.4]
    .io_b(x96_1_io_b),
    .io_result(x96_1_io_result)
  );
  RetimeWrapper_18 RetimeWrapper ( // @[package.scala 93:22:@2379.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_15 RetimeWrapper_1 ( // @[package.scala 93:22:@2414.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@2423.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@2436.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  assign _T_250 = io_sigsIn_done == 1'h0; // @[package.scala 100:49:@2275.4]
  assign b87_number = __io_result; // @[Math.scala 712:22:@2293.4 Math.scala 713:14:@2294.4]
  assign _T_268 = b87_number[31]; // @[FixedPoint.scala 50:25:@2299.4]
  assign _T_272 = _T_268 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@2301.4]
  assign _T_273 = b87_number[31:2]; // @[FixedPoint.scala 18:52:@2302.4]
  assign x92_number = x92_1_io_result; // @[Math.scala 712:22:@2333.4 Math.scala 713:14:@2334.4]
  assign x151_x90_D1_number = RetimeWrapper_io_out; // @[package.scala 96:25:@2384.4 package.scala 96:25:@2385.4]
  assign x96_number = x96_1_io_result; // @[Math.scala 712:22:@2375.4 Math.scala 713:14:@2376.4]
  assign x94_number = x94_1_io_result; // @[Math.scala 712:22:@2354.4 Math.scala 713:14:@2355.4]
  assign _T_350 = {x96_number,x94_number,x92_number,x151_x90_D1_number}; // @[Cat.scala 30:58:@2407.4]
  assign _T_365 = ~ io_sigsIn_break; // @[sm_x102_inr_Foreach.scala 94:95:@2433.4]
  assign _T_369 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@2441.4 package.scala 96:25:@2442.4]
  assign _T_371 = io_rr ? _T_369 : 1'h0; // @[implicits.scala 55:10:@2443.4]
  assign _T_372 = _T_365 & _T_371; // @[sm_x102_inr_Foreach.scala 94:112:@2444.4]
  assign _T_374 = _T_372 & _T_365; // @[sm_x102_inr_Foreach.scala 94:199:@2446.4]
  assign x153_b88_D1 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@2428.4 package.scala 96:25:@2429.4]
  assign x152_x89_D1_number = RetimeWrapper_1_io_out; // @[package.scala 96:25:@2419.4 package.scala 96:25:@2420.4]
  assign io_in_x84_a_0_wPort_0_ofs_0 = x152_x89_D1_number[3:0]; // @[MemInterfaceType.scala 89:54:@2450.4]
  assign io_in_x84_a_0_wPort_0_data_0 = {32'h0,_T_350}; // @[MemInterfaceType.scala 90:56:@2451.4]
  assign io_in_x84_a_0_wPort_0_en_0 = _T_374 & x153_b88_D1; // @[MemInterfaceType.scala 93:57:@2453.4]
  assign io_in_instrctrs_1_cycs = cycles_io_count; // @[Ledger.scala 282:21:@2280.4]
  assign io_in_instrctrs_1_iters = iters_io_count; // @[Ledger.scala 283:22:@2281.4]
  assign cycles_clock = clock; // @[:@2269.4]
  assign cycles_reset = reset; // @[:@2270.4]
  assign cycles_io_enable = io_sigsIn_baseEn; // @[sm_x102_inr_Foreach.scala 60:24:@2274.4]
  assign iters_clock = clock; // @[:@2272.4]
  assign iters_reset = reset; // @[:@2273.4]
  assign iters_io_enable = io_sigsIn_done & _T_253; // @[sm_x102_inr_Foreach.scala 61:23:@2279.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 710:17:@2291.4]
  assign x90_1_io_b = __io_result; // @[Math.scala 710:17:@2310.4]
  assign x91_sum_1_clock = clock; // @[:@2319.4]
  assign x91_sum_1_reset = reset; // @[:@2320.4]
  assign x91_sum_1_io_a = __io_result; // @[Math.scala 151:17:@2321.4]
  assign x91_sum_1_io_b = 32'h1; // @[Math.scala 152:17:@2322.4]
  assign x92_1_io_b = x91_sum_1_io_result; // @[Math.scala 710:17:@2331.4]
  assign x93_sum_1_clock = clock; // @[:@2340.4]
  assign x93_sum_1_reset = reset; // @[:@2341.4]
  assign x93_sum_1_io_a = __io_result; // @[Math.scala 151:17:@2342.4]
  assign x93_sum_1_io_b = 32'h2; // @[Math.scala 152:17:@2343.4]
  assign x94_1_io_b = x93_sum_1_io_result; // @[Math.scala 710:17:@2352.4]
  assign x95_sum_1_clock = clock; // @[:@2361.4]
  assign x95_sum_1_reset = reset; // @[:@2362.4]
  assign x95_sum_1_io_a = __io_result; // @[Math.scala 151:17:@2363.4]
  assign x95_sum_1_io_b = 32'h3; // @[Math.scala 152:17:@2364.4]
  assign x96_1_io_b = x95_sum_1_io_result; // @[Math.scala 710:17:@2373.4]
  assign RetimeWrapper_clock = clock; // @[:@2380.4]
  assign RetimeWrapper_reset = reset; // @[:@2381.4]
  assign RetimeWrapper_io_in = x90_1_io_result; // @[package.scala 94:16:@2382.4]
  assign RetimeWrapper_1_clock = clock; // @[:@2415.4]
  assign RetimeWrapper_1_reset = reset; // @[:@2416.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@2418.4]
  assign RetimeWrapper_1_io_in = {_T_272,_T_273}; // @[package.scala 94:16:@2417.4]
  assign RetimeWrapper_2_clock = clock; // @[:@2424.4]
  assign RetimeWrapper_2_reset = reset; // @[:@2425.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@2427.4]
  assign RetimeWrapper_2_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@2426.4]
  assign RetimeWrapper_3_clock = clock; // @[:@2437.4]
  assign RetimeWrapper_3_reset = reset; // @[:@2438.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@2440.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@2439.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_253 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_253 <= 1'h0;
    end else begin
      _T_253 <= _T_250;
    end
  end
endmodule
module x119_outr_UnitPipe_sm( // @[:@2654.2]
  input   clock, // @[:@2655.4]
  input   reset, // @[:@2656.4]
  input   io_enable, // @[:@2657.4]
  output  io_done, // @[:@2657.4]
  input   io_parentAck, // @[:@2657.4]
  input   io_doneIn_0, // @[:@2657.4]
  output  io_enableOut_0, // @[:@2657.4]
  output  io_childAck_0, // @[:@2657.4]
  input   io_ctrCopyDone_0 // @[:@2657.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@2660.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@2660.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@2660.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@2660.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@2660.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@2660.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@2663.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@2663.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@2663.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@2663.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@2663.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@2663.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@2680.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@2680.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@2680.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@2680.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@2680.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@2680.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@2711.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@2711.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@2711.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@2711.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@2711.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@2725.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@2725.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@2725.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@2725.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@2725.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@2743.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@2743.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@2743.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@2743.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@2743.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@2780.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@2780.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@2780.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@2780.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@2780.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@2797.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@2797.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@2797.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@2797.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@2797.4]
  wire  _T_105; // @[Controllers.scala 165:35:@2695.4]
  wire  _T_107; // @[Controllers.scala 165:60:@2696.4]
  wire  _T_108; // @[Controllers.scala 165:58:@2697.4]
  wire  _T_110; // @[Controllers.scala 165:76:@2698.4]
  wire  _T_111; // @[Controllers.scala 165:74:@2699.4]
  wire  _T_115; // @[Controllers.scala 165:109:@2702.4]
  wire  _T_118; // @[Controllers.scala 165:141:@2704.4]
  wire  _T_126; // @[package.scala 96:25:@2716.4 package.scala 96:25:@2717.4]
  wire  _T_130; // @[Controllers.scala 167:54:@2719.4]
  wire  _T_131; // @[Controllers.scala 167:52:@2720.4]
  wire  _T_138; // @[package.scala 96:25:@2730.4 package.scala 96:25:@2731.4]
  wire  _T_156; // @[package.scala 96:25:@2748.4 package.scala 96:25:@2749.4]
  wire  _T_160; // @[Controllers.scala 169:67:@2751.4]
  wire  _T_161; // @[Controllers.scala 169:86:@2752.4]
  wire  _T_174; // @[Controllers.scala 213:68:@2766.4]
  wire  _T_176; // @[Controllers.scala 213:90:@2768.4]
  wire  _T_178; // @[Controllers.scala 213:132:@2770.4]
  reg  _T_186; // @[package.scala 48:56:@2776.4]
  reg [31:0] _RAND_0;
  wire  _T_187; // @[package.scala 100:41:@2778.4]
  reg  _T_200; // @[package.scala 48:56:@2794.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@2660.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@2663.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@2680.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@2711.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@2725.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@2743.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@2780.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@2797.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_105 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@2695.4]
  assign _T_107 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@2696.4]
  assign _T_108 = _T_105 & _T_107; // @[Controllers.scala 165:58:@2697.4]
  assign _T_110 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@2698.4]
  assign _T_111 = _T_108 & _T_110; // @[Controllers.scala 165:74:@2699.4]
  assign _T_115 = _T_111 & io_enable; // @[Controllers.scala 165:109:@2702.4]
  assign _T_118 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@2704.4]
  assign _T_126 = RetimeWrapper_io_out; // @[package.scala 96:25:@2716.4 package.scala 96:25:@2717.4]
  assign _T_130 = _T_126 == 1'h0; // @[Controllers.scala 167:54:@2719.4]
  assign _T_131 = io_doneIn_0 | _T_130; // @[Controllers.scala 167:52:@2720.4]
  assign _T_138 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@2730.4 package.scala 96:25:@2731.4]
  assign _T_156 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@2748.4 package.scala 96:25:@2749.4]
  assign _T_160 = _T_156 == 1'h0; // @[Controllers.scala 169:67:@2751.4]
  assign _T_161 = _T_160 & io_enable; // @[Controllers.scala 169:86:@2752.4]
  assign _T_174 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@2766.4]
  assign _T_176 = _T_174 & _T_105; // @[Controllers.scala 213:90:@2768.4]
  assign _T_178 = ~ done_0_io_output; // @[Controllers.scala 213:132:@2770.4]
  assign _T_187 = done_0_io_output & _T_186; // @[package.scala 100:41:@2778.4]
  assign io_done = RetimeWrapper_4_io_out; // @[Controllers.scala 245:13:@2804.4]
  assign io_enableOut_0 = _T_176 & _T_178; // @[Controllers.scala 213:55:@2774.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@2765.4]
  assign active_0_clock = clock; // @[:@2661.4]
  assign active_0_reset = reset; // @[:@2662.4]
  assign active_0_io_input_set = _T_115 & _T_118; // @[Controllers.scala 165:32:@2706.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@2710.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@2668.4]
  assign done_0_clock = clock; // @[:@2664.4]
  assign done_0_reset = reset; // @[:@2665.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_161; // @[Controllers.scala 169:30:@2756.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@2678.4 Controllers.scala 170:32:@2763.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@2669.4]
  assign iterDone_0_clock = clock; // @[:@2681.4]
  assign iterDone_0_reset = reset; // @[:@2682.4]
  assign iterDone_0_io_input_set = _T_131 & io_enable; // @[Controllers.scala 167:34:@2724.4]
  assign iterDone_0_io_input_reset = _T_138 | io_parentAck; // @[Controllers.scala 92:37:@2692.4 Controllers.scala 168:36:@2740.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@2683.4]
  assign RetimeWrapper_clock = clock; // @[:@2712.4]
  assign RetimeWrapper_reset = reset; // @[:@2713.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@2715.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@2714.4]
  assign RetimeWrapper_1_clock = clock; // @[:@2726.4]
  assign RetimeWrapper_1_reset = reset; // @[:@2727.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@2729.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@2728.4]
  assign RetimeWrapper_2_clock = clock; // @[:@2744.4]
  assign RetimeWrapper_2_reset = reset; // @[:@2745.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@2747.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@2746.4]
  assign RetimeWrapper_3_clock = clock; // @[:@2781.4]
  assign RetimeWrapper_3_reset = reset; // @[:@2782.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@2784.4]
  assign RetimeWrapper_3_io_in = _T_187 | io_parentAck; // @[package.scala 94:16:@2783.4]
  assign RetimeWrapper_4_clock = clock; // @[:@2798.4]
  assign RetimeWrapper_4_reset = reset; // @[:@2799.4]
  assign RetimeWrapper_4_io_flow = io_enable; // @[package.scala 95:18:@2801.4]
  assign RetimeWrapper_4_io_in = done_0_io_output & _T_200; // @[package.scala 94:16:@2800.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_186 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_200 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_186 <= 1'h0;
    end else begin
      _T_186 <= _T_110;
    end
    if (reset) begin
      _T_200 <= 1'h0;
    end else begin
      _T_200 <= _T_110;
    end
  end
endmodule
module SingleCounter_2( // @[:@2948.2]
  input         clock, // @[:@2949.4]
  input         reset, // @[:@2950.4]
  input         io_input_reset, // @[:@2951.4]
  input         io_input_enable, // @[:@2951.4]
  output [31:0] io_output_count_0, // @[:@2951.4]
  output        io_output_oobs_0, // @[:@2951.4]
  output        io_output_done // @[:@2951.4]
);
  wire  bases_0_clock; // @[Counter.scala 253:53:@2964.4]
  wire  bases_0_reset; // @[Counter.scala 253:53:@2964.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 253:53:@2964.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 253:53:@2964.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 253:53:@2964.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 253:53:@2964.4]
  wire  SRFF_clock; // @[Counter.scala 255:22:@2980.4]
  wire  SRFF_reset; // @[Counter.scala 255:22:@2980.4]
  wire  SRFF_io_input_set; // @[Counter.scala 255:22:@2980.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 255:22:@2980.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 255:22:@2980.4]
  wire  SRFF_io_output; // @[Counter.scala 255:22:@2980.4]
  wire  _T_36; // @[Counter.scala 256:45:@2983.4]
  wire [31:0] _T_48; // @[Counter.scala 279:52:@3008.4]
  wire [32:0] _T_50; // @[Counter.scala 283:33:@3009.4]
  wire [31:0] _T_51; // @[Counter.scala 283:33:@3010.4]
  wire [31:0] _T_52; // @[Counter.scala 283:33:@3011.4]
  wire  _T_57; // @[Counter.scala 285:18:@3013.4]
  wire [31:0] _T_68; // @[Counter.scala 291:115:@3021.4]
  wire [31:0] _T_71; // @[Counter.scala 291:152:@3024.4]
  wire [31:0] _T_72; // @[Counter.scala 291:74:@3025.4]
  wire  _T_75; // @[Counter.scala 314:102:@3029.4]
  wire  _T_77; // @[Counter.scala 314:130:@3030.4]
  FF bases_0 ( // @[Counter.scala 253:53:@2964.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 255:22:@2980.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 256:45:@2983.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 279:52:@3008.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@3009.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@3010.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 283:33:@3011.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh8); // @[Counter.scala 285:18:@3013.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 291:115:@3021.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 291:152:@3024.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 291:74:@3025.4]
  assign _T_75 = $signed(_T_48) < $signed(32'sh0); // @[Counter.scala 314:102:@3029.4]
  assign _T_77 = $signed(_T_48) >= $signed(32'sh8); // @[Counter.scala 314:130:@3030.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 296:28:@3028.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 314:60:@3032.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 325:20:@3034.4]
  assign bases_0_clock = clock; // @[:@2965.4]
  assign bases_0_reset = reset; // @[:@2966.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 291:31:@3027.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 273:27:@3006.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 276:29:@3007.4]
  assign SRFF_clock = clock; // @[:@2981.4]
  assign SRFF_reset = reset; // @[:@2982.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 256:23:@2985.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 257:25:@2987.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 258:30:@2988.4]
endmodule
module x104_ctrchain( // @[:@3039.2]
  input         clock, // @[:@3040.4]
  input         reset, // @[:@3041.4]
  input         io_input_reset, // @[:@3042.4]
  input         io_input_enable, // @[:@3042.4]
  output [31:0] io_output_counts_0, // @[:@3042.4]
  output        io_output_oobs_0, // @[:@3042.4]
  output        io_output_done // @[:@3042.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 505:46:@3044.4]
  wire  ctrs_0_reset; // @[Counter.scala 505:46:@3044.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 505:46:@3044.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 505:46:@3044.4]
  wire [31:0] ctrs_0_io_output_count_0; // @[Counter.scala 505:46:@3044.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 505:46:@3044.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 505:46:@3044.4]
  reg  wasDone; // @[Counter.scala 534:24:@3053.4]
  reg [31:0] _RAND_0;
  wire  _T_45; // @[Counter.scala 538:69:@3059.4]
  wire  _T_47; // @[Counter.scala 538:80:@3060.4]
  reg  doneLatch; // @[Counter.scala 542:26:@3065.4]
  reg [31:0] _RAND_1;
  wire  _T_54; // @[Counter.scala 543:48:@3066.4]
  wire  _T_55; // @[Counter.scala 543:19:@3067.4]
  SingleCounter_2 ctrs_0 ( // @[Counter.scala 505:46:@3044.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done)
  );
  assign _T_45 = io_input_enable & ctrs_0_io_output_done; // @[Counter.scala 538:69:@3059.4]
  assign _T_47 = wasDone == 1'h0; // @[Counter.scala 538:80:@3060.4]
  assign _T_54 = ctrs_0_io_output_done ? 1'h1 : doneLatch; // @[Counter.scala 543:48:@3066.4]
  assign _T_55 = io_input_reset ? 1'h0 : _T_54; // @[Counter.scala 543:19:@3067.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 549:32:@3069.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 550:30:@3071.4]
  assign io_output_done = _T_45 & _T_47; // @[Counter.scala 538:18:@3062.4]
  assign ctrs_0_clock = clock; // @[:@3045.4]
  assign ctrs_0_reset = reset; // @[:@3046.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 512:24:@3050.4]
  assign ctrs_0_io_input_enable = io_input_enable; // @[Counter.scala 516:33:@3051.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= ctrs_0_io_output_done;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (ctrs_0_io_output_done) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module RetimeWrapper_37( // @[:@3568.2]
  input         clock, // @[:@3569.4]
  input         reset, // @[:@3570.4]
  input         io_flow, // @[:@3571.4]
  input  [63:0] io_in, // @[:@3571.4]
  output [63:0] io_out // @[:@3571.4]
);
  wire [63:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@3573.4]
  wire [63:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@3573.4]
  wire [63:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@3573.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3573.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3573.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3573.4]
  RetimeShiftRegister #(.WIDTH(64), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@3573.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3586.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3585.4]
  assign sr_init = 64'h0; // @[RetimeShiftRegister.scala 19:16:@3584.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3583.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3582.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3580.4]
endmodule
module x118_inr_Foreach_kernelx118_inr_Foreach_concrete1( // @[:@3684.2]
  input          clock, // @[:@3685.4]
  input          reset, // @[:@3686.4]
  output [3:0]   io_in_x84_a_0_rPort_0_ofs_0, // @[:@3687.4]
  output         io_in_x84_a_0_rPort_0_en_0, // @[:@3687.4]
  output         io_in_x84_a_0_rPort_0_backpressure, // @[:@3687.4]
  input  [63:0]  io_in_x84_a_0_rPort_0_output_0, // @[:@3687.4]
  output         io_in_x82_TVALID, // @[:@3687.4]
  input          io_in_x82_TREADY, // @[:@3687.4]
  output [511:0] io_in_x82_TDATA, // @[:@3687.4]
  output [63:0]  io_in_x82_TSTRB, // @[:@3687.4]
  output [63:0]  io_in_x82_TKEEP, // @[:@3687.4]
  output         io_in_x82_TLAST, // @[:@3687.4]
  output [7:0]   io_in_x82_TID, // @[:@3687.4]
  output [7:0]   io_in_x82_TDEST, // @[:@3687.4]
  output [31:0]  io_in_x82_TUSER, // @[:@3687.4]
  output [63:0]  io_in_instrctrs_3_cycs, // @[:@3687.4]
  output [63:0]  io_in_instrctrs_3_iters, // @[:@3687.4]
  output [63:0]  io_in_instrctrs_3_stalls, // @[:@3687.4]
  output [63:0]  io_in_instrctrs_3_idles, // @[:@3687.4]
  input          io_sigsIn_done, // @[:@3687.4]
  input          io_sigsIn_backpressure, // @[:@3687.4]
  input          io_sigsIn_datapathEn, // @[:@3687.4]
  input          io_sigsIn_baseEn, // @[:@3687.4]
  input          io_sigsIn_break, // @[:@3687.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_0, // @[:@3687.4]
  input          io_sigsIn_cchainOutputs_0_oobs_0, // @[:@3687.4]
  input          io_rr // @[:@3687.4]
);
  wire  cycles_clock; // @[sm_x118_inr_Foreach.scala 63:26:@3726.4]
  wire  cycles_reset; // @[sm_x118_inr_Foreach.scala 63:26:@3726.4]
  wire  cycles_io_enable; // @[sm_x118_inr_Foreach.scala 63:26:@3726.4]
  wire [63:0] cycles_io_count; // @[sm_x118_inr_Foreach.scala 63:26:@3726.4]
  wire  iters_clock; // @[sm_x118_inr_Foreach.scala 64:25:@3729.4]
  wire  iters_reset; // @[sm_x118_inr_Foreach.scala 64:25:@3729.4]
  wire  iters_io_enable; // @[sm_x118_inr_Foreach.scala 64:25:@3729.4]
  wire [63:0] iters_io_count; // @[sm_x118_inr_Foreach.scala 64:25:@3729.4]
  wire  stalls_clock; // @[sm_x118_inr_Foreach.scala 67:26:@3738.4]
  wire  stalls_reset; // @[sm_x118_inr_Foreach.scala 67:26:@3738.4]
  wire  stalls_io_enable; // @[sm_x118_inr_Foreach.scala 67:26:@3738.4]
  wire [63:0] stalls_io_count; // @[sm_x118_inr_Foreach.scala 67:26:@3738.4]
  wire  idles_clock; // @[sm_x118_inr_Foreach.scala 68:25:@3741.4]
  wire  idles_reset; // @[sm_x118_inr_Foreach.scala 68:25:@3741.4]
  wire  idles_io_enable; // @[sm_x118_inr_Foreach.scala 68:25:@3741.4]
  wire [63:0] idles_io_count; // @[sm_x118_inr_Foreach.scala 68:25:@3741.4]
  wire [31:0] __io_b; // @[Math.scala 709:24:@3758.4]
  wire [31:0] __io_result; // @[Math.scala 709:24:@3758.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@4001.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@4001.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@4001.4]
  wire [63:0] RetimeWrapper_io_in; // @[package.scala 93:22:@4001.4]
  wire [63:0] RetimeWrapper_io_out; // @[package.scala 93:22:@4001.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@4010.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@4010.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@4010.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@4010.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@4010.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@4035.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@4035.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@4035.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@4035.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@4035.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@4044.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@4044.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@4044.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@4044.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@4044.4]
  wire  _T_288; // @[package.scala 100:49:@3733.4]
  reg  _T_291; // @[package.scala 48:56:@3734.4]
  reg [31:0] _RAND_0;
  wire  _T_293; // @[sm_x118_inr_Foreach.scala 69:46:@3744.4]
  wire  b106; // @[sm_x118_inr_Foreach.scala 73:18:@3766.4]
  wire [31:0] b105_number; // @[Math.scala 712:22:@3763.4 Math.scala 713:14:@3764.4]
  wire [31:0] _T_311; // @[Math.scala 499:37:@3772.4]
  wire  x107; // @[Math.scala 499:44:@3774.4]
  wire  _T_334; // @[sm_x118_inr_Foreach.scala 84:123:@3786.4]
  wire  _T_338; // @[implicits.scala 55:10:@3789.4]
  wire  _T_339; // @[sm_x118_inr_Foreach.scala 84:140:@3790.4]
  wire  x114_0; // @[FixedPoint.scala 19:42:@3807.4]
  wire  x114_1; // @[FixedPoint.scala 19:42:@3809.4]
  wire  x114_2; // @[FixedPoint.scala 19:42:@3811.4]
  wire  x114_3; // @[FixedPoint.scala 19:42:@3813.4]
  wire  x114_4; // @[FixedPoint.scala 19:42:@3815.4]
  wire  x114_5; // @[FixedPoint.scala 19:42:@3817.4]
  wire  x114_6; // @[FixedPoint.scala 19:42:@3819.4]
  wire  x114_7; // @[FixedPoint.scala 19:42:@3821.4]
  wire  x114_8; // @[FixedPoint.scala 19:42:@3823.4]
  wire  x114_9; // @[FixedPoint.scala 19:42:@3825.4]
  wire  x114_10; // @[FixedPoint.scala 19:42:@3827.4]
  wire  x114_11; // @[FixedPoint.scala 19:42:@3829.4]
  wire  x114_12; // @[FixedPoint.scala 19:42:@3831.4]
  wire  x114_13; // @[FixedPoint.scala 19:42:@3833.4]
  wire  x114_14; // @[FixedPoint.scala 19:42:@3835.4]
  wire  x114_15; // @[FixedPoint.scala 19:42:@3837.4]
  wire  x114_16; // @[FixedPoint.scala 19:42:@3839.4]
  wire  x114_17; // @[FixedPoint.scala 19:42:@3841.4]
  wire  x114_18; // @[FixedPoint.scala 19:42:@3843.4]
  wire  x114_19; // @[FixedPoint.scala 19:42:@3845.4]
  wire  x114_20; // @[FixedPoint.scala 19:42:@3847.4]
  wire  x114_21; // @[FixedPoint.scala 19:42:@3849.4]
  wire  x114_22; // @[FixedPoint.scala 19:42:@3851.4]
  wire  x114_23; // @[FixedPoint.scala 19:42:@3853.4]
  wire  x114_24; // @[FixedPoint.scala 19:42:@3855.4]
  wire  x114_25; // @[FixedPoint.scala 19:42:@3857.4]
  wire  x114_26; // @[FixedPoint.scala 19:42:@3859.4]
  wire  x114_27; // @[FixedPoint.scala 19:42:@3861.4]
  wire  x114_28; // @[FixedPoint.scala 19:42:@3863.4]
  wire  x114_29; // @[FixedPoint.scala 19:42:@3865.4]
  wire  x114_30; // @[FixedPoint.scala 19:42:@3867.4]
  wire  x114_31; // @[FixedPoint.scala 19:42:@3869.4]
  wire  x114_32; // @[FixedPoint.scala 19:42:@3871.4]
  wire  x114_33; // @[FixedPoint.scala 19:42:@3873.4]
  wire  x114_34; // @[FixedPoint.scala 19:42:@3875.4]
  wire  x114_35; // @[FixedPoint.scala 19:42:@3877.4]
  wire  x114_36; // @[FixedPoint.scala 19:42:@3879.4]
  wire  x114_37; // @[FixedPoint.scala 19:42:@3881.4]
  wire  x114_38; // @[FixedPoint.scala 19:42:@3883.4]
  wire  x114_39; // @[FixedPoint.scala 19:42:@3885.4]
  wire  x114_40; // @[FixedPoint.scala 19:42:@3887.4]
  wire  x114_41; // @[FixedPoint.scala 19:42:@3889.4]
  wire  x114_42; // @[FixedPoint.scala 19:42:@3891.4]
  wire  x114_43; // @[FixedPoint.scala 19:42:@3893.4]
  wire  x114_44; // @[FixedPoint.scala 19:42:@3895.4]
  wire  x114_45; // @[FixedPoint.scala 19:42:@3897.4]
  wire  x114_46; // @[FixedPoint.scala 19:42:@3899.4]
  wire  x114_47; // @[FixedPoint.scala 19:42:@3901.4]
  wire  x114_48; // @[FixedPoint.scala 19:42:@3903.4]
  wire  x114_49; // @[FixedPoint.scala 19:42:@3905.4]
  wire  x114_50; // @[FixedPoint.scala 19:42:@3907.4]
  wire  x114_51; // @[FixedPoint.scala 19:42:@3909.4]
  wire  x114_52; // @[FixedPoint.scala 19:42:@3911.4]
  wire  x114_53; // @[FixedPoint.scala 19:42:@3913.4]
  wire  x114_54; // @[FixedPoint.scala 19:42:@3915.4]
  wire  x114_55; // @[FixedPoint.scala 19:42:@3917.4]
  wire  x114_56; // @[FixedPoint.scala 19:42:@3919.4]
  wire  x114_57; // @[FixedPoint.scala 19:42:@3921.4]
  wire  x114_58; // @[FixedPoint.scala 19:42:@3923.4]
  wire  x114_59; // @[FixedPoint.scala 19:42:@3925.4]
  wire  x114_60; // @[FixedPoint.scala 19:42:@3927.4]
  wire  x114_61; // @[FixedPoint.scala 19:42:@3929.4]
  wire  x114_62; // @[FixedPoint.scala 19:42:@3931.4]
  wire  x114_63; // @[FixedPoint.scala 19:42:@3933.4]
  wire [7:0] _T_490; // @[Cat.scala 30:58:@3942.4]
  wire [15:0] _T_498; // @[Cat.scala 30:58:@3950.4]
  wire [7:0] _T_505; // @[Cat.scala 30:58:@3957.4]
  wire [31:0] _T_514; // @[Cat.scala 30:58:@3966.4]
  wire [7:0] _T_521; // @[Cat.scala 30:58:@3973.4]
  wire [15:0] _T_529; // @[Cat.scala 30:58:@3981.4]
  wire [7:0] _T_536; // @[Cat.scala 30:58:@3988.4]
  wire [31:0] _T_545; // @[Cat.scala 30:58:@3997.4]
  wire [63:0] _T_546; // @[Cat.scala 30:58:@3998.4]
  wire [511:0] x115_number; // @[sm_x118_inr_Foreach.scala 91:22:@3935.4 sm_x118_inr_Foreach.scala 92:14:@3999.4]
  wire  x155_x113_D2; // @[package.scala 96:25:@4015.4 package.scala 96:25:@4016.4]
  wire [63:0] x154_x108_D2_number; // @[package.scala 96:25:@4006.4 package.scala 96:25:@4007.4]
  wire [720:0] x116_tuple; // @[Cat.scala 30:58:@4032.4]
  wire  _T_581; // @[package.scala 96:25:@4049.4 package.scala 96:25:@4050.4]
  wire  _T_583; // @[implicits.scala 55:10:@4051.4]
  wire  x156_b106_D2; // @[package.scala 96:25:@4040.4 package.scala 96:25:@4041.4]
  wire  _T_584; // @[sm_x118_inr_Foreach.scala 101:110:@4052.4]
  wire [8:0] _T_590; // @[sm_x118_inr_Foreach.scala 106:34:@4063.4]
  wire [62:0] _T_592; // @[sm_x118_inr_Foreach.scala 108:32:@4067.4]
  InstrumentationCounter cycles ( // @[sm_x118_inr_Foreach.scala 63:26:@3726.4]
    .clock(cycles_clock),
    .reset(cycles_reset),
    .io_enable(cycles_io_enable),
    .io_count(cycles_io_count)
  );
  InstrumentationCounter iters ( // @[sm_x118_inr_Foreach.scala 64:25:@3729.4]
    .clock(iters_clock),
    .reset(iters_reset),
    .io_enable(iters_io_enable),
    .io_count(iters_io_count)
  );
  InstrumentationCounter stalls ( // @[sm_x118_inr_Foreach.scala 67:26:@3738.4]
    .clock(stalls_clock),
    .reset(stalls_reset),
    .io_enable(stalls_io_enable),
    .io_count(stalls_io_count)
  );
  InstrumentationCounter idles ( // @[sm_x118_inr_Foreach.scala 68:25:@3741.4]
    .clock(idles_clock),
    .reset(idles_reset),
    .io_enable(idles_io_enable),
    .io_count(idles_io_count)
  );
  _ _ ( // @[Math.scala 709:24:@3758.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  RetimeWrapper_37 RetimeWrapper ( // @[package.scala 93:22:@4001.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@4010.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_2 ( // @[package.scala 93:22:@4035.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_3 ( // @[package.scala 93:22:@4044.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  assign _T_288 = io_sigsIn_done == 1'h0; // @[package.scala 100:49:@3733.4]
  assign _T_293 = ~ io_in_x82_TREADY; // @[sm_x118_inr_Foreach.scala 69:46:@3744.4]
  assign b106 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x118_inr_Foreach.scala 73:18:@3766.4]
  assign b105_number = __io_result; // @[Math.scala 712:22:@3763.4 Math.scala 713:14:@3764.4]
  assign _T_311 = $signed(b105_number); // @[Math.scala 499:37:@3772.4]
  assign x107 = $signed(_T_311) == $signed(32'sh0); // @[Math.scala 499:44:@3774.4]
  assign _T_334 = ~ io_sigsIn_break; // @[sm_x118_inr_Foreach.scala 84:123:@3786.4]
  assign _T_338 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 55:10:@3789.4]
  assign _T_339 = _T_334 & _T_338; // @[sm_x118_inr_Foreach.scala 84:140:@3790.4]
  assign x114_0 = io_in_x84_a_0_rPort_0_output_0[0]; // @[FixedPoint.scala 19:42:@3807.4]
  assign x114_1 = io_in_x84_a_0_rPort_0_output_0[1]; // @[FixedPoint.scala 19:42:@3809.4]
  assign x114_2 = io_in_x84_a_0_rPort_0_output_0[2]; // @[FixedPoint.scala 19:42:@3811.4]
  assign x114_3 = io_in_x84_a_0_rPort_0_output_0[3]; // @[FixedPoint.scala 19:42:@3813.4]
  assign x114_4 = io_in_x84_a_0_rPort_0_output_0[4]; // @[FixedPoint.scala 19:42:@3815.4]
  assign x114_5 = io_in_x84_a_0_rPort_0_output_0[5]; // @[FixedPoint.scala 19:42:@3817.4]
  assign x114_6 = io_in_x84_a_0_rPort_0_output_0[6]; // @[FixedPoint.scala 19:42:@3819.4]
  assign x114_7 = io_in_x84_a_0_rPort_0_output_0[7]; // @[FixedPoint.scala 19:42:@3821.4]
  assign x114_8 = io_in_x84_a_0_rPort_0_output_0[8]; // @[FixedPoint.scala 19:42:@3823.4]
  assign x114_9 = io_in_x84_a_0_rPort_0_output_0[9]; // @[FixedPoint.scala 19:42:@3825.4]
  assign x114_10 = io_in_x84_a_0_rPort_0_output_0[10]; // @[FixedPoint.scala 19:42:@3827.4]
  assign x114_11 = io_in_x84_a_0_rPort_0_output_0[11]; // @[FixedPoint.scala 19:42:@3829.4]
  assign x114_12 = io_in_x84_a_0_rPort_0_output_0[12]; // @[FixedPoint.scala 19:42:@3831.4]
  assign x114_13 = io_in_x84_a_0_rPort_0_output_0[13]; // @[FixedPoint.scala 19:42:@3833.4]
  assign x114_14 = io_in_x84_a_0_rPort_0_output_0[14]; // @[FixedPoint.scala 19:42:@3835.4]
  assign x114_15 = io_in_x84_a_0_rPort_0_output_0[15]; // @[FixedPoint.scala 19:42:@3837.4]
  assign x114_16 = io_in_x84_a_0_rPort_0_output_0[16]; // @[FixedPoint.scala 19:42:@3839.4]
  assign x114_17 = io_in_x84_a_0_rPort_0_output_0[17]; // @[FixedPoint.scala 19:42:@3841.4]
  assign x114_18 = io_in_x84_a_0_rPort_0_output_0[18]; // @[FixedPoint.scala 19:42:@3843.4]
  assign x114_19 = io_in_x84_a_0_rPort_0_output_0[19]; // @[FixedPoint.scala 19:42:@3845.4]
  assign x114_20 = io_in_x84_a_0_rPort_0_output_0[20]; // @[FixedPoint.scala 19:42:@3847.4]
  assign x114_21 = io_in_x84_a_0_rPort_0_output_0[21]; // @[FixedPoint.scala 19:42:@3849.4]
  assign x114_22 = io_in_x84_a_0_rPort_0_output_0[22]; // @[FixedPoint.scala 19:42:@3851.4]
  assign x114_23 = io_in_x84_a_0_rPort_0_output_0[23]; // @[FixedPoint.scala 19:42:@3853.4]
  assign x114_24 = io_in_x84_a_0_rPort_0_output_0[24]; // @[FixedPoint.scala 19:42:@3855.4]
  assign x114_25 = io_in_x84_a_0_rPort_0_output_0[25]; // @[FixedPoint.scala 19:42:@3857.4]
  assign x114_26 = io_in_x84_a_0_rPort_0_output_0[26]; // @[FixedPoint.scala 19:42:@3859.4]
  assign x114_27 = io_in_x84_a_0_rPort_0_output_0[27]; // @[FixedPoint.scala 19:42:@3861.4]
  assign x114_28 = io_in_x84_a_0_rPort_0_output_0[28]; // @[FixedPoint.scala 19:42:@3863.4]
  assign x114_29 = io_in_x84_a_0_rPort_0_output_0[29]; // @[FixedPoint.scala 19:42:@3865.4]
  assign x114_30 = io_in_x84_a_0_rPort_0_output_0[30]; // @[FixedPoint.scala 19:42:@3867.4]
  assign x114_31 = io_in_x84_a_0_rPort_0_output_0[31]; // @[FixedPoint.scala 19:42:@3869.4]
  assign x114_32 = io_in_x84_a_0_rPort_0_output_0[32]; // @[FixedPoint.scala 19:42:@3871.4]
  assign x114_33 = io_in_x84_a_0_rPort_0_output_0[33]; // @[FixedPoint.scala 19:42:@3873.4]
  assign x114_34 = io_in_x84_a_0_rPort_0_output_0[34]; // @[FixedPoint.scala 19:42:@3875.4]
  assign x114_35 = io_in_x84_a_0_rPort_0_output_0[35]; // @[FixedPoint.scala 19:42:@3877.4]
  assign x114_36 = io_in_x84_a_0_rPort_0_output_0[36]; // @[FixedPoint.scala 19:42:@3879.4]
  assign x114_37 = io_in_x84_a_0_rPort_0_output_0[37]; // @[FixedPoint.scala 19:42:@3881.4]
  assign x114_38 = io_in_x84_a_0_rPort_0_output_0[38]; // @[FixedPoint.scala 19:42:@3883.4]
  assign x114_39 = io_in_x84_a_0_rPort_0_output_0[39]; // @[FixedPoint.scala 19:42:@3885.4]
  assign x114_40 = io_in_x84_a_0_rPort_0_output_0[40]; // @[FixedPoint.scala 19:42:@3887.4]
  assign x114_41 = io_in_x84_a_0_rPort_0_output_0[41]; // @[FixedPoint.scala 19:42:@3889.4]
  assign x114_42 = io_in_x84_a_0_rPort_0_output_0[42]; // @[FixedPoint.scala 19:42:@3891.4]
  assign x114_43 = io_in_x84_a_0_rPort_0_output_0[43]; // @[FixedPoint.scala 19:42:@3893.4]
  assign x114_44 = io_in_x84_a_0_rPort_0_output_0[44]; // @[FixedPoint.scala 19:42:@3895.4]
  assign x114_45 = io_in_x84_a_0_rPort_0_output_0[45]; // @[FixedPoint.scala 19:42:@3897.4]
  assign x114_46 = io_in_x84_a_0_rPort_0_output_0[46]; // @[FixedPoint.scala 19:42:@3899.4]
  assign x114_47 = io_in_x84_a_0_rPort_0_output_0[47]; // @[FixedPoint.scala 19:42:@3901.4]
  assign x114_48 = io_in_x84_a_0_rPort_0_output_0[48]; // @[FixedPoint.scala 19:42:@3903.4]
  assign x114_49 = io_in_x84_a_0_rPort_0_output_0[49]; // @[FixedPoint.scala 19:42:@3905.4]
  assign x114_50 = io_in_x84_a_0_rPort_0_output_0[50]; // @[FixedPoint.scala 19:42:@3907.4]
  assign x114_51 = io_in_x84_a_0_rPort_0_output_0[51]; // @[FixedPoint.scala 19:42:@3909.4]
  assign x114_52 = io_in_x84_a_0_rPort_0_output_0[52]; // @[FixedPoint.scala 19:42:@3911.4]
  assign x114_53 = io_in_x84_a_0_rPort_0_output_0[53]; // @[FixedPoint.scala 19:42:@3913.4]
  assign x114_54 = io_in_x84_a_0_rPort_0_output_0[54]; // @[FixedPoint.scala 19:42:@3915.4]
  assign x114_55 = io_in_x84_a_0_rPort_0_output_0[55]; // @[FixedPoint.scala 19:42:@3917.4]
  assign x114_56 = io_in_x84_a_0_rPort_0_output_0[56]; // @[FixedPoint.scala 19:42:@3919.4]
  assign x114_57 = io_in_x84_a_0_rPort_0_output_0[57]; // @[FixedPoint.scala 19:42:@3921.4]
  assign x114_58 = io_in_x84_a_0_rPort_0_output_0[58]; // @[FixedPoint.scala 19:42:@3923.4]
  assign x114_59 = io_in_x84_a_0_rPort_0_output_0[59]; // @[FixedPoint.scala 19:42:@3925.4]
  assign x114_60 = io_in_x84_a_0_rPort_0_output_0[60]; // @[FixedPoint.scala 19:42:@3927.4]
  assign x114_61 = io_in_x84_a_0_rPort_0_output_0[61]; // @[FixedPoint.scala 19:42:@3929.4]
  assign x114_62 = io_in_x84_a_0_rPort_0_output_0[62]; // @[FixedPoint.scala 19:42:@3931.4]
  assign x114_63 = io_in_x84_a_0_rPort_0_output_0[63]; // @[FixedPoint.scala 19:42:@3933.4]
  assign _T_490 = {x114_7,x114_6,x114_5,x114_4,x114_3,x114_2,x114_1,x114_0}; // @[Cat.scala 30:58:@3942.4]
  assign _T_498 = {x114_15,x114_14,x114_13,x114_12,x114_11,x114_10,x114_9,x114_8,_T_490}; // @[Cat.scala 30:58:@3950.4]
  assign _T_505 = {x114_23,x114_22,x114_21,x114_20,x114_19,x114_18,x114_17,x114_16}; // @[Cat.scala 30:58:@3957.4]
  assign _T_514 = {x114_31,x114_30,x114_29,x114_28,x114_27,x114_26,x114_25,x114_24,_T_505,_T_498}; // @[Cat.scala 30:58:@3966.4]
  assign _T_521 = {x114_39,x114_38,x114_37,x114_36,x114_35,x114_34,x114_33,x114_32}; // @[Cat.scala 30:58:@3973.4]
  assign _T_529 = {x114_47,x114_46,x114_45,x114_44,x114_43,x114_42,x114_41,x114_40,_T_521}; // @[Cat.scala 30:58:@3981.4]
  assign _T_536 = {x114_55,x114_54,x114_53,x114_52,x114_51,x114_50,x114_49,x114_48}; // @[Cat.scala 30:58:@3988.4]
  assign _T_545 = {x114_63,x114_62,x114_61,x114_60,x114_59,x114_58,x114_57,x114_56,_T_536,_T_529}; // @[Cat.scala 30:58:@3997.4]
  assign _T_546 = {_T_545,_T_514}; // @[Cat.scala 30:58:@3998.4]
  assign x115_number = {{448'd0}, _T_546}; // @[sm_x118_inr_Foreach.scala 91:22:@3935.4 sm_x118_inr_Foreach.scala 92:14:@3999.4]
  assign x155_x113_D2 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@4015.4 package.scala 96:25:@4016.4]
  assign x154_x108_D2_number = RetimeWrapper_io_out; // @[package.scala 96:25:@4006.4 package.scala 96:25:@4007.4]
  assign x116_tuple = {x154_x108_D2_number,8'h0,8'h0,x155_x113_D2,128'h0,x115_number}; // @[Cat.scala 30:58:@4032.4]
  assign _T_581 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@4049.4 package.scala 96:25:@4050.4]
  assign _T_583 = io_rr ? _T_581 : 1'h0; // @[implicits.scala 55:10:@4051.4]
  assign x156_b106_D2 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@4040.4 package.scala 96:25:@4041.4]
  assign _T_584 = _T_583 & x156_b106_D2; // @[sm_x118_inr_Foreach.scala 101:110:@4052.4]
  assign _T_590 = x116_tuple[657:649]; // @[sm_x118_inr_Foreach.scala 106:34:@4063.4]
  assign _T_592 = x116_tuple[720:658]; // @[sm_x118_inr_Foreach.scala 108:32:@4067.4]
  assign io_in_x84_a_0_rPort_0_ofs_0 = b105_number[3:0]; // @[MemInterfaceType.scala 107:54:@3793.4]
  assign io_in_x84_a_0_rPort_0_en_0 = _T_339 & b106; // @[MemInterfaceType.scala 110:79:@3795.4]
  assign io_in_x84_a_0_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@3794.4]
  assign io_in_x82_TVALID = _T_584 & io_sigsIn_backpressure; // @[sm_x118_inr_Foreach.scala 101:17:@4054.4]
  assign io_in_x82_TDATA = x116_tuple[511:0]; // @[sm_x118_inr_Foreach.scala 102:19:@4056.4]
  assign io_in_x82_TSTRB = x116_tuple[575:512]; // @[sm_x118_inr_Foreach.scala 103:19:@4058.4]
  assign io_in_x82_TKEEP = x116_tuple[639:576]; // @[sm_x118_inr_Foreach.scala 104:19:@4060.4]
  assign io_in_x82_TLAST = x116_tuple[640]; // @[sm_x118_inr_Foreach.scala 107:17:@4066.4]
  assign io_in_x82_TID = x116_tuple[648:641]; // @[sm_x118_inr_Foreach.scala 105:17:@4062.4]
  assign io_in_x82_TDEST = _T_590[7:0]; // @[sm_x118_inr_Foreach.scala 106:19:@4064.4]
  assign io_in_x82_TUSER = _T_592[31:0]; // @[sm_x118_inr_Foreach.scala 108:17:@4068.4]
  assign io_in_instrctrs_3_cycs = cycles_io_count; // @[Ledger.scala 282:21:@3750.4]
  assign io_in_instrctrs_3_iters = iters_io_count; // @[Ledger.scala 283:22:@3751.4]
  assign io_in_instrctrs_3_stalls = stalls_io_count; // @[Ledger.scala 284:23:@3752.4]
  assign io_in_instrctrs_3_idles = idles_io_count; // @[Ledger.scala 285:22:@3753.4]
  assign cycles_clock = clock; // @[:@3727.4]
  assign cycles_reset = reset; // @[:@3728.4]
  assign cycles_io_enable = io_sigsIn_baseEn; // @[sm_x118_inr_Foreach.scala 65:24:@3732.4]
  assign iters_clock = clock; // @[:@3730.4]
  assign iters_reset = reset; // @[:@3731.4]
  assign iters_io_enable = io_sigsIn_done & _T_291; // @[sm_x118_inr_Foreach.scala 66:23:@3737.4]
  assign stalls_clock = clock; // @[:@3739.4]
  assign stalls_reset = reset; // @[:@3740.4]
  assign stalls_io_enable = io_sigsIn_baseEn & _T_293; // @[sm_x118_inr_Foreach.scala 69:24:@3746.4]
  assign idles_clock = clock; // @[:@3742.4]
  assign idles_reset = reset; // @[:@3743.4]
  assign idles_io_enable = 1'h0; // @[sm_x118_inr_Foreach.scala 70:23:@3749.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 710:17:@3761.4]
  assign RetimeWrapper_clock = clock; // @[:@4002.4]
  assign RetimeWrapper_reset = reset; // @[:@4003.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@4005.4]
  assign RetimeWrapper_io_in = x107 ? 64'h2 : 64'h0; // @[package.scala 94:16:@4004.4]
  assign RetimeWrapper_1_clock = clock; // @[:@4011.4]
  assign RetimeWrapper_1_reset = reset; // @[:@4012.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@4014.4]
  assign RetimeWrapper_1_io_in = $signed(_T_311) == $signed(32'sh7); // @[package.scala 94:16:@4013.4]
  assign RetimeWrapper_2_clock = clock; // @[:@4036.4]
  assign RetimeWrapper_2_reset = reset; // @[:@4037.4]
  assign RetimeWrapper_2_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@4039.4]
  assign RetimeWrapper_2_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@4038.4]
  assign RetimeWrapper_3_clock = clock; // @[:@4045.4]
  assign RetimeWrapper_3_reset = reset; // @[:@4046.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@4048.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@4047.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_291 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_291 <= 1'h0;
    end else begin
      _T_291 <= _T_288;
    end
  end
endmodule
module x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1( // @[:@4070.2]
  input          clock, // @[:@4071.4]
  input          reset, // @[:@4072.4]
  output [3:0]   io_in_x84_a_0_rPort_0_ofs_0, // @[:@4073.4]
  output         io_in_x84_a_0_rPort_0_en_0, // @[:@4073.4]
  output         io_in_x84_a_0_rPort_0_backpressure, // @[:@4073.4]
  input  [63:0]  io_in_x84_a_0_rPort_0_output_0, // @[:@4073.4]
  output         io_in_x82_TVALID, // @[:@4073.4]
  input          io_in_x82_TREADY, // @[:@4073.4]
  output [511:0] io_in_x82_TDATA, // @[:@4073.4]
  output [63:0]  io_in_x82_TSTRB, // @[:@4073.4]
  output [63:0]  io_in_x82_TKEEP, // @[:@4073.4]
  output         io_in_x82_TLAST, // @[:@4073.4]
  output [7:0]   io_in_x82_TID, // @[:@4073.4]
  output [7:0]   io_in_x82_TDEST, // @[:@4073.4]
  output [31:0]  io_in_x82_TUSER, // @[:@4073.4]
  output [63:0]  io_in_instrctrs_2_cycs, // @[:@4073.4]
  output [63:0]  io_in_instrctrs_2_iters, // @[:@4073.4]
  output [63:0]  io_in_instrctrs_3_cycs, // @[:@4073.4]
  output [63:0]  io_in_instrctrs_3_iters, // @[:@4073.4]
  output [63:0]  io_in_instrctrs_3_stalls, // @[:@4073.4]
  output [63:0]  io_in_instrctrs_3_idles, // @[:@4073.4]
  input          io_sigsIn_done, // @[:@4073.4]
  input          io_sigsIn_baseEn, // @[:@4073.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@4073.4]
  input          io_sigsIn_smChildAcks_0, // @[:@4073.4]
  output         io_sigsOut_smDoneIn_0, // @[:@4073.4]
  output         io_sigsOut_smCtrCopyDone_0, // @[:@4073.4]
  input          io_rr // @[:@4073.4]
);
  wire  cycles_clock; // @[sm_x119_outr_UnitPipe.scala 63:26:@4112.4]
  wire  cycles_reset; // @[sm_x119_outr_UnitPipe.scala 63:26:@4112.4]
  wire  cycles_io_enable; // @[sm_x119_outr_UnitPipe.scala 63:26:@4112.4]
  wire [63:0] cycles_io_count; // @[sm_x119_outr_UnitPipe.scala 63:26:@4112.4]
  wire  iters_clock; // @[sm_x119_outr_UnitPipe.scala 64:25:@4115.4]
  wire  iters_reset; // @[sm_x119_outr_UnitPipe.scala 64:25:@4115.4]
  wire  iters_io_enable; // @[sm_x119_outr_UnitPipe.scala 64:25:@4115.4]
  wire [63:0] iters_io_count; // @[sm_x119_outr_UnitPipe.scala 64:25:@4115.4]
  wire  x104_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@4128.4]
  wire  x104_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@4128.4]
  wire  x104_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@4128.4]
  wire  x104_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@4128.4]
  wire [31:0] x104_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@4128.4]
  wire  x104_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@4128.4]
  wire  x104_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@4128.4]
  wire  x118_inr_Foreach_sm_clock; // @[sm_x118_inr_Foreach.scala 33:18:@4180.4]
  wire  x118_inr_Foreach_sm_reset; // @[sm_x118_inr_Foreach.scala 33:18:@4180.4]
  wire  x118_inr_Foreach_sm_io_enable; // @[sm_x118_inr_Foreach.scala 33:18:@4180.4]
  wire  x118_inr_Foreach_sm_io_done; // @[sm_x118_inr_Foreach.scala 33:18:@4180.4]
  wire  x118_inr_Foreach_sm_io_doneLatch; // @[sm_x118_inr_Foreach.scala 33:18:@4180.4]
  wire  x118_inr_Foreach_sm_io_ctrDone; // @[sm_x118_inr_Foreach.scala 33:18:@4180.4]
  wire  x118_inr_Foreach_sm_io_datapathEn; // @[sm_x118_inr_Foreach.scala 33:18:@4180.4]
  wire  x118_inr_Foreach_sm_io_ctrInc; // @[sm_x118_inr_Foreach.scala 33:18:@4180.4]
  wire  x118_inr_Foreach_sm_io_ctrRst; // @[sm_x118_inr_Foreach.scala 33:18:@4180.4]
  wire  x118_inr_Foreach_sm_io_parentAck; // @[sm_x118_inr_Foreach.scala 33:18:@4180.4]
  wire  x118_inr_Foreach_sm_io_backpressure; // @[sm_x118_inr_Foreach.scala 33:18:@4180.4]
  wire  x118_inr_Foreach_sm_io_break; // @[sm_x118_inr_Foreach.scala 33:18:@4180.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@4208.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@4208.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@4208.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@4208.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@4208.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@4248.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@4248.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@4248.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@4248.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@4248.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@4256.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@4256.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@4256.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@4256.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@4256.4]
  wire  x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_clock; // @[sm_x118_inr_Foreach.scala 110:24:@4288.4]
  wire  x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_reset; // @[sm_x118_inr_Foreach.scala 110:24:@4288.4]
  wire [3:0] x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_x84_a_0_rPort_0_ofs_0; // @[sm_x118_inr_Foreach.scala 110:24:@4288.4]
  wire  x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_x84_a_0_rPort_0_en_0; // @[sm_x118_inr_Foreach.scala 110:24:@4288.4]
  wire  x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_x84_a_0_rPort_0_backpressure; // @[sm_x118_inr_Foreach.scala 110:24:@4288.4]
  wire [63:0] x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_x84_a_0_rPort_0_output_0; // @[sm_x118_inr_Foreach.scala 110:24:@4288.4]
  wire  x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_x82_TVALID; // @[sm_x118_inr_Foreach.scala 110:24:@4288.4]
  wire  x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_x82_TREADY; // @[sm_x118_inr_Foreach.scala 110:24:@4288.4]
  wire [511:0] x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_x82_TDATA; // @[sm_x118_inr_Foreach.scala 110:24:@4288.4]
  wire [63:0] x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_x82_TSTRB; // @[sm_x118_inr_Foreach.scala 110:24:@4288.4]
  wire [63:0] x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_x82_TKEEP; // @[sm_x118_inr_Foreach.scala 110:24:@4288.4]
  wire  x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_x82_TLAST; // @[sm_x118_inr_Foreach.scala 110:24:@4288.4]
  wire [7:0] x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_x82_TID; // @[sm_x118_inr_Foreach.scala 110:24:@4288.4]
  wire [7:0] x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_x82_TDEST; // @[sm_x118_inr_Foreach.scala 110:24:@4288.4]
  wire [31:0] x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_x82_TUSER; // @[sm_x118_inr_Foreach.scala 110:24:@4288.4]
  wire [63:0] x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_instrctrs_3_cycs; // @[sm_x118_inr_Foreach.scala 110:24:@4288.4]
  wire [63:0] x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_instrctrs_3_iters; // @[sm_x118_inr_Foreach.scala 110:24:@4288.4]
  wire [63:0] x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_instrctrs_3_stalls; // @[sm_x118_inr_Foreach.scala 110:24:@4288.4]
  wire [63:0] x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_instrctrs_3_idles; // @[sm_x118_inr_Foreach.scala 110:24:@4288.4]
  wire  x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_sigsIn_done; // @[sm_x118_inr_Foreach.scala 110:24:@4288.4]
  wire  x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_sigsIn_backpressure; // @[sm_x118_inr_Foreach.scala 110:24:@4288.4]
  wire  x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x118_inr_Foreach.scala 110:24:@4288.4]
  wire  x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_sigsIn_baseEn; // @[sm_x118_inr_Foreach.scala 110:24:@4288.4]
  wire  x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x118_inr_Foreach.scala 110:24:@4288.4]
  wire [31:0] x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x118_inr_Foreach.scala 110:24:@4288.4]
  wire  x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x118_inr_Foreach.scala 110:24:@4288.4]
  wire  x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_rr; // @[sm_x118_inr_Foreach.scala 110:24:@4288.4]
  wire  _T_288; // @[package.scala 100:49:@4119.4]
  reg  _T_291; // @[package.scala 48:56:@4120.4]
  reg [31:0] _RAND_0;
  wire  _T_355; // @[package.scala 96:25:@4213.4 package.scala 96:25:@4214.4]
  wire  _T_369; // @[package.scala 96:25:@4253.4 package.scala 96:25:@4254.4]
  wire  _T_375; // @[package.scala 96:25:@4261.4 package.scala 96:25:@4262.4]
  wire  _T_378; // @[SpatialBlocks.scala 110:93:@4264.4]
  wire  _T_380; // @[SpatialBlocks.scala 128:36:@4273.4]
  wire  _T_381; // @[SpatialBlocks.scala 128:78:@4274.4]
  InstrumentationCounter cycles ( // @[sm_x119_outr_UnitPipe.scala 63:26:@4112.4]
    .clock(cycles_clock),
    .reset(cycles_reset),
    .io_enable(cycles_io_enable),
    .io_count(cycles_io_count)
  );
  InstrumentationCounter iters ( // @[sm_x119_outr_UnitPipe.scala 64:25:@4115.4]
    .clock(iters_clock),
    .reset(iters_reset),
    .io_enable(iters_io_enable),
    .io_count(iters_io_count)
  );
  x104_ctrchain x104_ctrchain ( // @[SpatialBlocks.scala 37:22:@4128.4]
    .clock(x104_ctrchain_clock),
    .reset(x104_ctrchain_reset),
    .io_input_reset(x104_ctrchain_io_input_reset),
    .io_input_enable(x104_ctrchain_io_input_enable),
    .io_output_counts_0(x104_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x104_ctrchain_io_output_oobs_0),
    .io_output_done(x104_ctrchain_io_output_done)
  );
  x102_inr_Foreach_sm x118_inr_Foreach_sm ( // @[sm_x118_inr_Foreach.scala 33:18:@4180.4]
    .clock(x118_inr_Foreach_sm_clock),
    .reset(x118_inr_Foreach_sm_reset),
    .io_enable(x118_inr_Foreach_sm_io_enable),
    .io_done(x118_inr_Foreach_sm_io_done),
    .io_doneLatch(x118_inr_Foreach_sm_io_doneLatch),
    .io_ctrDone(x118_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x118_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x118_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x118_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x118_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x118_inr_Foreach_sm_io_backpressure),
    .io_break(x118_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@4208.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@4248.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@4256.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x118_inr_Foreach_kernelx118_inr_Foreach_concrete1 x118_inr_Foreach_kernelx118_inr_Foreach_concrete1 ( // @[sm_x118_inr_Foreach.scala 110:24:@4288.4]
    .clock(x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_clock),
    .reset(x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_reset),
    .io_in_x84_a_0_rPort_0_ofs_0(x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_x84_a_0_rPort_0_ofs_0),
    .io_in_x84_a_0_rPort_0_en_0(x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_x84_a_0_rPort_0_en_0),
    .io_in_x84_a_0_rPort_0_backpressure(x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_x84_a_0_rPort_0_backpressure),
    .io_in_x84_a_0_rPort_0_output_0(x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_x84_a_0_rPort_0_output_0),
    .io_in_x82_TVALID(x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_x82_TVALID),
    .io_in_x82_TREADY(x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_x82_TREADY),
    .io_in_x82_TDATA(x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_x82_TDATA),
    .io_in_x82_TSTRB(x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_x82_TSTRB),
    .io_in_x82_TKEEP(x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_x82_TKEEP),
    .io_in_x82_TLAST(x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_x82_TLAST),
    .io_in_x82_TID(x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_x82_TID),
    .io_in_x82_TDEST(x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_x82_TDEST),
    .io_in_x82_TUSER(x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_x82_TUSER),
    .io_in_instrctrs_3_cycs(x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_instrctrs_3_cycs),
    .io_in_instrctrs_3_iters(x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_instrctrs_3_iters),
    .io_in_instrctrs_3_stalls(x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_instrctrs_3_stalls),
    .io_in_instrctrs_3_idles(x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_instrctrs_3_idles),
    .io_sigsIn_done(x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_sigsIn_done),
    .io_sigsIn_backpressure(x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_baseEn(x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_sigsIn_baseEn),
    .io_sigsIn_break(x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_0(x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_rr(x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_rr)
  );
  assign _T_288 = io_sigsIn_done == 1'h0; // @[package.scala 100:49:@4119.4]
  assign _T_355 = RetimeWrapper_io_out; // @[package.scala 96:25:@4213.4 package.scala 96:25:@4214.4]
  assign _T_369 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@4253.4 package.scala 96:25:@4254.4]
  assign _T_375 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@4261.4 package.scala 96:25:@4262.4]
  assign _T_378 = ~ _T_375; // @[SpatialBlocks.scala 110:93:@4264.4]
  assign _T_380 = x118_inr_Foreach_sm_io_datapathEn; // @[SpatialBlocks.scala 128:36:@4273.4]
  assign _T_381 = ~ x118_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 128:78:@4274.4]
  assign io_in_x84_a_0_rPort_0_ofs_0 = x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_x84_a_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@4359.4]
  assign io_in_x84_a_0_rPort_0_en_0 = x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_x84_a_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@4358.4]
  assign io_in_x84_a_0_rPort_0_backpressure = x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_x84_a_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@4357.4]
  assign io_in_x82_TVALID = x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_x82_TVALID; // @[sm_x118_inr_Foreach.scala 51:22:@4369.4]
  assign io_in_x82_TDATA = x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_x82_TDATA; // @[sm_x118_inr_Foreach.scala 51:22:@4367.4]
  assign io_in_x82_TSTRB = x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_x82_TSTRB; // @[sm_x118_inr_Foreach.scala 51:22:@4366.4]
  assign io_in_x82_TKEEP = x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_x82_TKEEP; // @[sm_x118_inr_Foreach.scala 51:22:@4365.4]
  assign io_in_x82_TLAST = x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_x82_TLAST; // @[sm_x118_inr_Foreach.scala 51:22:@4364.4]
  assign io_in_x82_TID = x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_x82_TID; // @[sm_x118_inr_Foreach.scala 51:22:@4363.4]
  assign io_in_x82_TDEST = x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_x82_TDEST; // @[sm_x118_inr_Foreach.scala 51:22:@4362.4]
  assign io_in_x82_TUSER = x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_x82_TUSER; // @[sm_x118_inr_Foreach.scala 51:22:@4361.4]
  assign io_in_instrctrs_2_cycs = cycles_io_count; // @[Ledger.scala 282:21:@4124.4]
  assign io_in_instrctrs_2_iters = iters_io_count; // @[Ledger.scala 283:22:@4125.4]
  assign io_in_instrctrs_3_cycs = x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_instrctrs_3_cycs; // @[Ledger.scala 291:78:@4373.4]
  assign io_in_instrctrs_3_iters = x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_instrctrs_3_iters; // @[Ledger.scala 291:78:@4372.4]
  assign io_in_instrctrs_3_stalls = x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_instrctrs_3_stalls; // @[Ledger.scala 291:78:@4371.4]
  assign io_in_instrctrs_3_idles = x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_instrctrs_3_idles; // @[Ledger.scala 291:78:@4370.4]
  assign io_sigsOut_smDoneIn_0 = x118_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 127:53:@4271.4]
  assign io_sigsOut_smCtrCopyDone_0 = x118_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 139:125:@4287.4]
  assign cycles_clock = clock; // @[:@4113.4]
  assign cycles_reset = reset; // @[:@4114.4]
  assign cycles_io_enable = io_sigsIn_baseEn; // @[sm_x119_outr_UnitPipe.scala 65:24:@4118.4]
  assign iters_clock = clock; // @[:@4116.4]
  assign iters_reset = reset; // @[:@4117.4]
  assign iters_io_enable = io_sigsIn_done & _T_291; // @[sm_x119_outr_UnitPipe.scala 66:23:@4123.4]
  assign x104_ctrchain_clock = clock; // @[:@4129.4]
  assign x104_ctrchain_reset = reset; // @[:@4130.4]
  assign x104_ctrchain_io_input_reset = x118_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 130:103:@4286.4]
  assign x104_ctrchain_io_input_enable = x118_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 104:75:@4241.4 SpatialBlocks.scala 130:45:@4285.4]
  assign x118_inr_Foreach_sm_clock = clock; // @[:@4181.4]
  assign x118_inr_Foreach_sm_reset = reset; // @[:@4182.4]
  assign x118_inr_Foreach_sm_io_enable = _T_369 & _T_378; // @[SpatialBlocks.scala 112:18:@4268.4]
  assign x118_inr_Foreach_sm_io_ctrDone = io_rr ? _T_355 : 1'h0; // @[sm_x119_outr_UnitPipe.scala 73:38:@4216.4]
  assign x118_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 114:21:@4270.4]
  assign x118_inr_Foreach_sm_io_backpressure = io_in_x82_TREADY | x118_inr_Foreach_sm_io_doneLatch; // @[SpatialBlocks.scala 105:24:@4242.4]
  assign x118_inr_Foreach_sm_io_break = 1'h0; // @[sm_x119_outr_UnitPipe.scala 77:36:@4222.4]
  assign RetimeWrapper_clock = clock; // @[:@4209.4]
  assign RetimeWrapper_reset = reset; // @[:@4210.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@4212.4]
  assign RetimeWrapper_io_in = x104_ctrchain_io_output_done; // @[package.scala 94:16:@4211.4]
  assign RetimeWrapper_1_clock = clock; // @[:@4249.4]
  assign RetimeWrapper_1_reset = reset; // @[:@4250.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@4252.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@4251.4]
  assign RetimeWrapper_2_clock = clock; // @[:@4257.4]
  assign RetimeWrapper_2_reset = reset; // @[:@4258.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@4260.4]
  assign RetimeWrapper_2_io_in = x118_inr_Foreach_sm_io_done; // @[package.scala 94:16:@4259.4]
  assign x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_clock = clock; // @[:@4289.4]
  assign x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_reset = reset; // @[:@4290.4]
  assign x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_x84_a_0_rPort_0_output_0 = io_in_x84_a_0_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@4356.4]
  assign x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_in_x82_TREADY = io_in_x82_TREADY; // @[sm_x118_inr_Foreach.scala 51:22:@4368.4]
  assign x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_sigsIn_done = x118_inr_Foreach_sm_io_done; // @[sm_x118_inr_Foreach.scala 115:22:@4392.4]
  assign x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_sigsIn_backpressure = io_in_x82_TREADY | x118_inr_Foreach_sm_io_doneLatch; // @[sm_x118_inr_Foreach.scala 115:22:@4388.4]
  assign x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_380 & _T_381; // @[sm_x118_inr_Foreach.scala 115:22:@4386.4]
  assign x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_sigsIn_baseEn = _T_369 & _T_378; // @[sm_x118_inr_Foreach.scala 115:22:@4385.4]
  assign x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_sigsIn_break = x118_inr_Foreach_sm_io_break; // @[sm_x118_inr_Foreach.scala 115:22:@4384.4]
  assign x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = x104_ctrchain_io_output_counts_0; // @[sm_x118_inr_Foreach.scala 115:22:@4379.4]
  assign x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x104_ctrchain_io_output_oobs_0; // @[sm_x118_inr_Foreach.scala 115:22:@4378.4]
  assign x118_inr_Foreach_kernelx118_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x118_inr_Foreach.scala 114:18:@4374.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_291 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_291 <= 1'h0;
    end else begin
      _T_291 <= _T_288;
    end
  end
endmodule
module RootController_kernelRootController_concrete1( // @[:@4401.2]
  input          clock, // @[:@4402.4]
  input          reset, // @[:@4403.4]
  output         io_in_x82_TVALID, // @[:@4404.4]
  input          io_in_x82_TREADY, // @[:@4404.4]
  output [511:0] io_in_x82_TDATA, // @[:@4404.4]
  output [63:0]  io_in_x82_TSTRB, // @[:@4404.4]
  output [63:0]  io_in_x82_TKEEP, // @[:@4404.4]
  output         io_in_x82_TLAST, // @[:@4404.4]
  output [7:0]   io_in_x82_TID, // @[:@4404.4]
  output [7:0]   io_in_x82_TDEST, // @[:@4404.4]
  output [31:0]  io_in_x82_TUSER, // @[:@4404.4]
  output [63:0]  io_in_instrctrs_0_cycs, // @[:@4404.4]
  output [63:0]  io_in_instrctrs_0_iters, // @[:@4404.4]
  output [63:0]  io_in_instrctrs_1_cycs, // @[:@4404.4]
  output [63:0]  io_in_instrctrs_1_iters, // @[:@4404.4]
  output [63:0]  io_in_instrctrs_2_cycs, // @[:@4404.4]
  output [63:0]  io_in_instrctrs_2_iters, // @[:@4404.4]
  output [63:0]  io_in_instrctrs_3_cycs, // @[:@4404.4]
  output [63:0]  io_in_instrctrs_3_iters, // @[:@4404.4]
  output [63:0]  io_in_instrctrs_3_stalls, // @[:@4404.4]
  output [63:0]  io_in_instrctrs_3_idles, // @[:@4404.4]
  input          io_sigsIn_done, // @[:@4404.4]
  input          io_sigsIn_baseEn, // @[:@4404.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@4404.4]
  input          io_sigsIn_smEnableOuts_1, // @[:@4404.4]
  input          io_sigsIn_smChildAcks_0, // @[:@4404.4]
  input          io_sigsIn_smChildAcks_1, // @[:@4404.4]
  output         io_sigsOut_smDoneIn_0, // @[:@4404.4]
  output         io_sigsOut_smDoneIn_1, // @[:@4404.4]
  input          io_rr // @[:@4404.4]
);
  wire  cycles_clock; // @[sm_RootController.scala 58:26:@4432.4]
  wire  cycles_reset; // @[sm_RootController.scala 58:26:@4432.4]
  wire  cycles_io_enable; // @[sm_RootController.scala 58:26:@4432.4]
  wire [63:0] cycles_io_count; // @[sm_RootController.scala 58:26:@4432.4]
  wire  iters_clock; // @[sm_RootController.scala 59:25:@4435.4]
  wire  iters_reset; // @[sm_RootController.scala 59:25:@4435.4]
  wire  iters_io_enable; // @[sm_RootController.scala 59:25:@4435.4]
  wire [63:0] iters_io_count; // @[sm_RootController.scala 59:25:@4435.4]
  wire  x84_a_0_clock; // @[m_x84_a_0.scala 27:17:@4448.4]
  wire  x84_a_0_reset; // @[m_x84_a_0.scala 27:17:@4448.4]
  wire [3:0] x84_a_0_io_rPort_0_ofs_0; // @[m_x84_a_0.scala 27:17:@4448.4]
  wire  x84_a_0_io_rPort_0_en_0; // @[m_x84_a_0.scala 27:17:@4448.4]
  wire  x84_a_0_io_rPort_0_backpressure; // @[m_x84_a_0.scala 27:17:@4448.4]
  wire [63:0] x84_a_0_io_rPort_0_output_0; // @[m_x84_a_0.scala 27:17:@4448.4]
  wire [3:0] x84_a_0_io_wPort_0_ofs_0; // @[m_x84_a_0.scala 27:17:@4448.4]
  wire [63:0] x84_a_0_io_wPort_0_data_0; // @[m_x84_a_0.scala 27:17:@4448.4]
  wire  x84_a_0_io_wPort_0_en_0; // @[m_x84_a_0.scala 27:17:@4448.4]
  wire  x86_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@4465.4]
  wire  x86_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@4465.4]
  wire  x86_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@4465.4]
  wire  x86_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@4465.4]
  wire [31:0] x86_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@4465.4]
  wire  x86_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@4465.4]
  wire  x86_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@4465.4]
  wire  x102_inr_Foreach_sm_clock; // @[sm_x102_inr_Foreach.scala 32:18:@4517.4]
  wire  x102_inr_Foreach_sm_reset; // @[sm_x102_inr_Foreach.scala 32:18:@4517.4]
  wire  x102_inr_Foreach_sm_io_enable; // @[sm_x102_inr_Foreach.scala 32:18:@4517.4]
  wire  x102_inr_Foreach_sm_io_done; // @[sm_x102_inr_Foreach.scala 32:18:@4517.4]
  wire  x102_inr_Foreach_sm_io_doneLatch; // @[sm_x102_inr_Foreach.scala 32:18:@4517.4]
  wire  x102_inr_Foreach_sm_io_ctrDone; // @[sm_x102_inr_Foreach.scala 32:18:@4517.4]
  wire  x102_inr_Foreach_sm_io_datapathEn; // @[sm_x102_inr_Foreach.scala 32:18:@4517.4]
  wire  x102_inr_Foreach_sm_io_ctrInc; // @[sm_x102_inr_Foreach.scala 32:18:@4517.4]
  wire  x102_inr_Foreach_sm_io_ctrRst; // @[sm_x102_inr_Foreach.scala 32:18:@4517.4]
  wire  x102_inr_Foreach_sm_io_parentAck; // @[sm_x102_inr_Foreach.scala 32:18:@4517.4]
  wire  x102_inr_Foreach_sm_io_backpressure; // @[sm_x102_inr_Foreach.scala 32:18:@4517.4]
  wire  x102_inr_Foreach_sm_io_break; // @[sm_x102_inr_Foreach.scala 32:18:@4517.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@4545.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@4545.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@4545.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@4545.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@4545.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@4585.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@4585.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@4585.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@4585.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@4585.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@4593.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@4593.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@4593.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@4593.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@4593.4]
  wire  x102_inr_Foreach_kernelx102_inr_Foreach_concrete1_clock; // @[sm_x102_inr_Foreach.scala 96:24:@4624.4]
  wire  x102_inr_Foreach_kernelx102_inr_Foreach_concrete1_reset; // @[sm_x102_inr_Foreach.scala 96:24:@4624.4]
  wire [3:0] x102_inr_Foreach_kernelx102_inr_Foreach_concrete1_io_in_x84_a_0_wPort_0_ofs_0; // @[sm_x102_inr_Foreach.scala 96:24:@4624.4]
  wire [63:0] x102_inr_Foreach_kernelx102_inr_Foreach_concrete1_io_in_x84_a_0_wPort_0_data_0; // @[sm_x102_inr_Foreach.scala 96:24:@4624.4]
  wire  x102_inr_Foreach_kernelx102_inr_Foreach_concrete1_io_in_x84_a_0_wPort_0_en_0; // @[sm_x102_inr_Foreach.scala 96:24:@4624.4]
  wire [63:0] x102_inr_Foreach_kernelx102_inr_Foreach_concrete1_io_in_instrctrs_1_cycs; // @[sm_x102_inr_Foreach.scala 96:24:@4624.4]
  wire [63:0] x102_inr_Foreach_kernelx102_inr_Foreach_concrete1_io_in_instrctrs_1_iters; // @[sm_x102_inr_Foreach.scala 96:24:@4624.4]
  wire  x102_inr_Foreach_kernelx102_inr_Foreach_concrete1_io_sigsIn_done; // @[sm_x102_inr_Foreach.scala 96:24:@4624.4]
  wire  x102_inr_Foreach_kernelx102_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x102_inr_Foreach.scala 96:24:@4624.4]
  wire  x102_inr_Foreach_kernelx102_inr_Foreach_concrete1_io_sigsIn_baseEn; // @[sm_x102_inr_Foreach.scala 96:24:@4624.4]
  wire  x102_inr_Foreach_kernelx102_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x102_inr_Foreach.scala 96:24:@4624.4]
  wire [31:0] x102_inr_Foreach_kernelx102_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x102_inr_Foreach.scala 96:24:@4624.4]
  wire  x102_inr_Foreach_kernelx102_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x102_inr_Foreach.scala 96:24:@4624.4]
  wire  x102_inr_Foreach_kernelx102_inr_Foreach_concrete1_io_rr; // @[sm_x102_inr_Foreach.scala 96:24:@4624.4]
  wire  x119_outr_UnitPipe_sm_clock; // @[sm_x119_outr_UnitPipe.scala 33:18:@4755.4]
  wire  x119_outr_UnitPipe_sm_reset; // @[sm_x119_outr_UnitPipe.scala 33:18:@4755.4]
  wire  x119_outr_UnitPipe_sm_io_enable; // @[sm_x119_outr_UnitPipe.scala 33:18:@4755.4]
  wire  x119_outr_UnitPipe_sm_io_done; // @[sm_x119_outr_UnitPipe.scala 33:18:@4755.4]
  wire  x119_outr_UnitPipe_sm_io_parentAck; // @[sm_x119_outr_UnitPipe.scala 33:18:@4755.4]
  wire  x119_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x119_outr_UnitPipe.scala 33:18:@4755.4]
  wire  x119_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x119_outr_UnitPipe.scala 33:18:@4755.4]
  wire  x119_outr_UnitPipe_sm_io_childAck_0; // @[sm_x119_outr_UnitPipe.scala 33:18:@4755.4]
  wire  x119_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x119_outr_UnitPipe.scala 33:18:@4755.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@4807.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@4807.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@4807.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@4807.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@4807.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@4815.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@4815.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@4815.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@4815.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@4815.4]
  wire  x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_clock; // @[sm_x119_outr_UnitPipe.scala 82:24:@4842.4]
  wire  x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_reset; // @[sm_x119_outr_UnitPipe.scala 82:24:@4842.4]
  wire [3:0] x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_x84_a_0_rPort_0_ofs_0; // @[sm_x119_outr_UnitPipe.scala 82:24:@4842.4]
  wire  x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_x84_a_0_rPort_0_en_0; // @[sm_x119_outr_UnitPipe.scala 82:24:@4842.4]
  wire  x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_x84_a_0_rPort_0_backpressure; // @[sm_x119_outr_UnitPipe.scala 82:24:@4842.4]
  wire [63:0] x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_x84_a_0_rPort_0_output_0; // @[sm_x119_outr_UnitPipe.scala 82:24:@4842.4]
  wire  x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_x82_TVALID; // @[sm_x119_outr_UnitPipe.scala 82:24:@4842.4]
  wire  x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_x82_TREADY; // @[sm_x119_outr_UnitPipe.scala 82:24:@4842.4]
  wire [511:0] x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_x82_TDATA; // @[sm_x119_outr_UnitPipe.scala 82:24:@4842.4]
  wire [63:0] x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_x82_TSTRB; // @[sm_x119_outr_UnitPipe.scala 82:24:@4842.4]
  wire [63:0] x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_x82_TKEEP; // @[sm_x119_outr_UnitPipe.scala 82:24:@4842.4]
  wire  x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_x82_TLAST; // @[sm_x119_outr_UnitPipe.scala 82:24:@4842.4]
  wire [7:0] x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_x82_TID; // @[sm_x119_outr_UnitPipe.scala 82:24:@4842.4]
  wire [7:0] x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_x82_TDEST; // @[sm_x119_outr_UnitPipe.scala 82:24:@4842.4]
  wire [31:0] x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_x82_TUSER; // @[sm_x119_outr_UnitPipe.scala 82:24:@4842.4]
  wire [63:0] x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_instrctrs_2_cycs; // @[sm_x119_outr_UnitPipe.scala 82:24:@4842.4]
  wire [63:0] x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_instrctrs_2_iters; // @[sm_x119_outr_UnitPipe.scala 82:24:@4842.4]
  wire [63:0] x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_instrctrs_3_cycs; // @[sm_x119_outr_UnitPipe.scala 82:24:@4842.4]
  wire [63:0] x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_instrctrs_3_iters; // @[sm_x119_outr_UnitPipe.scala 82:24:@4842.4]
  wire [63:0] x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_instrctrs_3_stalls; // @[sm_x119_outr_UnitPipe.scala 82:24:@4842.4]
  wire [63:0] x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_instrctrs_3_idles; // @[sm_x119_outr_UnitPipe.scala 82:24:@4842.4]
  wire  x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_sigsIn_done; // @[sm_x119_outr_UnitPipe.scala 82:24:@4842.4]
  wire  x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_sigsIn_baseEn; // @[sm_x119_outr_UnitPipe.scala 82:24:@4842.4]
  wire  x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x119_outr_UnitPipe.scala 82:24:@4842.4]
  wire  x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x119_outr_UnitPipe.scala 82:24:@4842.4]
  wire  x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x119_outr_UnitPipe.scala 82:24:@4842.4]
  wire  x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x119_outr_UnitPipe.scala 82:24:@4842.4]
  wire  x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_rr; // @[sm_x119_outr_UnitPipe.scala 82:24:@4842.4]
  wire  _T_162; // @[package.scala 100:49:@4439.4]
  reg  _T_165; // @[package.scala 48:56:@4440.4]
  reg [31:0] _RAND_0;
  wire  _T_230; // @[package.scala 96:25:@4550.4 package.scala 96:25:@4551.4]
  wire  _T_245; // @[package.scala 96:25:@4590.4 package.scala 96:25:@4591.4]
  wire  _T_251; // @[package.scala 96:25:@4598.4 package.scala 96:25:@4599.4]
  wire  _T_254; // @[SpatialBlocks.scala 110:93:@4601.4]
  wire  _T_256; // @[SpatialBlocks.scala 128:36:@4610.4]
  wire  _T_257; // @[SpatialBlocks.scala 128:78:@4611.4]
  wire  _T_333; // @[package.scala 96:25:@4812.4 package.scala 96:25:@4813.4]
  wire  _T_339; // @[package.scala 96:25:@4820.4 package.scala 96:25:@4821.4]
  wire  _T_342; // @[SpatialBlocks.scala 110:93:@4823.4]
  InstrumentationCounter cycles ( // @[sm_RootController.scala 58:26:@4432.4]
    .clock(cycles_clock),
    .reset(cycles_reset),
    .io_enable(cycles_io_enable),
    .io_count(cycles_io_count)
  );
  InstrumentationCounter iters ( // @[sm_RootController.scala 59:25:@4435.4]
    .clock(iters_clock),
    .reset(iters_reset),
    .io_enable(iters_io_enable),
    .io_count(iters_io_count)
  );
  x84_a_0 x84_a_0 ( // @[m_x84_a_0.scala 27:17:@4448.4]
    .clock(x84_a_0_clock),
    .reset(x84_a_0_reset),
    .io_rPort_0_ofs_0(x84_a_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x84_a_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x84_a_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x84_a_0_io_rPort_0_output_0),
    .io_wPort_0_ofs_0(x84_a_0_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x84_a_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x84_a_0_io_wPort_0_en_0)
  );
  x86_ctrchain x86_ctrchain ( // @[SpatialBlocks.scala 37:22:@4465.4]
    .clock(x86_ctrchain_clock),
    .reset(x86_ctrchain_reset),
    .io_input_reset(x86_ctrchain_io_input_reset),
    .io_input_enable(x86_ctrchain_io_input_enable),
    .io_output_counts_0(x86_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x86_ctrchain_io_output_oobs_0),
    .io_output_done(x86_ctrchain_io_output_done)
  );
  x102_inr_Foreach_sm x102_inr_Foreach_sm ( // @[sm_x102_inr_Foreach.scala 32:18:@4517.4]
    .clock(x102_inr_Foreach_sm_clock),
    .reset(x102_inr_Foreach_sm_reset),
    .io_enable(x102_inr_Foreach_sm_io_enable),
    .io_done(x102_inr_Foreach_sm_io_done),
    .io_doneLatch(x102_inr_Foreach_sm_io_doneLatch),
    .io_ctrDone(x102_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x102_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x102_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x102_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x102_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x102_inr_Foreach_sm_io_backpressure),
    .io_break(x102_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@4545.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@4585.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@4593.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x102_inr_Foreach_kernelx102_inr_Foreach_concrete1 x102_inr_Foreach_kernelx102_inr_Foreach_concrete1 ( // @[sm_x102_inr_Foreach.scala 96:24:@4624.4]
    .clock(x102_inr_Foreach_kernelx102_inr_Foreach_concrete1_clock),
    .reset(x102_inr_Foreach_kernelx102_inr_Foreach_concrete1_reset),
    .io_in_x84_a_0_wPort_0_ofs_0(x102_inr_Foreach_kernelx102_inr_Foreach_concrete1_io_in_x84_a_0_wPort_0_ofs_0),
    .io_in_x84_a_0_wPort_0_data_0(x102_inr_Foreach_kernelx102_inr_Foreach_concrete1_io_in_x84_a_0_wPort_0_data_0),
    .io_in_x84_a_0_wPort_0_en_0(x102_inr_Foreach_kernelx102_inr_Foreach_concrete1_io_in_x84_a_0_wPort_0_en_0),
    .io_in_instrctrs_1_cycs(x102_inr_Foreach_kernelx102_inr_Foreach_concrete1_io_in_instrctrs_1_cycs),
    .io_in_instrctrs_1_iters(x102_inr_Foreach_kernelx102_inr_Foreach_concrete1_io_in_instrctrs_1_iters),
    .io_sigsIn_done(x102_inr_Foreach_kernelx102_inr_Foreach_concrete1_io_sigsIn_done),
    .io_sigsIn_datapathEn(x102_inr_Foreach_kernelx102_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_baseEn(x102_inr_Foreach_kernelx102_inr_Foreach_concrete1_io_sigsIn_baseEn),
    .io_sigsIn_break(x102_inr_Foreach_kernelx102_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_0(x102_inr_Foreach_kernelx102_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x102_inr_Foreach_kernelx102_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_rr(x102_inr_Foreach_kernelx102_inr_Foreach_concrete1_io_rr)
  );
  x119_outr_UnitPipe_sm x119_outr_UnitPipe_sm ( // @[sm_x119_outr_UnitPipe.scala 33:18:@4755.4]
    .clock(x119_outr_UnitPipe_sm_clock),
    .reset(x119_outr_UnitPipe_sm_reset),
    .io_enable(x119_outr_UnitPipe_sm_io_enable),
    .io_done(x119_outr_UnitPipe_sm_io_done),
    .io_parentAck(x119_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x119_outr_UnitPipe_sm_io_doneIn_0),
    .io_enableOut_0(x119_outr_UnitPipe_sm_io_enableOut_0),
    .io_childAck_0(x119_outr_UnitPipe_sm_io_childAck_0),
    .io_ctrCopyDone_0(x119_outr_UnitPipe_sm_io_ctrCopyDone_0)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@4807.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@4815.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1 x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1 ( // @[sm_x119_outr_UnitPipe.scala 82:24:@4842.4]
    .clock(x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_clock),
    .reset(x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_reset),
    .io_in_x84_a_0_rPort_0_ofs_0(x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_x84_a_0_rPort_0_ofs_0),
    .io_in_x84_a_0_rPort_0_en_0(x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_x84_a_0_rPort_0_en_0),
    .io_in_x84_a_0_rPort_0_backpressure(x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_x84_a_0_rPort_0_backpressure),
    .io_in_x84_a_0_rPort_0_output_0(x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_x84_a_0_rPort_0_output_0),
    .io_in_x82_TVALID(x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_x82_TVALID),
    .io_in_x82_TREADY(x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_x82_TREADY),
    .io_in_x82_TDATA(x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_x82_TDATA),
    .io_in_x82_TSTRB(x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_x82_TSTRB),
    .io_in_x82_TKEEP(x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_x82_TKEEP),
    .io_in_x82_TLAST(x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_x82_TLAST),
    .io_in_x82_TID(x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_x82_TID),
    .io_in_x82_TDEST(x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_x82_TDEST),
    .io_in_x82_TUSER(x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_x82_TUSER),
    .io_in_instrctrs_2_cycs(x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_instrctrs_2_cycs),
    .io_in_instrctrs_2_iters(x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_instrctrs_2_iters),
    .io_in_instrctrs_3_cycs(x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_instrctrs_3_cycs),
    .io_in_instrctrs_3_iters(x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_instrctrs_3_iters),
    .io_in_instrctrs_3_stalls(x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_instrctrs_3_stalls),
    .io_in_instrctrs_3_idles(x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_instrctrs_3_idles),
    .io_sigsIn_done(x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_sigsIn_done),
    .io_sigsIn_baseEn(x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_sigsIn_baseEn),
    .io_sigsIn_smEnableOuts_0(x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smCtrCopyDone_0(x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_rr(x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_rr)
  );
  assign _T_162 = io_sigsIn_done == 1'h0; // @[package.scala 100:49:@4439.4]
  assign _T_230 = RetimeWrapper_io_out; // @[package.scala 96:25:@4550.4 package.scala 96:25:@4551.4]
  assign _T_245 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@4590.4 package.scala 96:25:@4591.4]
  assign _T_251 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@4598.4 package.scala 96:25:@4599.4]
  assign _T_254 = ~ _T_251; // @[SpatialBlocks.scala 110:93:@4601.4]
  assign _T_256 = x102_inr_Foreach_sm_io_datapathEn; // @[SpatialBlocks.scala 128:36:@4610.4]
  assign _T_257 = ~ x102_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 128:78:@4611.4]
  assign _T_333 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@4812.4 package.scala 96:25:@4813.4]
  assign _T_339 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@4820.4 package.scala 96:25:@4821.4]
  assign _T_342 = ~ _T_339; // @[SpatialBlocks.scala 110:93:@4823.4]
  assign io_in_x82_TVALID = x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_x82_TVALID; // @[sm_x119_outr_UnitPipe.scala 51:22:@4923.4]
  assign io_in_x82_TDATA = x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_x82_TDATA; // @[sm_x119_outr_UnitPipe.scala 51:22:@4921.4]
  assign io_in_x82_TSTRB = x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_x82_TSTRB; // @[sm_x119_outr_UnitPipe.scala 51:22:@4920.4]
  assign io_in_x82_TKEEP = x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_x82_TKEEP; // @[sm_x119_outr_UnitPipe.scala 51:22:@4919.4]
  assign io_in_x82_TLAST = x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_x82_TLAST; // @[sm_x119_outr_UnitPipe.scala 51:22:@4918.4]
  assign io_in_x82_TID = x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_x82_TID; // @[sm_x119_outr_UnitPipe.scala 51:22:@4917.4]
  assign io_in_x82_TDEST = x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_x82_TDEST; // @[sm_x119_outr_UnitPipe.scala 51:22:@4916.4]
  assign io_in_x82_TUSER = x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_x82_TUSER; // @[sm_x119_outr_UnitPipe.scala 51:22:@4915.4]
  assign io_in_instrctrs_0_cycs = cycles_io_count; // @[Ledger.scala 282:21:@4444.4]
  assign io_in_instrctrs_0_iters = iters_io_count; // @[Ledger.scala 283:22:@4445.4]
  assign io_in_instrctrs_1_cycs = x102_inr_Foreach_kernelx102_inr_Foreach_concrete1_io_in_instrctrs_1_cycs; // @[Ledger.scala 291:78:@4693.4]
  assign io_in_instrctrs_1_iters = x102_inr_Foreach_kernelx102_inr_Foreach_concrete1_io_in_instrctrs_1_iters; // @[Ledger.scala 291:78:@4692.4]
  assign io_in_instrctrs_2_cycs = x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_instrctrs_2_cycs; // @[Ledger.scala 291:78:@4927.4]
  assign io_in_instrctrs_2_iters = x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_instrctrs_2_iters; // @[Ledger.scala 291:78:@4926.4]
  assign io_in_instrctrs_3_cycs = x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_instrctrs_3_cycs; // @[Ledger.scala 291:78:@4931.4]
  assign io_in_instrctrs_3_iters = x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_instrctrs_3_iters; // @[Ledger.scala 291:78:@4930.4]
  assign io_in_instrctrs_3_stalls = x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_instrctrs_3_stalls; // @[Ledger.scala 291:78:@4929.4]
  assign io_in_instrctrs_3_idles = x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_instrctrs_3_idles; // @[Ledger.scala 291:78:@4928.4]
  assign io_sigsOut_smDoneIn_0 = x102_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 127:53:@4608.4]
  assign io_sigsOut_smDoneIn_1 = x119_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 127:53:@4830.4]
  assign cycles_clock = clock; // @[:@4433.4]
  assign cycles_reset = reset; // @[:@4434.4]
  assign cycles_io_enable = io_sigsIn_baseEn; // @[sm_RootController.scala 60:24:@4438.4]
  assign iters_clock = clock; // @[:@4436.4]
  assign iters_reset = reset; // @[:@4437.4]
  assign iters_io_enable = io_sigsIn_done & _T_165; // @[sm_RootController.scala 61:23:@4443.4]
  assign x84_a_0_clock = clock; // @[:@4449.4]
  assign x84_a_0_reset = reset; // @[:@4450.4]
  assign x84_a_0_io_rPort_0_ofs_0 = x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_x84_a_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@4913.4]
  assign x84_a_0_io_rPort_0_en_0 = x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_x84_a_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@4912.4]
  assign x84_a_0_io_rPort_0_backpressure = x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_x84_a_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@4911.4]
  assign x84_a_0_io_wPort_0_ofs_0 = x102_inr_Foreach_kernelx102_inr_Foreach_concrete1_io_in_x84_a_0_wPort_0_ofs_0; // @[MemInterfaceType.scala 67:44:@4688.4]
  assign x84_a_0_io_wPort_0_data_0 = x102_inr_Foreach_kernelx102_inr_Foreach_concrete1_io_in_x84_a_0_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@4687.4]
  assign x84_a_0_io_wPort_0_en_0 = x102_inr_Foreach_kernelx102_inr_Foreach_concrete1_io_in_x84_a_0_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@4683.4]
  assign x86_ctrchain_clock = clock; // @[:@4466.4]
  assign x86_ctrchain_reset = reset; // @[:@4467.4]
  assign x86_ctrchain_io_input_reset = x102_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 130:103:@4623.4]
  assign x86_ctrchain_io_input_enable = x102_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 104:75:@4578.4 SpatialBlocks.scala 130:45:@4622.4]
  assign x102_inr_Foreach_sm_clock = clock; // @[:@4518.4]
  assign x102_inr_Foreach_sm_reset = reset; // @[:@4519.4]
  assign x102_inr_Foreach_sm_io_enable = _T_245 & _T_254; // @[SpatialBlocks.scala 112:18:@4605.4]
  assign x102_inr_Foreach_sm_io_ctrDone = io_rr ? _T_230 : 1'h0; // @[sm_RootController.scala 69:38:@4553.4]
  assign x102_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 114:21:@4607.4]
  assign x102_inr_Foreach_sm_io_backpressure = 1'h1; // @[SpatialBlocks.scala 105:24:@4579.4]
  assign x102_inr_Foreach_sm_io_break = 1'h0; // @[sm_RootController.scala 73:36:@4559.4]
  assign RetimeWrapper_clock = clock; // @[:@4546.4]
  assign RetimeWrapper_reset = reset; // @[:@4547.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@4549.4]
  assign RetimeWrapper_io_in = x86_ctrchain_io_output_done; // @[package.scala 94:16:@4548.4]
  assign RetimeWrapper_1_clock = clock; // @[:@4586.4]
  assign RetimeWrapper_1_reset = reset; // @[:@4587.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@4589.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@4588.4]
  assign RetimeWrapper_2_clock = clock; // @[:@4594.4]
  assign RetimeWrapper_2_reset = reset; // @[:@4595.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@4597.4]
  assign RetimeWrapper_2_io_in = x102_inr_Foreach_sm_io_done; // @[package.scala 94:16:@4596.4]
  assign x102_inr_Foreach_kernelx102_inr_Foreach_concrete1_clock = clock; // @[:@4625.4]
  assign x102_inr_Foreach_kernelx102_inr_Foreach_concrete1_reset = reset; // @[:@4626.4]
  assign x102_inr_Foreach_kernelx102_inr_Foreach_concrete1_io_sigsIn_done = x102_inr_Foreach_sm_io_done; // @[sm_x102_inr_Foreach.scala 101:22:@4712.4]
  assign x102_inr_Foreach_kernelx102_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_256 & _T_257; // @[sm_x102_inr_Foreach.scala 101:22:@4706.4]
  assign x102_inr_Foreach_kernelx102_inr_Foreach_concrete1_io_sigsIn_baseEn = _T_245 & _T_254; // @[sm_x102_inr_Foreach.scala 101:22:@4705.4]
  assign x102_inr_Foreach_kernelx102_inr_Foreach_concrete1_io_sigsIn_break = x102_inr_Foreach_sm_io_break; // @[sm_x102_inr_Foreach.scala 101:22:@4704.4]
  assign x102_inr_Foreach_kernelx102_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = x86_ctrchain_io_output_counts_0; // @[sm_x102_inr_Foreach.scala 101:22:@4699.4]
  assign x102_inr_Foreach_kernelx102_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x86_ctrchain_io_output_oobs_0; // @[sm_x102_inr_Foreach.scala 101:22:@4698.4]
  assign x102_inr_Foreach_kernelx102_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x102_inr_Foreach.scala 100:18:@4694.4]
  assign x119_outr_UnitPipe_sm_clock = clock; // @[:@4756.4]
  assign x119_outr_UnitPipe_sm_reset = reset; // @[:@4757.4]
  assign x119_outr_UnitPipe_sm_io_enable = _T_333 & _T_342; // @[SpatialBlocks.scala 112:18:@4827.4]
  assign x119_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 114:21:@4829.4]
  assign x119_outr_UnitPipe_sm_io_doneIn_0 = x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 102:67:@4799.4]
  assign x119_outr_UnitPipe_sm_io_ctrCopyDone_0 = x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 132:80:@4841.4]
  assign RetimeWrapper_3_clock = clock; // @[:@4808.4]
  assign RetimeWrapper_3_reset = reset; // @[:@4809.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@4811.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@4810.4]
  assign RetimeWrapper_4_clock = clock; // @[:@4816.4]
  assign RetimeWrapper_4_reset = reset; // @[:@4817.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@4819.4]
  assign RetimeWrapper_4_io_in = x119_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@4818.4]
  assign x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_clock = clock; // @[:@4843.4]
  assign x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_reset = reset; // @[:@4844.4]
  assign x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_x84_a_0_rPort_0_output_0 = x84_a_0_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@4910.4]
  assign x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_in_x82_TREADY = io_in_x82_TREADY; // @[sm_x119_outr_UnitPipe.scala 51:22:@4922.4]
  assign x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_sigsIn_done = x119_outr_UnitPipe_sm_io_done; // @[sm_x119_outr_UnitPipe.scala 87:22:@4950.4]
  assign x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_sigsIn_baseEn = _T_333 & _T_342; // @[sm_x119_outr_UnitPipe.scala 87:22:@4943.4]
  assign x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x119_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x119_outr_UnitPipe.scala 87:22:@4940.4]
  assign x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x119_outr_UnitPipe_sm_io_childAck_0; // @[sm_x119_outr_UnitPipe.scala 87:22:@4938.4]
  assign x119_outr_UnitPipe_kernelx119_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x119_outr_UnitPipe.scala 86:18:@4932.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_165 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_165 <= 1'h0;
    end else begin
      _T_165 <= _T_162;
    end
  end
endmodule
module AccelUnit( // @[:@4959.2]
  input          clock, // @[:@4960.4]
  input          reset, // @[:@4961.4]
  input          io_enable, // @[:@4962.4]
  output         io_done, // @[:@4962.4]
  input          io_reset, // @[:@4962.4]
  input          io_memStreams_loads_0_cmd_ready, // @[:@4962.4]
  output         io_memStreams_loads_0_cmd_valid, // @[:@4962.4]
  output [63:0]  io_memStreams_loads_0_cmd_bits_addr, // @[:@4962.4]
  output [31:0]  io_memStreams_loads_0_cmd_bits_size, // @[:@4962.4]
  output         io_memStreams_loads_0_data_ready, // @[:@4962.4]
  input          io_memStreams_loads_0_data_valid, // @[:@4962.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_0, // @[:@4962.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_1, // @[:@4962.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_2, // @[:@4962.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_3, // @[:@4962.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_4, // @[:@4962.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_5, // @[:@4962.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_6, // @[:@4962.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_7, // @[:@4962.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_8, // @[:@4962.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_9, // @[:@4962.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_10, // @[:@4962.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_11, // @[:@4962.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_12, // @[:@4962.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_13, // @[:@4962.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_14, // @[:@4962.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_15, // @[:@4962.4]
  input          io_memStreams_stores_0_cmd_ready, // @[:@4962.4]
  output         io_memStreams_stores_0_cmd_valid, // @[:@4962.4]
  output [63:0]  io_memStreams_stores_0_cmd_bits_addr, // @[:@4962.4]
  output [31:0]  io_memStreams_stores_0_cmd_bits_size, // @[:@4962.4]
  input          io_memStreams_stores_0_data_ready, // @[:@4962.4]
  output         io_memStreams_stores_0_data_valid, // @[:@4962.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_0, // @[:@4962.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_1, // @[:@4962.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_2, // @[:@4962.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_3, // @[:@4962.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_4, // @[:@4962.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_5, // @[:@4962.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_6, // @[:@4962.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_7, // @[:@4962.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_8, // @[:@4962.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_9, // @[:@4962.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_10, // @[:@4962.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_11, // @[:@4962.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_12, // @[:@4962.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_13, // @[:@4962.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_14, // @[:@4962.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_15, // @[:@4962.4]
  output [15:0]  io_memStreams_stores_0_data_bits_wstrb, // @[:@4962.4]
  output         io_memStreams_stores_0_wresp_ready, // @[:@4962.4]
  input          io_memStreams_stores_0_wresp_valid, // @[:@4962.4]
  input          io_memStreams_stores_0_wresp_bits, // @[:@4962.4]
  input          io_memStreams_gathers_0_cmd_ready, // @[:@4962.4]
  output         io_memStreams_gathers_0_cmd_valid, // @[:@4962.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_0, // @[:@4962.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_1, // @[:@4962.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_2, // @[:@4962.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_3, // @[:@4962.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_4, // @[:@4962.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_5, // @[:@4962.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_6, // @[:@4962.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_7, // @[:@4962.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_8, // @[:@4962.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_9, // @[:@4962.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_10, // @[:@4962.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_11, // @[:@4962.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_12, // @[:@4962.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_13, // @[:@4962.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_14, // @[:@4962.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_15, // @[:@4962.4]
  output         io_memStreams_gathers_0_data_ready, // @[:@4962.4]
  input          io_memStreams_gathers_0_data_valid, // @[:@4962.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_0, // @[:@4962.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_1, // @[:@4962.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_2, // @[:@4962.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_3, // @[:@4962.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_4, // @[:@4962.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_5, // @[:@4962.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_6, // @[:@4962.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_7, // @[:@4962.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_8, // @[:@4962.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_9, // @[:@4962.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_10, // @[:@4962.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_11, // @[:@4962.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_12, // @[:@4962.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_13, // @[:@4962.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_14, // @[:@4962.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_15, // @[:@4962.4]
  input          io_memStreams_scatters_0_cmd_ready, // @[:@4962.4]
  output         io_memStreams_scatters_0_cmd_valid, // @[:@4962.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_0, // @[:@4962.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_1, // @[:@4962.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_2, // @[:@4962.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_3, // @[:@4962.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_4, // @[:@4962.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_5, // @[:@4962.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_6, // @[:@4962.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_7, // @[:@4962.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_8, // @[:@4962.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_9, // @[:@4962.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_10, // @[:@4962.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_11, // @[:@4962.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_12, // @[:@4962.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_13, // @[:@4962.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_14, // @[:@4962.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_15, // @[:@4962.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_0, // @[:@4962.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_1, // @[:@4962.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_2, // @[:@4962.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_3, // @[:@4962.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_4, // @[:@4962.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_5, // @[:@4962.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_6, // @[:@4962.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_7, // @[:@4962.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_8, // @[:@4962.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_9, // @[:@4962.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_10, // @[:@4962.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_11, // @[:@4962.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_12, // @[:@4962.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_13, // @[:@4962.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_14, // @[:@4962.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_15, // @[:@4962.4]
  output         io_memStreams_scatters_0_wresp_ready, // @[:@4962.4]
  input          io_memStreams_scatters_0_wresp_valid, // @[:@4962.4]
  input          io_memStreams_scatters_0_wresp_bits, // @[:@4962.4]
  input          io_axiStreamsIn_0_TVALID, // @[:@4962.4]
  output         io_axiStreamsIn_0_TREADY, // @[:@4962.4]
  input  [255:0] io_axiStreamsIn_0_TDATA, // @[:@4962.4]
  input  [31:0]  io_axiStreamsIn_0_TSTRB, // @[:@4962.4]
  input  [31:0]  io_axiStreamsIn_0_TKEEP, // @[:@4962.4]
  input          io_axiStreamsIn_0_TLAST, // @[:@4962.4]
  input  [7:0]   io_axiStreamsIn_0_TID, // @[:@4962.4]
  input  [7:0]   io_axiStreamsIn_0_TDEST, // @[:@4962.4]
  input  [31:0]  io_axiStreamsIn_0_TUSER, // @[:@4962.4]
  output         io_axiStreamsOut_0_TVALID, // @[:@4962.4]
  input          io_axiStreamsOut_0_TREADY, // @[:@4962.4]
  output [511:0] io_axiStreamsOut_0_TDATA, // @[:@4962.4]
  output [63:0]  io_axiStreamsOut_0_TSTRB, // @[:@4962.4]
  output [63:0]  io_axiStreamsOut_0_TKEEP, // @[:@4962.4]
  output         io_axiStreamsOut_0_TLAST, // @[:@4962.4]
  output [7:0]   io_axiStreamsOut_0_TID, // @[:@4962.4]
  output [7:0]   io_axiStreamsOut_0_TDEST, // @[:@4962.4]
  output [31:0]  io_axiStreamsOut_0_TUSER, // @[:@4962.4]
  output         io_heap_0_req_valid, // @[:@4962.4]
  output         io_heap_0_req_bits_allocDealloc, // @[:@4962.4]
  output [63:0]  io_heap_0_req_bits_sizeAddr, // @[:@4962.4]
  input          io_heap_0_resp_valid, // @[:@4962.4]
  input          io_heap_0_resp_bits_allocDealloc, // @[:@4962.4]
  input  [63:0]  io_heap_0_resp_bits_sizeAddr, // @[:@4962.4]
  input  [63:0]  io_argIns_0, // @[:@4962.4]
  input          io_argOuts_0_port_ready, // @[:@4962.4]
  output         io_argOuts_0_port_valid, // @[:@4962.4]
  output [63:0]  io_argOuts_0_port_bits, // @[:@4962.4]
  input  [63:0]  io_argOuts_0_echo, // @[:@4962.4]
  input          io_argOuts_1_port_ready, // @[:@4962.4]
  output         io_argOuts_1_port_valid, // @[:@4962.4]
  output [63:0]  io_argOuts_1_port_bits, // @[:@4962.4]
  input  [63:0]  io_argOuts_1_echo, // @[:@4962.4]
  input          io_argOuts_2_port_ready, // @[:@4962.4]
  output         io_argOuts_2_port_valid, // @[:@4962.4]
  output [63:0]  io_argOuts_2_port_bits, // @[:@4962.4]
  input  [63:0]  io_argOuts_2_echo, // @[:@4962.4]
  input          io_argOuts_3_port_ready, // @[:@4962.4]
  output         io_argOuts_3_port_valid, // @[:@4962.4]
  output [63:0]  io_argOuts_3_port_bits, // @[:@4962.4]
  input  [63:0]  io_argOuts_3_echo, // @[:@4962.4]
  input          io_argOuts_4_port_ready, // @[:@4962.4]
  output         io_argOuts_4_port_valid, // @[:@4962.4]
  output [63:0]  io_argOuts_4_port_bits, // @[:@4962.4]
  input  [63:0]  io_argOuts_4_echo, // @[:@4962.4]
  input          io_argOuts_5_port_ready, // @[:@4962.4]
  output         io_argOuts_5_port_valid, // @[:@4962.4]
  output [63:0]  io_argOuts_5_port_bits, // @[:@4962.4]
  input  [63:0]  io_argOuts_5_echo, // @[:@4962.4]
  input          io_argOuts_6_port_ready, // @[:@4962.4]
  output         io_argOuts_6_port_valid, // @[:@4962.4]
  output [63:0]  io_argOuts_6_port_bits, // @[:@4962.4]
  input  [63:0]  io_argOuts_6_echo, // @[:@4962.4]
  input          io_argOuts_7_port_ready, // @[:@4962.4]
  output         io_argOuts_7_port_valid, // @[:@4962.4]
  output [63:0]  io_argOuts_7_port_bits, // @[:@4962.4]
  input  [63:0]  io_argOuts_7_echo, // @[:@4962.4]
  input          io_argOuts_8_port_ready, // @[:@4962.4]
  output         io_argOuts_8_port_valid, // @[:@4962.4]
  output [63:0]  io_argOuts_8_port_bits, // @[:@4962.4]
  input  [63:0]  io_argOuts_8_echo, // @[:@4962.4]
  input          io_argOuts_9_port_ready, // @[:@4962.4]
  output         io_argOuts_9_port_valid, // @[:@4962.4]
  output [63:0]  io_argOuts_9_port_bits, // @[:@4962.4]
  input  [63:0]  io_argOuts_9_echo // @[:@4962.4]
);
  wire  SingleCounter_clock; // @[Main.scala 28:32:@5156.4]
  wire  SingleCounter_reset; // @[Main.scala 28:32:@5156.4]
  wire  SingleCounter_io_input_reset; // @[Main.scala 28:32:@5156.4]
  wire  SingleCounter_io_output_done; // @[Main.scala 28:32:@5156.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@5174.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@5174.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@5174.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@5174.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@5174.4]
  wire  SRFF_clock; // @[Main.scala 33:28:@5187.4]
  wire  SRFF_reset; // @[Main.scala 33:28:@5187.4]
  wire  SRFF_io_input_set; // @[Main.scala 33:28:@5187.4]
  wire  SRFF_io_input_reset; // @[Main.scala 33:28:@5187.4]
  wire  SRFF_io_input_asyn_reset; // @[Main.scala 33:28:@5187.4]
  wire  SRFF_io_output; // @[Main.scala 33:28:@5187.4]
  wire  RootController_sm_clock; // @[sm_RootController.scala 32:18:@5230.4]
  wire  RootController_sm_reset; // @[sm_RootController.scala 32:18:@5230.4]
  wire  RootController_sm_io_enable; // @[sm_RootController.scala 32:18:@5230.4]
  wire  RootController_sm_io_done; // @[sm_RootController.scala 32:18:@5230.4]
  wire  RootController_sm_io_rst; // @[sm_RootController.scala 32:18:@5230.4]
  wire  RootController_sm_io_ctrDone; // @[sm_RootController.scala 32:18:@5230.4]
  wire  RootController_sm_io_ctrInc; // @[sm_RootController.scala 32:18:@5230.4]
  wire  RootController_sm_io_doneIn_0; // @[sm_RootController.scala 32:18:@5230.4]
  wire  RootController_sm_io_doneIn_1; // @[sm_RootController.scala 32:18:@5230.4]
  wire  RootController_sm_io_enableOut_0; // @[sm_RootController.scala 32:18:@5230.4]
  wire  RootController_sm_io_enableOut_1; // @[sm_RootController.scala 32:18:@5230.4]
  wire  RootController_sm_io_childAck_0; // @[sm_RootController.scala 32:18:@5230.4]
  wire  RootController_sm_io_childAck_1; // @[sm_RootController.scala 32:18:@5230.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@5267.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@5267.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@5267.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@5267.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@5267.4]
  wire  RootController_kernelRootController_concrete1_clock; // @[sm_RootController.scala 86:24:@5331.4]
  wire  RootController_kernelRootController_concrete1_reset; // @[sm_RootController.scala 86:24:@5331.4]
  wire  RootController_kernelRootController_concrete1_io_in_x82_TVALID; // @[sm_RootController.scala 86:24:@5331.4]
  wire  RootController_kernelRootController_concrete1_io_in_x82_TREADY; // @[sm_RootController.scala 86:24:@5331.4]
  wire [511:0] RootController_kernelRootController_concrete1_io_in_x82_TDATA; // @[sm_RootController.scala 86:24:@5331.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x82_TSTRB; // @[sm_RootController.scala 86:24:@5331.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x82_TKEEP; // @[sm_RootController.scala 86:24:@5331.4]
  wire  RootController_kernelRootController_concrete1_io_in_x82_TLAST; // @[sm_RootController.scala 86:24:@5331.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x82_TID; // @[sm_RootController.scala 86:24:@5331.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x82_TDEST; // @[sm_RootController.scala 86:24:@5331.4]
  wire [31:0] RootController_kernelRootController_concrete1_io_in_x82_TUSER; // @[sm_RootController.scala 86:24:@5331.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_0_cycs; // @[sm_RootController.scala 86:24:@5331.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_0_iters; // @[sm_RootController.scala 86:24:@5331.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_1_cycs; // @[sm_RootController.scala 86:24:@5331.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_1_iters; // @[sm_RootController.scala 86:24:@5331.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_2_cycs; // @[sm_RootController.scala 86:24:@5331.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_2_iters; // @[sm_RootController.scala 86:24:@5331.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_3_cycs; // @[sm_RootController.scala 86:24:@5331.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_3_iters; // @[sm_RootController.scala 86:24:@5331.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_3_stalls; // @[sm_RootController.scala 86:24:@5331.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_3_idles; // @[sm_RootController.scala 86:24:@5331.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_done; // @[sm_RootController.scala 86:24:@5331.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_baseEn; // @[sm_RootController.scala 86:24:@5331.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_RootController.scala 86:24:@5331.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_RootController.scala 86:24:@5331.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0; // @[sm_RootController.scala 86:24:@5331.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_1; // @[sm_RootController.scala 86:24:@5331.4]
  wire  RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[sm_RootController.scala 86:24:@5331.4]
  wire  RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_1; // @[sm_RootController.scala 86:24:@5331.4]
  wire  RootController_kernelRootController_concrete1_io_rr; // @[sm_RootController.scala 86:24:@5331.4]
  wire  _T_665; // @[package.scala 96:25:@5179.4 package.scala 96:25:@5180.4]
  wire  _T_738; // @[Main.scala 35:50:@5263.4]
  wire  _T_739; // @[Main.scala 35:59:@5264.4]
  wire  _T_751; // @[package.scala 100:49:@5284.4]
  reg  _T_754; // @[package.scala 48:56:@5285.4]
  reg [31:0] _RAND_0;
  SingleCounter SingleCounter ( // @[Main.scala 28:32:@5156.4]
    .clock(SingleCounter_clock),
    .reset(SingleCounter_reset),
    .io_input_reset(SingleCounter_io_input_reset),
    .io_output_done(SingleCounter_io_output_done)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@5174.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  SRFF SRFF ( // @[Main.scala 33:28:@5187.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  RootController_sm RootController_sm ( // @[sm_RootController.scala 32:18:@5230.4]
    .clock(RootController_sm_clock),
    .reset(RootController_sm_reset),
    .io_enable(RootController_sm_io_enable),
    .io_done(RootController_sm_io_done),
    .io_rst(RootController_sm_io_rst),
    .io_ctrDone(RootController_sm_io_ctrDone),
    .io_ctrInc(RootController_sm_io_ctrInc),
    .io_doneIn_0(RootController_sm_io_doneIn_0),
    .io_doneIn_1(RootController_sm_io_doneIn_1),
    .io_enableOut_0(RootController_sm_io_enableOut_0),
    .io_enableOut_1(RootController_sm_io_enableOut_1),
    .io_childAck_0(RootController_sm_io_childAck_0),
    .io_childAck_1(RootController_sm_io_childAck_1)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@5267.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RootController_kernelRootController_concrete1 RootController_kernelRootController_concrete1 ( // @[sm_RootController.scala 86:24:@5331.4]
    .clock(RootController_kernelRootController_concrete1_clock),
    .reset(RootController_kernelRootController_concrete1_reset),
    .io_in_x82_TVALID(RootController_kernelRootController_concrete1_io_in_x82_TVALID),
    .io_in_x82_TREADY(RootController_kernelRootController_concrete1_io_in_x82_TREADY),
    .io_in_x82_TDATA(RootController_kernelRootController_concrete1_io_in_x82_TDATA),
    .io_in_x82_TSTRB(RootController_kernelRootController_concrete1_io_in_x82_TSTRB),
    .io_in_x82_TKEEP(RootController_kernelRootController_concrete1_io_in_x82_TKEEP),
    .io_in_x82_TLAST(RootController_kernelRootController_concrete1_io_in_x82_TLAST),
    .io_in_x82_TID(RootController_kernelRootController_concrete1_io_in_x82_TID),
    .io_in_x82_TDEST(RootController_kernelRootController_concrete1_io_in_x82_TDEST),
    .io_in_x82_TUSER(RootController_kernelRootController_concrete1_io_in_x82_TUSER),
    .io_in_instrctrs_0_cycs(RootController_kernelRootController_concrete1_io_in_instrctrs_0_cycs),
    .io_in_instrctrs_0_iters(RootController_kernelRootController_concrete1_io_in_instrctrs_0_iters),
    .io_in_instrctrs_1_cycs(RootController_kernelRootController_concrete1_io_in_instrctrs_1_cycs),
    .io_in_instrctrs_1_iters(RootController_kernelRootController_concrete1_io_in_instrctrs_1_iters),
    .io_in_instrctrs_2_cycs(RootController_kernelRootController_concrete1_io_in_instrctrs_2_cycs),
    .io_in_instrctrs_2_iters(RootController_kernelRootController_concrete1_io_in_instrctrs_2_iters),
    .io_in_instrctrs_3_cycs(RootController_kernelRootController_concrete1_io_in_instrctrs_3_cycs),
    .io_in_instrctrs_3_iters(RootController_kernelRootController_concrete1_io_in_instrctrs_3_iters),
    .io_in_instrctrs_3_stalls(RootController_kernelRootController_concrete1_io_in_instrctrs_3_stalls),
    .io_in_instrctrs_3_idles(RootController_kernelRootController_concrete1_io_in_instrctrs_3_idles),
    .io_sigsIn_done(RootController_kernelRootController_concrete1_io_sigsIn_done),
    .io_sigsIn_baseEn(RootController_kernelRootController_concrete1_io_sigsIn_baseEn),
    .io_sigsIn_smEnableOuts_0(RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smChildAcks_0(RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsOut_smDoneIn_0(RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_1),
    .io_rr(RootController_kernelRootController_concrete1_io_rr)
  );
  assign _T_665 = RetimeWrapper_io_out; // @[package.scala 96:25:@5179.4 package.scala 96:25:@5180.4]
  assign _T_738 = io_enable & _T_665; // @[Main.scala 35:50:@5263.4]
  assign _T_739 = ~ SRFF_io_output; // @[Main.scala 35:59:@5264.4]
  assign _T_751 = RootController_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@5284.4]
  assign io_done = SRFF_io_output; // @[Main.scala 42:23:@5283.4]
  assign io_memStreams_loads_0_cmd_valid = 1'h0;
  assign io_memStreams_loads_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_loads_0_cmd_bits_size = 32'h0;
  assign io_memStreams_loads_0_data_ready = 1'h0;
  assign io_memStreams_stores_0_cmd_valid = 1'h0;
  assign io_memStreams_stores_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_stores_0_cmd_bits_size = 32'h0;
  assign io_memStreams_stores_0_data_valid = 1'h0;
  assign io_memStreams_stores_0_data_bits_wdata_0 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_1 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_2 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_3 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_4 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_5 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_6 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_7 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_8 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_9 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_10 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_11 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_12 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_13 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_14 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_15 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wstrb = 16'h0;
  assign io_memStreams_stores_0_wresp_ready = 1'h0;
  assign io_memStreams_gathers_0_cmd_valid = 1'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_0 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_1 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_2 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_3 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_4 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_5 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_6 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_7 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_8 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_9 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_10 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_11 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_12 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_13 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_14 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_15 = 64'h0;
  assign io_memStreams_gathers_0_data_ready = 1'h0;
  assign io_memStreams_scatters_0_cmd_valid = 1'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_0 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_1 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_2 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_3 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_4 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_5 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_6 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_7 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_8 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_9 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_10 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_11 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_12 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_13 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_14 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_15 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_0 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_1 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_2 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_3 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_4 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_5 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_6 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_7 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_8 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_9 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_10 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_11 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_12 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_13 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_14 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_15 = 32'h0;
  assign io_memStreams_scatters_0_wresp_ready = 1'h0;
  assign io_axiStreamsIn_0_TREADY = 1'h0;
  assign io_axiStreamsOut_0_TVALID = RootController_kernelRootController_concrete1_io_in_x82_TVALID; // @[sm_RootController.scala 47:22:@5399.4]
  assign io_axiStreamsOut_0_TDATA = RootController_kernelRootController_concrete1_io_in_x82_TDATA; // @[sm_RootController.scala 47:22:@5397.4]
  assign io_axiStreamsOut_0_TSTRB = RootController_kernelRootController_concrete1_io_in_x82_TSTRB; // @[sm_RootController.scala 47:22:@5396.4]
  assign io_axiStreamsOut_0_TKEEP = RootController_kernelRootController_concrete1_io_in_x82_TKEEP; // @[sm_RootController.scala 47:22:@5395.4]
  assign io_axiStreamsOut_0_TLAST = RootController_kernelRootController_concrete1_io_in_x82_TLAST; // @[sm_RootController.scala 47:22:@5394.4]
  assign io_axiStreamsOut_0_TID = RootController_kernelRootController_concrete1_io_in_x82_TID; // @[sm_RootController.scala 47:22:@5393.4]
  assign io_axiStreamsOut_0_TDEST = RootController_kernelRootController_concrete1_io_in_x82_TDEST; // @[sm_RootController.scala 47:22:@5392.4]
  assign io_axiStreamsOut_0_TUSER = RootController_kernelRootController_concrete1_io_in_x82_TUSER; // @[sm_RootController.scala 47:22:@5391.4]
  assign io_heap_0_req_valid = 1'h0;
  assign io_heap_0_req_bits_allocDealloc = 1'h0;
  assign io_heap_0_req_bits_sizeAddr = 64'h0;
  assign io_argOuts_0_port_valid = io_enable; // @[Instrument.scala 27:57:@5449.4]
  assign io_argOuts_0_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_0_cycs; // @[Instrument.scala 26:56:@5448.4]
  assign io_argOuts_1_port_valid = io_enable; // @[Instrument.scala 29:56:@5451.4]
  assign io_argOuts_1_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_0_iters; // @[Instrument.scala 28:55:@5450.4]
  assign io_argOuts_2_port_valid = io_enable; // @[Instrument.scala 31:58:@5453.4]
  assign io_argOuts_2_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_1_cycs; // @[Instrument.scala 30:57:@5452.4]
  assign io_argOuts_3_port_valid = io_enable; // @[Instrument.scala 33:57:@5455.4]
  assign io_argOuts_3_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_1_iters; // @[Instrument.scala 32:56:@5454.4]
  assign io_argOuts_4_port_valid = io_enable; // @[Instrument.scala 35:58:@5457.4]
  assign io_argOuts_4_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_2_cycs; // @[Instrument.scala 34:57:@5456.4]
  assign io_argOuts_5_port_valid = io_enable; // @[Instrument.scala 37:57:@5459.4]
  assign io_argOuts_5_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_2_iters; // @[Instrument.scala 36:56:@5458.4]
  assign io_argOuts_6_port_valid = io_enable; // @[Instrument.scala 39:58:@5461.4]
  assign io_argOuts_6_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_3_cycs; // @[Instrument.scala 38:57:@5460.4]
  assign io_argOuts_7_port_valid = io_enable; // @[Instrument.scala 41:57:@5463.4]
  assign io_argOuts_7_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_3_iters; // @[Instrument.scala 40:56:@5462.4]
  assign io_argOuts_8_port_valid = io_enable; // @[Instrument.scala 43:59:@5465.4]
  assign io_argOuts_8_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_3_stalls; // @[Instrument.scala 42:58:@5464.4]
  assign io_argOuts_9_port_valid = io_enable; // @[Instrument.scala 45:56:@5467.4]
  assign io_argOuts_9_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_3_idles; // @[Instrument.scala 44:55:@5466.4]
  assign SingleCounter_clock = clock; // @[:@5157.4]
  assign SingleCounter_reset = reset; // @[:@5158.4]
  assign SingleCounter_io_input_reset = reset; // @[Main.scala 29:79:@5172.4]
  assign RetimeWrapper_clock = clock; // @[:@5175.4]
  assign RetimeWrapper_reset = reset; // @[:@5176.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@5178.4]
  assign RetimeWrapper_io_in = SingleCounter_io_output_done; // @[package.scala 94:16:@5177.4]
  assign SRFF_clock = clock; // @[:@5188.4]
  assign SRFF_reset = reset; // @[:@5189.4]
  assign SRFF_io_input_set = RootController_sm_io_done; // @[Main.scala 51:29:@5447.4]
  assign SRFF_io_input_reset = RetimeWrapper_1_io_out; // @[Main.scala 40:31:@5281.4]
  assign SRFF_io_input_asyn_reset = RetimeWrapper_1_io_out; // @[Main.scala 41:36:@5282.4]
  assign RootController_sm_clock = clock; // @[:@5231.4]
  assign RootController_sm_reset = reset; // @[:@5232.4]
  assign RootController_sm_io_enable = _T_738 & _T_739; // @[Main.scala 39:33:@5280.4 SpatialBlocks.scala 112:18:@5319.4]
  assign RootController_sm_io_rst = RetimeWrapper_1_io_out; // @[SpatialBlocks.scala 106:15:@5313.4]
  assign RootController_sm_io_ctrDone = RootController_sm_io_ctrInc & _T_754; // @[Main.scala 43:34:@5288.4]
  assign RootController_sm_io_doneIn_0 = RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 102:67:@5308.4]
  assign RootController_sm_io_doneIn_1 = RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 102:67:@5309.4]
  assign RetimeWrapper_1_clock = clock; // @[:@5268.4]
  assign RetimeWrapper_1_reset = reset; // @[:@5269.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@5271.4]
  assign RetimeWrapper_1_io_in = reset | io_reset; // @[package.scala 94:16:@5270.4]
  assign RootController_kernelRootController_concrete1_clock = clock; // @[:@5332.4]
  assign RootController_kernelRootController_concrete1_reset = reset; // @[:@5333.4]
  assign RootController_kernelRootController_concrete1_io_in_x82_TREADY = io_axiStreamsOut_0_TREADY; // @[sm_RootController.scala 47:22:@5398.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_done = RootController_sm_io_done; // @[sm_RootController.scala 91:22:@5437.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_baseEn = _T_738 & _T_739; // @[sm_RootController.scala 91:22:@5430.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0 = RootController_sm_io_enableOut_0; // @[sm_RootController.scala 91:22:@5426.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_1 = RootController_sm_io_enableOut_1; // @[sm_RootController.scala 91:22:@5427.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0 = RootController_sm_io_childAck_0; // @[sm_RootController.scala 91:22:@5422.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_1 = RootController_sm_io_childAck_1; // @[sm_RootController.scala 91:22:@5423.4]
  assign RootController_kernelRootController_concrete1_io_rr = RetimeWrapper_io_out; // @[sm_RootController.scala 90:18:@5416.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_754 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_754 <= 1'h0;
    end else begin
      _T_754 <= _T_751;
    end
  end
endmodule
module DRAMHeap( // @[:@6374.2]
  input         io_accel_0_req_valid, // @[:@6377.4]
  input         io_accel_0_req_bits_allocDealloc, // @[:@6377.4]
  input  [63:0] io_accel_0_req_bits_sizeAddr, // @[:@6377.4]
  output        io_accel_0_resp_valid, // @[:@6377.4]
  output        io_accel_0_resp_bits_allocDealloc, // @[:@6377.4]
  output [63:0] io_accel_0_resp_bits_sizeAddr, // @[:@6377.4]
  output        io_host_0_req_valid, // @[:@6377.4]
  output        io_host_0_req_bits_allocDealloc, // @[:@6377.4]
  output [63:0] io_host_0_req_bits_sizeAddr, // @[:@6377.4]
  input         io_host_0_resp_valid, // @[:@6377.4]
  input         io_host_0_resp_bits_allocDealloc, // @[:@6377.4]
  input  [63:0] io_host_0_resp_bits_sizeAddr // @[:@6377.4]
);
  assign io_accel_0_resp_valid = io_host_0_resp_valid; // @[DRAMHeap.scala 24:18:@6384.4]
  assign io_accel_0_resp_bits_allocDealloc = io_host_0_resp_bits_allocDealloc; // @[DRAMHeap.scala 25:17:@6386.4]
  assign io_accel_0_resp_bits_sizeAddr = io_host_0_resp_bits_sizeAddr; // @[DRAMHeap.scala 25:17:@6385.4]
  assign io_host_0_req_valid = io_accel_0_req_valid; // @[DRAMHeap.scala 21:18:@6381.4]
  assign io_host_0_req_bits_allocDealloc = io_accel_0_req_bits_allocDealloc; // @[DRAMHeap.scala 21:18:@6380.4]
  assign io_host_0_req_bits_sizeAddr = io_accel_0_req_bits_sizeAddr; // @[DRAMHeap.scala 21:18:@6379.4]
endmodule
module RetimeWrapper_41( // @[:@6400.2]
  input         clock, // @[:@6401.4]
  input         reset, // @[:@6402.4]
  input         io_flow, // @[:@6403.4]
  input  [63:0] io_in, // @[:@6403.4]
  output [63:0] io_out // @[:@6403.4]
);
  wire [63:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@6405.4]
  wire [63:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@6405.4]
  wire [63:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@6405.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@6405.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@6405.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@6405.4]
  RetimeShiftRegister #(.WIDTH(64), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@6405.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@6418.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@6417.4]
  assign sr_init = 64'h0; // @[RetimeShiftRegister.scala 19:16:@6416.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@6415.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@6414.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@6412.4]
endmodule
module FringeFF( // @[:@6420.2]
  input         clock, // @[:@6421.4]
  input         reset, // @[:@6422.4]
  input  [63:0] io_in, // @[:@6423.4]
  input         io_reset, // @[:@6423.4]
  output [63:0] io_out, // @[:@6423.4]
  input         io_enable // @[:@6423.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@6426.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@6426.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@6426.4]
  wire [63:0] RetimeWrapper_io_in; // @[package.scala 93:22:@6426.4]
  wire [63:0] RetimeWrapper_io_out; // @[package.scala 93:22:@6426.4]
  wire [63:0] _T_18; // @[package.scala 96:25:@6431.4 package.scala 96:25:@6432.4]
  wire [63:0] _GEN_0; // @[FringeFF.scala 21:27:@6437.6]
  RetimeWrapper_41 RetimeWrapper ( // @[package.scala 93:22:@6426.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@6431.4 package.scala 96:25:@6432.4]
  assign _GEN_0 = io_reset ? 64'h0 : _T_18; // @[FringeFF.scala 21:27:@6437.6]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@6443.4]
  assign RetimeWrapper_clock = clock; // @[:@6427.4]
  assign RetimeWrapper_reset = reset; // @[:@6428.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@6430.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _GEN_0; // @[package.scala 94:16:@6429.4]
endmodule
module MuxN( // @[:@35572.2]
  input  [63:0] io_ins_0, // @[:@35575.4]
  input  [63:0] io_ins_1, // @[:@35575.4]
  input  [63:0] io_ins_2, // @[:@35575.4]
  input  [63:0] io_ins_3, // @[:@35575.4]
  input  [63:0] io_ins_4, // @[:@35575.4]
  input  [63:0] io_ins_5, // @[:@35575.4]
  input  [63:0] io_ins_6, // @[:@35575.4]
  input  [63:0] io_ins_7, // @[:@35575.4]
  input  [63:0] io_ins_8, // @[:@35575.4]
  input  [63:0] io_ins_9, // @[:@35575.4]
  input  [63:0] io_ins_10, // @[:@35575.4]
  input  [63:0] io_ins_11, // @[:@35575.4]
  input  [63:0] io_ins_12, // @[:@35575.4]
  input  [63:0] io_ins_13, // @[:@35575.4]
  input  [63:0] io_ins_14, // @[:@35575.4]
  input  [63:0] io_ins_15, // @[:@35575.4]
  input  [63:0] io_ins_16, // @[:@35575.4]
  input  [63:0] io_ins_17, // @[:@35575.4]
  input  [63:0] io_ins_18, // @[:@35575.4]
  input  [63:0] io_ins_19, // @[:@35575.4]
  input  [63:0] io_ins_20, // @[:@35575.4]
  input  [63:0] io_ins_21, // @[:@35575.4]
  input  [63:0] io_ins_22, // @[:@35575.4]
  input  [63:0] io_ins_23, // @[:@35575.4]
  input  [63:0] io_ins_24, // @[:@35575.4]
  input  [63:0] io_ins_25, // @[:@35575.4]
  input  [63:0] io_ins_26, // @[:@35575.4]
  input  [63:0] io_ins_27, // @[:@35575.4]
  input  [63:0] io_ins_28, // @[:@35575.4]
  input  [63:0] io_ins_29, // @[:@35575.4]
  input  [63:0] io_ins_30, // @[:@35575.4]
  input  [63:0] io_ins_31, // @[:@35575.4]
  input  [63:0] io_ins_32, // @[:@35575.4]
  input  [63:0] io_ins_33, // @[:@35575.4]
  input  [63:0] io_ins_34, // @[:@35575.4]
  input  [63:0] io_ins_35, // @[:@35575.4]
  input  [63:0] io_ins_36, // @[:@35575.4]
  input  [63:0] io_ins_37, // @[:@35575.4]
  input  [63:0] io_ins_38, // @[:@35575.4]
  input  [63:0] io_ins_39, // @[:@35575.4]
  input  [63:0] io_ins_40, // @[:@35575.4]
  input  [63:0] io_ins_41, // @[:@35575.4]
  input  [63:0] io_ins_42, // @[:@35575.4]
  input  [63:0] io_ins_43, // @[:@35575.4]
  input  [63:0] io_ins_44, // @[:@35575.4]
  input  [63:0] io_ins_45, // @[:@35575.4]
  input  [63:0] io_ins_46, // @[:@35575.4]
  input  [63:0] io_ins_47, // @[:@35575.4]
  input  [63:0] io_ins_48, // @[:@35575.4]
  input  [63:0] io_ins_49, // @[:@35575.4]
  input  [63:0] io_ins_50, // @[:@35575.4]
  input  [63:0] io_ins_51, // @[:@35575.4]
  input  [63:0] io_ins_52, // @[:@35575.4]
  input  [63:0] io_ins_53, // @[:@35575.4]
  input  [63:0] io_ins_54, // @[:@35575.4]
  input  [63:0] io_ins_55, // @[:@35575.4]
  input  [63:0] io_ins_56, // @[:@35575.4]
  input  [63:0] io_ins_57, // @[:@35575.4]
  input  [63:0] io_ins_58, // @[:@35575.4]
  input  [63:0] io_ins_59, // @[:@35575.4]
  input  [63:0] io_ins_60, // @[:@35575.4]
  input  [63:0] io_ins_61, // @[:@35575.4]
  input  [63:0] io_ins_62, // @[:@35575.4]
  input  [63:0] io_ins_63, // @[:@35575.4]
  input  [63:0] io_ins_64, // @[:@35575.4]
  input  [63:0] io_ins_65, // @[:@35575.4]
  input  [63:0] io_ins_66, // @[:@35575.4]
  input  [63:0] io_ins_67, // @[:@35575.4]
  input  [63:0] io_ins_68, // @[:@35575.4]
  input  [63:0] io_ins_69, // @[:@35575.4]
  input  [63:0] io_ins_70, // @[:@35575.4]
  input  [63:0] io_ins_71, // @[:@35575.4]
  input  [63:0] io_ins_72, // @[:@35575.4]
  input  [63:0] io_ins_73, // @[:@35575.4]
  input  [63:0] io_ins_74, // @[:@35575.4]
  input  [63:0] io_ins_75, // @[:@35575.4]
  input  [63:0] io_ins_76, // @[:@35575.4]
  input  [63:0] io_ins_77, // @[:@35575.4]
  input  [63:0] io_ins_78, // @[:@35575.4]
  input  [63:0] io_ins_79, // @[:@35575.4]
  input  [63:0] io_ins_80, // @[:@35575.4]
  input  [63:0] io_ins_81, // @[:@35575.4]
  input  [63:0] io_ins_82, // @[:@35575.4]
  input  [63:0] io_ins_83, // @[:@35575.4]
  input  [63:0] io_ins_84, // @[:@35575.4]
  input  [63:0] io_ins_85, // @[:@35575.4]
  input  [63:0] io_ins_86, // @[:@35575.4]
  input  [63:0] io_ins_87, // @[:@35575.4]
  input  [63:0] io_ins_88, // @[:@35575.4]
  input  [63:0] io_ins_89, // @[:@35575.4]
  input  [63:0] io_ins_90, // @[:@35575.4]
  input  [63:0] io_ins_91, // @[:@35575.4]
  input  [63:0] io_ins_92, // @[:@35575.4]
  input  [63:0] io_ins_93, // @[:@35575.4]
  input  [63:0] io_ins_94, // @[:@35575.4]
  input  [63:0] io_ins_95, // @[:@35575.4]
  input  [63:0] io_ins_96, // @[:@35575.4]
  input  [63:0] io_ins_97, // @[:@35575.4]
  input  [63:0] io_ins_98, // @[:@35575.4]
  input  [63:0] io_ins_99, // @[:@35575.4]
  input  [63:0] io_ins_100, // @[:@35575.4]
  input  [63:0] io_ins_101, // @[:@35575.4]
  input  [63:0] io_ins_102, // @[:@35575.4]
  input  [63:0] io_ins_103, // @[:@35575.4]
  input  [63:0] io_ins_104, // @[:@35575.4]
  input  [63:0] io_ins_105, // @[:@35575.4]
  input  [63:0] io_ins_106, // @[:@35575.4]
  input  [63:0] io_ins_107, // @[:@35575.4]
  input  [63:0] io_ins_108, // @[:@35575.4]
  input  [63:0] io_ins_109, // @[:@35575.4]
  input  [63:0] io_ins_110, // @[:@35575.4]
  input  [63:0] io_ins_111, // @[:@35575.4]
  input  [63:0] io_ins_112, // @[:@35575.4]
  input  [63:0] io_ins_113, // @[:@35575.4]
  input  [63:0] io_ins_114, // @[:@35575.4]
  input  [63:0] io_ins_115, // @[:@35575.4]
  input  [63:0] io_ins_116, // @[:@35575.4]
  input  [63:0] io_ins_117, // @[:@35575.4]
  input  [63:0] io_ins_118, // @[:@35575.4]
  input  [63:0] io_ins_119, // @[:@35575.4]
  input  [63:0] io_ins_120, // @[:@35575.4]
  input  [63:0] io_ins_121, // @[:@35575.4]
  input  [63:0] io_ins_122, // @[:@35575.4]
  input  [63:0] io_ins_123, // @[:@35575.4]
  input  [63:0] io_ins_124, // @[:@35575.4]
  input  [63:0] io_ins_125, // @[:@35575.4]
  input  [63:0] io_ins_126, // @[:@35575.4]
  input  [63:0] io_ins_127, // @[:@35575.4]
  input  [63:0] io_ins_128, // @[:@35575.4]
  input  [63:0] io_ins_129, // @[:@35575.4]
  input  [63:0] io_ins_130, // @[:@35575.4]
  input  [63:0] io_ins_131, // @[:@35575.4]
  input  [63:0] io_ins_132, // @[:@35575.4]
  input  [63:0] io_ins_133, // @[:@35575.4]
  input  [63:0] io_ins_134, // @[:@35575.4]
  input  [63:0] io_ins_135, // @[:@35575.4]
  input  [63:0] io_ins_136, // @[:@35575.4]
  input  [63:0] io_ins_137, // @[:@35575.4]
  input  [63:0] io_ins_138, // @[:@35575.4]
  input  [63:0] io_ins_139, // @[:@35575.4]
  input  [63:0] io_ins_140, // @[:@35575.4]
  input  [63:0] io_ins_141, // @[:@35575.4]
  input  [63:0] io_ins_142, // @[:@35575.4]
  input  [63:0] io_ins_143, // @[:@35575.4]
  input  [63:0] io_ins_144, // @[:@35575.4]
  input  [63:0] io_ins_145, // @[:@35575.4]
  input  [63:0] io_ins_146, // @[:@35575.4]
  input  [63:0] io_ins_147, // @[:@35575.4]
  input  [63:0] io_ins_148, // @[:@35575.4]
  input  [63:0] io_ins_149, // @[:@35575.4]
  input  [63:0] io_ins_150, // @[:@35575.4]
  input  [63:0] io_ins_151, // @[:@35575.4]
  input  [63:0] io_ins_152, // @[:@35575.4]
  input  [63:0] io_ins_153, // @[:@35575.4]
  input  [63:0] io_ins_154, // @[:@35575.4]
  input  [63:0] io_ins_155, // @[:@35575.4]
  input  [63:0] io_ins_156, // @[:@35575.4]
  input  [63:0] io_ins_157, // @[:@35575.4]
  input  [63:0] io_ins_158, // @[:@35575.4]
  input  [63:0] io_ins_159, // @[:@35575.4]
  input  [63:0] io_ins_160, // @[:@35575.4]
  input  [63:0] io_ins_161, // @[:@35575.4]
  input  [63:0] io_ins_162, // @[:@35575.4]
  input  [63:0] io_ins_163, // @[:@35575.4]
  input  [63:0] io_ins_164, // @[:@35575.4]
  input  [63:0] io_ins_165, // @[:@35575.4]
  input  [63:0] io_ins_166, // @[:@35575.4]
  input  [63:0] io_ins_167, // @[:@35575.4]
  input  [63:0] io_ins_168, // @[:@35575.4]
  input  [63:0] io_ins_169, // @[:@35575.4]
  input  [63:0] io_ins_170, // @[:@35575.4]
  input  [63:0] io_ins_171, // @[:@35575.4]
  input  [63:0] io_ins_172, // @[:@35575.4]
  input  [63:0] io_ins_173, // @[:@35575.4]
  input  [63:0] io_ins_174, // @[:@35575.4]
  input  [63:0] io_ins_175, // @[:@35575.4]
  input  [63:0] io_ins_176, // @[:@35575.4]
  input  [63:0] io_ins_177, // @[:@35575.4]
  input  [63:0] io_ins_178, // @[:@35575.4]
  input  [63:0] io_ins_179, // @[:@35575.4]
  input  [63:0] io_ins_180, // @[:@35575.4]
  input  [63:0] io_ins_181, // @[:@35575.4]
  input  [63:0] io_ins_182, // @[:@35575.4]
  input  [63:0] io_ins_183, // @[:@35575.4]
  input  [63:0] io_ins_184, // @[:@35575.4]
  input  [63:0] io_ins_185, // @[:@35575.4]
  input  [63:0] io_ins_186, // @[:@35575.4]
  input  [63:0] io_ins_187, // @[:@35575.4]
  input  [63:0] io_ins_188, // @[:@35575.4]
  input  [63:0] io_ins_189, // @[:@35575.4]
  input  [63:0] io_ins_190, // @[:@35575.4]
  input  [63:0] io_ins_191, // @[:@35575.4]
  input  [63:0] io_ins_192, // @[:@35575.4]
  input  [63:0] io_ins_193, // @[:@35575.4]
  input  [63:0] io_ins_194, // @[:@35575.4]
  input  [63:0] io_ins_195, // @[:@35575.4]
  input  [63:0] io_ins_196, // @[:@35575.4]
  input  [63:0] io_ins_197, // @[:@35575.4]
  input  [63:0] io_ins_198, // @[:@35575.4]
  input  [63:0] io_ins_199, // @[:@35575.4]
  input  [63:0] io_ins_200, // @[:@35575.4]
  input  [63:0] io_ins_201, // @[:@35575.4]
  input  [63:0] io_ins_202, // @[:@35575.4]
  input  [63:0] io_ins_203, // @[:@35575.4]
  input  [63:0] io_ins_204, // @[:@35575.4]
  input  [63:0] io_ins_205, // @[:@35575.4]
  input  [63:0] io_ins_206, // @[:@35575.4]
  input  [63:0] io_ins_207, // @[:@35575.4]
  input  [63:0] io_ins_208, // @[:@35575.4]
  input  [63:0] io_ins_209, // @[:@35575.4]
  input  [63:0] io_ins_210, // @[:@35575.4]
  input  [63:0] io_ins_211, // @[:@35575.4]
  input  [63:0] io_ins_212, // @[:@35575.4]
  input  [63:0] io_ins_213, // @[:@35575.4]
  input  [63:0] io_ins_214, // @[:@35575.4]
  input  [63:0] io_ins_215, // @[:@35575.4]
  input  [63:0] io_ins_216, // @[:@35575.4]
  input  [63:0] io_ins_217, // @[:@35575.4]
  input  [63:0] io_ins_218, // @[:@35575.4]
  input  [63:0] io_ins_219, // @[:@35575.4]
  input  [63:0] io_ins_220, // @[:@35575.4]
  input  [63:0] io_ins_221, // @[:@35575.4]
  input  [63:0] io_ins_222, // @[:@35575.4]
  input  [63:0] io_ins_223, // @[:@35575.4]
  input  [63:0] io_ins_224, // @[:@35575.4]
  input  [63:0] io_ins_225, // @[:@35575.4]
  input  [63:0] io_ins_226, // @[:@35575.4]
  input  [63:0] io_ins_227, // @[:@35575.4]
  input  [63:0] io_ins_228, // @[:@35575.4]
  input  [63:0] io_ins_229, // @[:@35575.4]
  input  [63:0] io_ins_230, // @[:@35575.4]
  input  [63:0] io_ins_231, // @[:@35575.4]
  input  [63:0] io_ins_232, // @[:@35575.4]
  input  [63:0] io_ins_233, // @[:@35575.4]
  input  [63:0] io_ins_234, // @[:@35575.4]
  input  [63:0] io_ins_235, // @[:@35575.4]
  input  [63:0] io_ins_236, // @[:@35575.4]
  input  [63:0] io_ins_237, // @[:@35575.4]
  input  [63:0] io_ins_238, // @[:@35575.4]
  input  [63:0] io_ins_239, // @[:@35575.4]
  input  [63:0] io_ins_240, // @[:@35575.4]
  input  [63:0] io_ins_241, // @[:@35575.4]
  input  [63:0] io_ins_242, // @[:@35575.4]
  input  [63:0] io_ins_243, // @[:@35575.4]
  input  [63:0] io_ins_244, // @[:@35575.4]
  input  [63:0] io_ins_245, // @[:@35575.4]
  input  [63:0] io_ins_246, // @[:@35575.4]
  input  [63:0] io_ins_247, // @[:@35575.4]
  input  [63:0] io_ins_248, // @[:@35575.4]
  input  [63:0] io_ins_249, // @[:@35575.4]
  input  [63:0] io_ins_250, // @[:@35575.4]
  input  [63:0] io_ins_251, // @[:@35575.4]
  input  [63:0] io_ins_252, // @[:@35575.4]
  input  [63:0] io_ins_253, // @[:@35575.4]
  input  [63:0] io_ins_254, // @[:@35575.4]
  input  [63:0] io_ins_255, // @[:@35575.4]
  input  [63:0] io_ins_256, // @[:@35575.4]
  input  [63:0] io_ins_257, // @[:@35575.4]
  input  [63:0] io_ins_258, // @[:@35575.4]
  input  [63:0] io_ins_259, // @[:@35575.4]
  input  [63:0] io_ins_260, // @[:@35575.4]
  input  [63:0] io_ins_261, // @[:@35575.4]
  input  [63:0] io_ins_262, // @[:@35575.4]
  input  [63:0] io_ins_263, // @[:@35575.4]
  input  [63:0] io_ins_264, // @[:@35575.4]
  input  [63:0] io_ins_265, // @[:@35575.4]
  input  [63:0] io_ins_266, // @[:@35575.4]
  input  [63:0] io_ins_267, // @[:@35575.4]
  input  [63:0] io_ins_268, // @[:@35575.4]
  input  [63:0] io_ins_269, // @[:@35575.4]
  input  [63:0] io_ins_270, // @[:@35575.4]
  input  [63:0] io_ins_271, // @[:@35575.4]
  input  [63:0] io_ins_272, // @[:@35575.4]
  input  [63:0] io_ins_273, // @[:@35575.4]
  input  [63:0] io_ins_274, // @[:@35575.4]
  input  [63:0] io_ins_275, // @[:@35575.4]
  input  [63:0] io_ins_276, // @[:@35575.4]
  input  [63:0] io_ins_277, // @[:@35575.4]
  input  [63:0] io_ins_278, // @[:@35575.4]
  input  [63:0] io_ins_279, // @[:@35575.4]
  input  [63:0] io_ins_280, // @[:@35575.4]
  input  [63:0] io_ins_281, // @[:@35575.4]
  input  [63:0] io_ins_282, // @[:@35575.4]
  input  [63:0] io_ins_283, // @[:@35575.4]
  input  [63:0] io_ins_284, // @[:@35575.4]
  input  [63:0] io_ins_285, // @[:@35575.4]
  input  [63:0] io_ins_286, // @[:@35575.4]
  input  [63:0] io_ins_287, // @[:@35575.4]
  input  [63:0] io_ins_288, // @[:@35575.4]
  input  [63:0] io_ins_289, // @[:@35575.4]
  input  [63:0] io_ins_290, // @[:@35575.4]
  input  [63:0] io_ins_291, // @[:@35575.4]
  input  [63:0] io_ins_292, // @[:@35575.4]
  input  [63:0] io_ins_293, // @[:@35575.4]
  input  [63:0] io_ins_294, // @[:@35575.4]
  input  [63:0] io_ins_295, // @[:@35575.4]
  input  [63:0] io_ins_296, // @[:@35575.4]
  input  [63:0] io_ins_297, // @[:@35575.4]
  input  [63:0] io_ins_298, // @[:@35575.4]
  input  [63:0] io_ins_299, // @[:@35575.4]
  input  [63:0] io_ins_300, // @[:@35575.4]
  input  [63:0] io_ins_301, // @[:@35575.4]
  input  [63:0] io_ins_302, // @[:@35575.4]
  input  [63:0] io_ins_303, // @[:@35575.4]
  input  [63:0] io_ins_304, // @[:@35575.4]
  input  [63:0] io_ins_305, // @[:@35575.4]
  input  [63:0] io_ins_306, // @[:@35575.4]
  input  [63:0] io_ins_307, // @[:@35575.4]
  input  [63:0] io_ins_308, // @[:@35575.4]
  input  [63:0] io_ins_309, // @[:@35575.4]
  input  [63:0] io_ins_310, // @[:@35575.4]
  input  [63:0] io_ins_311, // @[:@35575.4]
  input  [63:0] io_ins_312, // @[:@35575.4]
  input  [63:0] io_ins_313, // @[:@35575.4]
  input  [63:0] io_ins_314, // @[:@35575.4]
  input  [63:0] io_ins_315, // @[:@35575.4]
  input  [63:0] io_ins_316, // @[:@35575.4]
  input  [63:0] io_ins_317, // @[:@35575.4]
  input  [63:0] io_ins_318, // @[:@35575.4]
  input  [63:0] io_ins_319, // @[:@35575.4]
  input  [63:0] io_ins_320, // @[:@35575.4]
  input  [63:0] io_ins_321, // @[:@35575.4]
  input  [63:0] io_ins_322, // @[:@35575.4]
  input  [63:0] io_ins_323, // @[:@35575.4]
  input  [63:0] io_ins_324, // @[:@35575.4]
  input  [63:0] io_ins_325, // @[:@35575.4]
  input  [63:0] io_ins_326, // @[:@35575.4]
  input  [63:0] io_ins_327, // @[:@35575.4]
  input  [63:0] io_ins_328, // @[:@35575.4]
  input  [63:0] io_ins_329, // @[:@35575.4]
  input  [63:0] io_ins_330, // @[:@35575.4]
  input  [63:0] io_ins_331, // @[:@35575.4]
  input  [63:0] io_ins_332, // @[:@35575.4]
  input  [63:0] io_ins_333, // @[:@35575.4]
  input  [63:0] io_ins_334, // @[:@35575.4]
  input  [63:0] io_ins_335, // @[:@35575.4]
  input  [63:0] io_ins_336, // @[:@35575.4]
  input  [63:0] io_ins_337, // @[:@35575.4]
  input  [63:0] io_ins_338, // @[:@35575.4]
  input  [63:0] io_ins_339, // @[:@35575.4]
  input  [63:0] io_ins_340, // @[:@35575.4]
  input  [63:0] io_ins_341, // @[:@35575.4]
  input  [63:0] io_ins_342, // @[:@35575.4]
  input  [63:0] io_ins_343, // @[:@35575.4]
  input  [63:0] io_ins_344, // @[:@35575.4]
  input  [63:0] io_ins_345, // @[:@35575.4]
  input  [63:0] io_ins_346, // @[:@35575.4]
  input  [63:0] io_ins_347, // @[:@35575.4]
  input  [63:0] io_ins_348, // @[:@35575.4]
  input  [63:0] io_ins_349, // @[:@35575.4]
  input  [63:0] io_ins_350, // @[:@35575.4]
  input  [63:0] io_ins_351, // @[:@35575.4]
  input  [63:0] io_ins_352, // @[:@35575.4]
  input  [63:0] io_ins_353, // @[:@35575.4]
  input  [63:0] io_ins_354, // @[:@35575.4]
  input  [63:0] io_ins_355, // @[:@35575.4]
  input  [63:0] io_ins_356, // @[:@35575.4]
  input  [63:0] io_ins_357, // @[:@35575.4]
  input  [63:0] io_ins_358, // @[:@35575.4]
  input  [63:0] io_ins_359, // @[:@35575.4]
  input  [63:0] io_ins_360, // @[:@35575.4]
  input  [63:0] io_ins_361, // @[:@35575.4]
  input  [63:0] io_ins_362, // @[:@35575.4]
  input  [63:0] io_ins_363, // @[:@35575.4]
  input  [63:0] io_ins_364, // @[:@35575.4]
  input  [63:0] io_ins_365, // @[:@35575.4]
  input  [63:0] io_ins_366, // @[:@35575.4]
  input  [63:0] io_ins_367, // @[:@35575.4]
  input  [63:0] io_ins_368, // @[:@35575.4]
  input  [63:0] io_ins_369, // @[:@35575.4]
  input  [63:0] io_ins_370, // @[:@35575.4]
  input  [63:0] io_ins_371, // @[:@35575.4]
  input  [63:0] io_ins_372, // @[:@35575.4]
  input  [63:0] io_ins_373, // @[:@35575.4]
  input  [63:0] io_ins_374, // @[:@35575.4]
  input  [63:0] io_ins_375, // @[:@35575.4]
  input  [63:0] io_ins_376, // @[:@35575.4]
  input  [63:0] io_ins_377, // @[:@35575.4]
  input  [63:0] io_ins_378, // @[:@35575.4]
  input  [63:0] io_ins_379, // @[:@35575.4]
  input  [63:0] io_ins_380, // @[:@35575.4]
  input  [63:0] io_ins_381, // @[:@35575.4]
  input  [63:0] io_ins_382, // @[:@35575.4]
  input  [63:0] io_ins_383, // @[:@35575.4]
  input  [63:0] io_ins_384, // @[:@35575.4]
  input  [63:0] io_ins_385, // @[:@35575.4]
  input  [63:0] io_ins_386, // @[:@35575.4]
  input  [63:0] io_ins_387, // @[:@35575.4]
  input  [63:0] io_ins_388, // @[:@35575.4]
  input  [63:0] io_ins_389, // @[:@35575.4]
  input  [63:0] io_ins_390, // @[:@35575.4]
  input  [63:0] io_ins_391, // @[:@35575.4]
  input  [63:0] io_ins_392, // @[:@35575.4]
  input  [63:0] io_ins_393, // @[:@35575.4]
  input  [63:0] io_ins_394, // @[:@35575.4]
  input  [63:0] io_ins_395, // @[:@35575.4]
  input  [63:0] io_ins_396, // @[:@35575.4]
  input  [63:0] io_ins_397, // @[:@35575.4]
  input  [63:0] io_ins_398, // @[:@35575.4]
  input  [63:0] io_ins_399, // @[:@35575.4]
  input  [63:0] io_ins_400, // @[:@35575.4]
  input  [63:0] io_ins_401, // @[:@35575.4]
  input  [63:0] io_ins_402, // @[:@35575.4]
  input  [63:0] io_ins_403, // @[:@35575.4]
  input  [63:0] io_ins_404, // @[:@35575.4]
  input  [63:0] io_ins_405, // @[:@35575.4]
  input  [63:0] io_ins_406, // @[:@35575.4]
  input  [63:0] io_ins_407, // @[:@35575.4]
  input  [63:0] io_ins_408, // @[:@35575.4]
  input  [63:0] io_ins_409, // @[:@35575.4]
  input  [63:0] io_ins_410, // @[:@35575.4]
  input  [63:0] io_ins_411, // @[:@35575.4]
  input  [63:0] io_ins_412, // @[:@35575.4]
  input  [63:0] io_ins_413, // @[:@35575.4]
  input  [63:0] io_ins_414, // @[:@35575.4]
  input  [63:0] io_ins_415, // @[:@35575.4]
  input  [63:0] io_ins_416, // @[:@35575.4]
  input  [63:0] io_ins_417, // @[:@35575.4]
  input  [63:0] io_ins_418, // @[:@35575.4]
  input  [63:0] io_ins_419, // @[:@35575.4]
  input  [63:0] io_ins_420, // @[:@35575.4]
  input  [63:0] io_ins_421, // @[:@35575.4]
  input  [63:0] io_ins_422, // @[:@35575.4]
  input  [63:0] io_ins_423, // @[:@35575.4]
  input  [63:0] io_ins_424, // @[:@35575.4]
  input  [63:0] io_ins_425, // @[:@35575.4]
  input  [63:0] io_ins_426, // @[:@35575.4]
  input  [63:0] io_ins_427, // @[:@35575.4]
  input  [63:0] io_ins_428, // @[:@35575.4]
  input  [63:0] io_ins_429, // @[:@35575.4]
  input  [63:0] io_ins_430, // @[:@35575.4]
  input  [63:0] io_ins_431, // @[:@35575.4]
  input  [63:0] io_ins_432, // @[:@35575.4]
  input  [63:0] io_ins_433, // @[:@35575.4]
  input  [63:0] io_ins_434, // @[:@35575.4]
  input  [63:0] io_ins_435, // @[:@35575.4]
  input  [63:0] io_ins_436, // @[:@35575.4]
  input  [63:0] io_ins_437, // @[:@35575.4]
  input  [63:0] io_ins_438, // @[:@35575.4]
  input  [63:0] io_ins_439, // @[:@35575.4]
  input  [63:0] io_ins_440, // @[:@35575.4]
  input  [63:0] io_ins_441, // @[:@35575.4]
  input  [63:0] io_ins_442, // @[:@35575.4]
  input  [63:0] io_ins_443, // @[:@35575.4]
  input  [63:0] io_ins_444, // @[:@35575.4]
  input  [63:0] io_ins_445, // @[:@35575.4]
  input  [63:0] io_ins_446, // @[:@35575.4]
  input  [63:0] io_ins_447, // @[:@35575.4]
  input  [63:0] io_ins_448, // @[:@35575.4]
  input  [63:0] io_ins_449, // @[:@35575.4]
  input  [63:0] io_ins_450, // @[:@35575.4]
  input  [63:0] io_ins_451, // @[:@35575.4]
  input  [63:0] io_ins_452, // @[:@35575.4]
  input  [63:0] io_ins_453, // @[:@35575.4]
  input  [63:0] io_ins_454, // @[:@35575.4]
  input  [63:0] io_ins_455, // @[:@35575.4]
  input  [63:0] io_ins_456, // @[:@35575.4]
  input  [63:0] io_ins_457, // @[:@35575.4]
  input  [63:0] io_ins_458, // @[:@35575.4]
  input  [63:0] io_ins_459, // @[:@35575.4]
  input  [63:0] io_ins_460, // @[:@35575.4]
  input  [63:0] io_ins_461, // @[:@35575.4]
  input  [63:0] io_ins_462, // @[:@35575.4]
  input  [63:0] io_ins_463, // @[:@35575.4]
  input  [63:0] io_ins_464, // @[:@35575.4]
  input  [63:0] io_ins_465, // @[:@35575.4]
  input  [63:0] io_ins_466, // @[:@35575.4]
  input  [63:0] io_ins_467, // @[:@35575.4]
  input  [63:0] io_ins_468, // @[:@35575.4]
  input  [63:0] io_ins_469, // @[:@35575.4]
  input  [63:0] io_ins_470, // @[:@35575.4]
  input  [63:0] io_ins_471, // @[:@35575.4]
  input  [63:0] io_ins_472, // @[:@35575.4]
  input  [63:0] io_ins_473, // @[:@35575.4]
  input  [63:0] io_ins_474, // @[:@35575.4]
  input  [63:0] io_ins_475, // @[:@35575.4]
  input  [63:0] io_ins_476, // @[:@35575.4]
  input  [63:0] io_ins_477, // @[:@35575.4]
  input  [63:0] io_ins_478, // @[:@35575.4]
  input  [63:0] io_ins_479, // @[:@35575.4]
  input  [63:0] io_ins_480, // @[:@35575.4]
  input  [63:0] io_ins_481, // @[:@35575.4]
  input  [63:0] io_ins_482, // @[:@35575.4]
  input  [63:0] io_ins_483, // @[:@35575.4]
  input  [63:0] io_ins_484, // @[:@35575.4]
  input  [63:0] io_ins_485, // @[:@35575.4]
  input  [63:0] io_ins_486, // @[:@35575.4]
  input  [63:0] io_ins_487, // @[:@35575.4]
  input  [63:0] io_ins_488, // @[:@35575.4]
  input  [63:0] io_ins_489, // @[:@35575.4]
  input  [63:0] io_ins_490, // @[:@35575.4]
  input  [63:0] io_ins_491, // @[:@35575.4]
  input  [63:0] io_ins_492, // @[:@35575.4]
  input  [63:0] io_ins_493, // @[:@35575.4]
  input  [63:0] io_ins_494, // @[:@35575.4]
  input  [63:0] io_ins_495, // @[:@35575.4]
  input  [63:0] io_ins_496, // @[:@35575.4]
  input  [63:0] io_ins_497, // @[:@35575.4]
  input  [63:0] io_ins_498, // @[:@35575.4]
  input  [63:0] io_ins_499, // @[:@35575.4]
  input  [63:0] io_ins_500, // @[:@35575.4]
  input  [63:0] io_ins_501, // @[:@35575.4]
  input  [63:0] io_ins_502, // @[:@35575.4]
  input  [63:0] io_ins_503, // @[:@35575.4]
  input  [63:0] io_ins_504, // @[:@35575.4]
  input  [63:0] io_ins_505, // @[:@35575.4]
  input  [63:0] io_ins_506, // @[:@35575.4]
  input  [63:0] io_ins_507, // @[:@35575.4]
  input  [63:0] io_ins_508, // @[:@35575.4]
  input  [63:0] io_ins_509, // @[:@35575.4]
  input  [63:0] io_ins_510, // @[:@35575.4]
  input  [63:0] io_ins_511, // @[:@35575.4]
  input  [8:0]  io_sel, // @[:@35575.4]
  output [63:0] io_out // @[:@35575.4]
);
  wire [63:0] _GEN_1; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_2; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_3; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_4; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_5; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_6; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_7; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_8; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_9; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_10; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_11; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_12; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_13; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_14; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_15; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_16; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_17; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_18; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_19; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_20; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_21; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_22; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_23; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_24; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_25; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_26; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_27; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_28; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_29; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_30; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_31; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_32; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_33; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_34; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_35; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_36; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_37; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_38; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_39; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_40; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_41; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_42; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_43; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_44; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_45; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_46; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_47; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_48; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_49; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_50; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_51; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_52; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_53; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_54; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_55; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_56; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_57; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_58; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_59; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_60; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_61; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_62; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_63; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_64; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_65; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_66; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_67; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_68; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_69; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_70; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_71; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_72; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_73; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_74; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_75; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_76; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_77; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_78; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_79; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_80; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_81; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_82; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_83; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_84; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_85; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_86; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_87; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_88; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_89; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_90; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_91; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_92; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_93; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_94; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_95; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_96; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_97; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_98; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_99; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_100; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_101; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_102; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_103; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_104; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_105; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_106; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_107; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_108; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_109; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_110; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_111; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_112; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_113; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_114; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_115; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_116; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_117; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_118; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_119; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_120; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_121; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_122; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_123; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_124; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_125; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_126; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_127; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_128; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_129; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_130; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_131; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_132; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_133; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_134; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_135; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_136; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_137; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_138; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_139; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_140; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_141; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_142; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_143; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_144; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_145; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_146; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_147; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_148; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_149; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_150; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_151; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_152; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_153; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_154; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_155; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_156; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_157; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_158; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_159; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_160; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_161; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_162; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_163; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_164; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_165; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_166; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_167; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_168; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_169; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_170; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_171; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_172; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_173; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_174; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_175; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_176; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_177; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_178; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_179; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_180; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_181; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_182; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_183; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_184; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_185; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_186; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_187; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_188; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_189; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_190; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_191; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_192; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_193; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_194; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_195; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_196; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_197; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_198; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_199; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_200; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_201; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_202; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_203; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_204; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_205; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_206; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_207; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_208; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_209; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_210; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_211; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_212; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_213; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_214; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_215; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_216; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_217; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_218; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_219; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_220; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_221; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_222; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_223; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_224; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_225; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_226; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_227; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_228; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_229; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_230; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_231; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_232; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_233; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_234; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_235; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_236; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_237; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_238; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_239; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_240; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_241; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_242; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_243; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_244; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_245; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_246; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_247; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_248; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_249; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_250; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_251; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_252; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_253; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_254; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_255; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_256; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_257; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_258; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_259; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_260; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_261; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_262; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_263; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_264; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_265; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_266; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_267; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_268; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_269; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_270; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_271; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_272; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_273; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_274; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_275; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_276; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_277; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_278; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_279; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_280; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_281; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_282; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_283; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_284; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_285; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_286; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_287; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_288; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_289; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_290; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_291; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_292; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_293; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_294; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_295; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_296; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_297; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_298; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_299; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_300; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_301; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_302; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_303; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_304; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_305; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_306; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_307; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_308; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_309; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_310; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_311; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_312; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_313; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_314; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_315; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_316; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_317; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_318; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_319; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_320; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_321; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_322; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_323; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_324; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_325; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_326; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_327; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_328; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_329; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_330; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_331; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_332; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_333; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_334; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_335; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_336; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_337; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_338; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_339; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_340; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_341; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_342; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_343; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_344; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_345; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_346; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_347; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_348; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_349; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_350; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_351; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_352; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_353; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_354; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_355; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_356; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_357; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_358; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_359; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_360; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_361; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_362; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_363; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_364; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_365; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_366; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_367; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_368; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_369; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_370; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_371; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_372; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_373; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_374; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_375; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_376; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_377; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_378; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_379; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_380; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_381; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_382; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_383; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_384; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_385; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_386; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_387; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_388; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_389; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_390; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_391; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_392; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_393; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_394; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_395; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_396; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_397; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_398; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_399; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_400; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_401; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_402; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_403; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_404; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_405; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_406; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_407; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_408; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_409; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_410; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_411; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_412; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_413; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_414; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_415; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_416; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_417; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_418; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_419; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_420; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_421; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_422; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_423; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_424; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_425; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_426; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_427; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_428; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_429; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_430; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_431; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_432; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_433; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_434; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_435; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_436; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_437; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_438; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_439; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_440; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_441; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_442; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_443; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_444; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_445; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_446; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_447; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_448; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_449; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_450; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_451; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_452; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_453; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_454; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_455; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_456; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_457; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_458; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_459; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_460; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_461; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_462; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_463; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_464; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_465; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_466; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_467; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_468; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_469; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_470; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_471; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_472; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_473; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_474; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_475; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_476; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_477; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_478; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_479; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_480; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_481; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_482; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_483; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_484; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_485; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_486; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_487; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_488; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_489; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_490; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_491; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_492; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_493; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_494; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_495; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_496; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_497; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_498; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_499; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_500; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_501; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_502; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_503; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_504; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_505; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_506; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_507; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_508; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_509; // @[MuxN.scala 16:10:@35577.4]
  wire [63:0] _GEN_510; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_1 = 9'h1 == io_sel ? io_ins_1 : io_ins_0; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_2 = 9'h2 == io_sel ? io_ins_2 : _GEN_1; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_3 = 9'h3 == io_sel ? io_ins_3 : _GEN_2; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_4 = 9'h4 == io_sel ? io_ins_4 : _GEN_3; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_5 = 9'h5 == io_sel ? io_ins_5 : _GEN_4; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_6 = 9'h6 == io_sel ? io_ins_6 : _GEN_5; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_7 = 9'h7 == io_sel ? io_ins_7 : _GEN_6; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_8 = 9'h8 == io_sel ? io_ins_8 : _GEN_7; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_9 = 9'h9 == io_sel ? io_ins_9 : _GEN_8; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_10 = 9'ha == io_sel ? io_ins_10 : _GEN_9; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_11 = 9'hb == io_sel ? io_ins_11 : _GEN_10; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_12 = 9'hc == io_sel ? io_ins_12 : _GEN_11; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_13 = 9'hd == io_sel ? io_ins_13 : _GEN_12; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_14 = 9'he == io_sel ? io_ins_14 : _GEN_13; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_15 = 9'hf == io_sel ? io_ins_15 : _GEN_14; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_16 = 9'h10 == io_sel ? io_ins_16 : _GEN_15; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_17 = 9'h11 == io_sel ? io_ins_17 : _GEN_16; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_18 = 9'h12 == io_sel ? io_ins_18 : _GEN_17; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_19 = 9'h13 == io_sel ? io_ins_19 : _GEN_18; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_20 = 9'h14 == io_sel ? io_ins_20 : _GEN_19; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_21 = 9'h15 == io_sel ? io_ins_21 : _GEN_20; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_22 = 9'h16 == io_sel ? io_ins_22 : _GEN_21; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_23 = 9'h17 == io_sel ? io_ins_23 : _GEN_22; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_24 = 9'h18 == io_sel ? io_ins_24 : _GEN_23; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_25 = 9'h19 == io_sel ? io_ins_25 : _GEN_24; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_26 = 9'h1a == io_sel ? io_ins_26 : _GEN_25; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_27 = 9'h1b == io_sel ? io_ins_27 : _GEN_26; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_28 = 9'h1c == io_sel ? io_ins_28 : _GEN_27; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_29 = 9'h1d == io_sel ? io_ins_29 : _GEN_28; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_30 = 9'h1e == io_sel ? io_ins_30 : _GEN_29; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_31 = 9'h1f == io_sel ? io_ins_31 : _GEN_30; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_32 = 9'h20 == io_sel ? io_ins_32 : _GEN_31; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_33 = 9'h21 == io_sel ? io_ins_33 : _GEN_32; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_34 = 9'h22 == io_sel ? io_ins_34 : _GEN_33; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_35 = 9'h23 == io_sel ? io_ins_35 : _GEN_34; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_36 = 9'h24 == io_sel ? io_ins_36 : _GEN_35; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_37 = 9'h25 == io_sel ? io_ins_37 : _GEN_36; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_38 = 9'h26 == io_sel ? io_ins_38 : _GEN_37; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_39 = 9'h27 == io_sel ? io_ins_39 : _GEN_38; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_40 = 9'h28 == io_sel ? io_ins_40 : _GEN_39; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_41 = 9'h29 == io_sel ? io_ins_41 : _GEN_40; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_42 = 9'h2a == io_sel ? io_ins_42 : _GEN_41; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_43 = 9'h2b == io_sel ? io_ins_43 : _GEN_42; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_44 = 9'h2c == io_sel ? io_ins_44 : _GEN_43; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_45 = 9'h2d == io_sel ? io_ins_45 : _GEN_44; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_46 = 9'h2e == io_sel ? io_ins_46 : _GEN_45; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_47 = 9'h2f == io_sel ? io_ins_47 : _GEN_46; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_48 = 9'h30 == io_sel ? io_ins_48 : _GEN_47; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_49 = 9'h31 == io_sel ? io_ins_49 : _GEN_48; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_50 = 9'h32 == io_sel ? io_ins_50 : _GEN_49; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_51 = 9'h33 == io_sel ? io_ins_51 : _GEN_50; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_52 = 9'h34 == io_sel ? io_ins_52 : _GEN_51; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_53 = 9'h35 == io_sel ? io_ins_53 : _GEN_52; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_54 = 9'h36 == io_sel ? io_ins_54 : _GEN_53; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_55 = 9'h37 == io_sel ? io_ins_55 : _GEN_54; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_56 = 9'h38 == io_sel ? io_ins_56 : _GEN_55; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_57 = 9'h39 == io_sel ? io_ins_57 : _GEN_56; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_58 = 9'h3a == io_sel ? io_ins_58 : _GEN_57; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_59 = 9'h3b == io_sel ? io_ins_59 : _GEN_58; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_60 = 9'h3c == io_sel ? io_ins_60 : _GEN_59; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_61 = 9'h3d == io_sel ? io_ins_61 : _GEN_60; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_62 = 9'h3e == io_sel ? io_ins_62 : _GEN_61; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_63 = 9'h3f == io_sel ? io_ins_63 : _GEN_62; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_64 = 9'h40 == io_sel ? io_ins_64 : _GEN_63; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_65 = 9'h41 == io_sel ? io_ins_65 : _GEN_64; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_66 = 9'h42 == io_sel ? io_ins_66 : _GEN_65; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_67 = 9'h43 == io_sel ? io_ins_67 : _GEN_66; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_68 = 9'h44 == io_sel ? io_ins_68 : _GEN_67; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_69 = 9'h45 == io_sel ? io_ins_69 : _GEN_68; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_70 = 9'h46 == io_sel ? io_ins_70 : _GEN_69; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_71 = 9'h47 == io_sel ? io_ins_71 : _GEN_70; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_72 = 9'h48 == io_sel ? io_ins_72 : _GEN_71; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_73 = 9'h49 == io_sel ? io_ins_73 : _GEN_72; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_74 = 9'h4a == io_sel ? io_ins_74 : _GEN_73; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_75 = 9'h4b == io_sel ? io_ins_75 : _GEN_74; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_76 = 9'h4c == io_sel ? io_ins_76 : _GEN_75; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_77 = 9'h4d == io_sel ? io_ins_77 : _GEN_76; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_78 = 9'h4e == io_sel ? io_ins_78 : _GEN_77; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_79 = 9'h4f == io_sel ? io_ins_79 : _GEN_78; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_80 = 9'h50 == io_sel ? io_ins_80 : _GEN_79; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_81 = 9'h51 == io_sel ? io_ins_81 : _GEN_80; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_82 = 9'h52 == io_sel ? io_ins_82 : _GEN_81; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_83 = 9'h53 == io_sel ? io_ins_83 : _GEN_82; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_84 = 9'h54 == io_sel ? io_ins_84 : _GEN_83; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_85 = 9'h55 == io_sel ? io_ins_85 : _GEN_84; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_86 = 9'h56 == io_sel ? io_ins_86 : _GEN_85; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_87 = 9'h57 == io_sel ? io_ins_87 : _GEN_86; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_88 = 9'h58 == io_sel ? io_ins_88 : _GEN_87; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_89 = 9'h59 == io_sel ? io_ins_89 : _GEN_88; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_90 = 9'h5a == io_sel ? io_ins_90 : _GEN_89; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_91 = 9'h5b == io_sel ? io_ins_91 : _GEN_90; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_92 = 9'h5c == io_sel ? io_ins_92 : _GEN_91; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_93 = 9'h5d == io_sel ? io_ins_93 : _GEN_92; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_94 = 9'h5e == io_sel ? io_ins_94 : _GEN_93; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_95 = 9'h5f == io_sel ? io_ins_95 : _GEN_94; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_96 = 9'h60 == io_sel ? io_ins_96 : _GEN_95; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_97 = 9'h61 == io_sel ? io_ins_97 : _GEN_96; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_98 = 9'h62 == io_sel ? io_ins_98 : _GEN_97; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_99 = 9'h63 == io_sel ? io_ins_99 : _GEN_98; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_100 = 9'h64 == io_sel ? io_ins_100 : _GEN_99; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_101 = 9'h65 == io_sel ? io_ins_101 : _GEN_100; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_102 = 9'h66 == io_sel ? io_ins_102 : _GEN_101; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_103 = 9'h67 == io_sel ? io_ins_103 : _GEN_102; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_104 = 9'h68 == io_sel ? io_ins_104 : _GEN_103; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_105 = 9'h69 == io_sel ? io_ins_105 : _GEN_104; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_106 = 9'h6a == io_sel ? io_ins_106 : _GEN_105; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_107 = 9'h6b == io_sel ? io_ins_107 : _GEN_106; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_108 = 9'h6c == io_sel ? io_ins_108 : _GEN_107; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_109 = 9'h6d == io_sel ? io_ins_109 : _GEN_108; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_110 = 9'h6e == io_sel ? io_ins_110 : _GEN_109; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_111 = 9'h6f == io_sel ? io_ins_111 : _GEN_110; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_112 = 9'h70 == io_sel ? io_ins_112 : _GEN_111; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_113 = 9'h71 == io_sel ? io_ins_113 : _GEN_112; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_114 = 9'h72 == io_sel ? io_ins_114 : _GEN_113; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_115 = 9'h73 == io_sel ? io_ins_115 : _GEN_114; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_116 = 9'h74 == io_sel ? io_ins_116 : _GEN_115; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_117 = 9'h75 == io_sel ? io_ins_117 : _GEN_116; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_118 = 9'h76 == io_sel ? io_ins_118 : _GEN_117; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_119 = 9'h77 == io_sel ? io_ins_119 : _GEN_118; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_120 = 9'h78 == io_sel ? io_ins_120 : _GEN_119; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_121 = 9'h79 == io_sel ? io_ins_121 : _GEN_120; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_122 = 9'h7a == io_sel ? io_ins_122 : _GEN_121; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_123 = 9'h7b == io_sel ? io_ins_123 : _GEN_122; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_124 = 9'h7c == io_sel ? io_ins_124 : _GEN_123; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_125 = 9'h7d == io_sel ? io_ins_125 : _GEN_124; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_126 = 9'h7e == io_sel ? io_ins_126 : _GEN_125; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_127 = 9'h7f == io_sel ? io_ins_127 : _GEN_126; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_128 = 9'h80 == io_sel ? io_ins_128 : _GEN_127; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_129 = 9'h81 == io_sel ? io_ins_129 : _GEN_128; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_130 = 9'h82 == io_sel ? io_ins_130 : _GEN_129; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_131 = 9'h83 == io_sel ? io_ins_131 : _GEN_130; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_132 = 9'h84 == io_sel ? io_ins_132 : _GEN_131; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_133 = 9'h85 == io_sel ? io_ins_133 : _GEN_132; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_134 = 9'h86 == io_sel ? io_ins_134 : _GEN_133; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_135 = 9'h87 == io_sel ? io_ins_135 : _GEN_134; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_136 = 9'h88 == io_sel ? io_ins_136 : _GEN_135; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_137 = 9'h89 == io_sel ? io_ins_137 : _GEN_136; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_138 = 9'h8a == io_sel ? io_ins_138 : _GEN_137; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_139 = 9'h8b == io_sel ? io_ins_139 : _GEN_138; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_140 = 9'h8c == io_sel ? io_ins_140 : _GEN_139; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_141 = 9'h8d == io_sel ? io_ins_141 : _GEN_140; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_142 = 9'h8e == io_sel ? io_ins_142 : _GEN_141; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_143 = 9'h8f == io_sel ? io_ins_143 : _GEN_142; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_144 = 9'h90 == io_sel ? io_ins_144 : _GEN_143; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_145 = 9'h91 == io_sel ? io_ins_145 : _GEN_144; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_146 = 9'h92 == io_sel ? io_ins_146 : _GEN_145; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_147 = 9'h93 == io_sel ? io_ins_147 : _GEN_146; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_148 = 9'h94 == io_sel ? io_ins_148 : _GEN_147; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_149 = 9'h95 == io_sel ? io_ins_149 : _GEN_148; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_150 = 9'h96 == io_sel ? io_ins_150 : _GEN_149; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_151 = 9'h97 == io_sel ? io_ins_151 : _GEN_150; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_152 = 9'h98 == io_sel ? io_ins_152 : _GEN_151; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_153 = 9'h99 == io_sel ? io_ins_153 : _GEN_152; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_154 = 9'h9a == io_sel ? io_ins_154 : _GEN_153; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_155 = 9'h9b == io_sel ? io_ins_155 : _GEN_154; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_156 = 9'h9c == io_sel ? io_ins_156 : _GEN_155; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_157 = 9'h9d == io_sel ? io_ins_157 : _GEN_156; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_158 = 9'h9e == io_sel ? io_ins_158 : _GEN_157; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_159 = 9'h9f == io_sel ? io_ins_159 : _GEN_158; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_160 = 9'ha0 == io_sel ? io_ins_160 : _GEN_159; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_161 = 9'ha1 == io_sel ? io_ins_161 : _GEN_160; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_162 = 9'ha2 == io_sel ? io_ins_162 : _GEN_161; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_163 = 9'ha3 == io_sel ? io_ins_163 : _GEN_162; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_164 = 9'ha4 == io_sel ? io_ins_164 : _GEN_163; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_165 = 9'ha5 == io_sel ? io_ins_165 : _GEN_164; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_166 = 9'ha6 == io_sel ? io_ins_166 : _GEN_165; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_167 = 9'ha7 == io_sel ? io_ins_167 : _GEN_166; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_168 = 9'ha8 == io_sel ? io_ins_168 : _GEN_167; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_169 = 9'ha9 == io_sel ? io_ins_169 : _GEN_168; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_170 = 9'haa == io_sel ? io_ins_170 : _GEN_169; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_171 = 9'hab == io_sel ? io_ins_171 : _GEN_170; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_172 = 9'hac == io_sel ? io_ins_172 : _GEN_171; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_173 = 9'had == io_sel ? io_ins_173 : _GEN_172; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_174 = 9'hae == io_sel ? io_ins_174 : _GEN_173; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_175 = 9'haf == io_sel ? io_ins_175 : _GEN_174; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_176 = 9'hb0 == io_sel ? io_ins_176 : _GEN_175; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_177 = 9'hb1 == io_sel ? io_ins_177 : _GEN_176; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_178 = 9'hb2 == io_sel ? io_ins_178 : _GEN_177; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_179 = 9'hb3 == io_sel ? io_ins_179 : _GEN_178; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_180 = 9'hb4 == io_sel ? io_ins_180 : _GEN_179; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_181 = 9'hb5 == io_sel ? io_ins_181 : _GEN_180; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_182 = 9'hb6 == io_sel ? io_ins_182 : _GEN_181; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_183 = 9'hb7 == io_sel ? io_ins_183 : _GEN_182; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_184 = 9'hb8 == io_sel ? io_ins_184 : _GEN_183; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_185 = 9'hb9 == io_sel ? io_ins_185 : _GEN_184; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_186 = 9'hba == io_sel ? io_ins_186 : _GEN_185; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_187 = 9'hbb == io_sel ? io_ins_187 : _GEN_186; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_188 = 9'hbc == io_sel ? io_ins_188 : _GEN_187; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_189 = 9'hbd == io_sel ? io_ins_189 : _GEN_188; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_190 = 9'hbe == io_sel ? io_ins_190 : _GEN_189; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_191 = 9'hbf == io_sel ? io_ins_191 : _GEN_190; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_192 = 9'hc0 == io_sel ? io_ins_192 : _GEN_191; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_193 = 9'hc1 == io_sel ? io_ins_193 : _GEN_192; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_194 = 9'hc2 == io_sel ? io_ins_194 : _GEN_193; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_195 = 9'hc3 == io_sel ? io_ins_195 : _GEN_194; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_196 = 9'hc4 == io_sel ? io_ins_196 : _GEN_195; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_197 = 9'hc5 == io_sel ? io_ins_197 : _GEN_196; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_198 = 9'hc6 == io_sel ? io_ins_198 : _GEN_197; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_199 = 9'hc7 == io_sel ? io_ins_199 : _GEN_198; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_200 = 9'hc8 == io_sel ? io_ins_200 : _GEN_199; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_201 = 9'hc9 == io_sel ? io_ins_201 : _GEN_200; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_202 = 9'hca == io_sel ? io_ins_202 : _GEN_201; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_203 = 9'hcb == io_sel ? io_ins_203 : _GEN_202; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_204 = 9'hcc == io_sel ? io_ins_204 : _GEN_203; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_205 = 9'hcd == io_sel ? io_ins_205 : _GEN_204; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_206 = 9'hce == io_sel ? io_ins_206 : _GEN_205; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_207 = 9'hcf == io_sel ? io_ins_207 : _GEN_206; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_208 = 9'hd0 == io_sel ? io_ins_208 : _GEN_207; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_209 = 9'hd1 == io_sel ? io_ins_209 : _GEN_208; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_210 = 9'hd2 == io_sel ? io_ins_210 : _GEN_209; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_211 = 9'hd3 == io_sel ? io_ins_211 : _GEN_210; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_212 = 9'hd4 == io_sel ? io_ins_212 : _GEN_211; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_213 = 9'hd5 == io_sel ? io_ins_213 : _GEN_212; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_214 = 9'hd6 == io_sel ? io_ins_214 : _GEN_213; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_215 = 9'hd7 == io_sel ? io_ins_215 : _GEN_214; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_216 = 9'hd8 == io_sel ? io_ins_216 : _GEN_215; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_217 = 9'hd9 == io_sel ? io_ins_217 : _GEN_216; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_218 = 9'hda == io_sel ? io_ins_218 : _GEN_217; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_219 = 9'hdb == io_sel ? io_ins_219 : _GEN_218; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_220 = 9'hdc == io_sel ? io_ins_220 : _GEN_219; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_221 = 9'hdd == io_sel ? io_ins_221 : _GEN_220; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_222 = 9'hde == io_sel ? io_ins_222 : _GEN_221; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_223 = 9'hdf == io_sel ? io_ins_223 : _GEN_222; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_224 = 9'he0 == io_sel ? io_ins_224 : _GEN_223; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_225 = 9'he1 == io_sel ? io_ins_225 : _GEN_224; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_226 = 9'he2 == io_sel ? io_ins_226 : _GEN_225; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_227 = 9'he3 == io_sel ? io_ins_227 : _GEN_226; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_228 = 9'he4 == io_sel ? io_ins_228 : _GEN_227; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_229 = 9'he5 == io_sel ? io_ins_229 : _GEN_228; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_230 = 9'he6 == io_sel ? io_ins_230 : _GEN_229; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_231 = 9'he7 == io_sel ? io_ins_231 : _GEN_230; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_232 = 9'he8 == io_sel ? io_ins_232 : _GEN_231; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_233 = 9'he9 == io_sel ? io_ins_233 : _GEN_232; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_234 = 9'hea == io_sel ? io_ins_234 : _GEN_233; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_235 = 9'heb == io_sel ? io_ins_235 : _GEN_234; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_236 = 9'hec == io_sel ? io_ins_236 : _GEN_235; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_237 = 9'hed == io_sel ? io_ins_237 : _GEN_236; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_238 = 9'hee == io_sel ? io_ins_238 : _GEN_237; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_239 = 9'hef == io_sel ? io_ins_239 : _GEN_238; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_240 = 9'hf0 == io_sel ? io_ins_240 : _GEN_239; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_241 = 9'hf1 == io_sel ? io_ins_241 : _GEN_240; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_242 = 9'hf2 == io_sel ? io_ins_242 : _GEN_241; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_243 = 9'hf3 == io_sel ? io_ins_243 : _GEN_242; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_244 = 9'hf4 == io_sel ? io_ins_244 : _GEN_243; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_245 = 9'hf5 == io_sel ? io_ins_245 : _GEN_244; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_246 = 9'hf6 == io_sel ? io_ins_246 : _GEN_245; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_247 = 9'hf7 == io_sel ? io_ins_247 : _GEN_246; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_248 = 9'hf8 == io_sel ? io_ins_248 : _GEN_247; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_249 = 9'hf9 == io_sel ? io_ins_249 : _GEN_248; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_250 = 9'hfa == io_sel ? io_ins_250 : _GEN_249; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_251 = 9'hfb == io_sel ? io_ins_251 : _GEN_250; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_252 = 9'hfc == io_sel ? io_ins_252 : _GEN_251; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_253 = 9'hfd == io_sel ? io_ins_253 : _GEN_252; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_254 = 9'hfe == io_sel ? io_ins_254 : _GEN_253; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_255 = 9'hff == io_sel ? io_ins_255 : _GEN_254; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_256 = 9'h100 == io_sel ? io_ins_256 : _GEN_255; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_257 = 9'h101 == io_sel ? io_ins_257 : _GEN_256; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_258 = 9'h102 == io_sel ? io_ins_258 : _GEN_257; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_259 = 9'h103 == io_sel ? io_ins_259 : _GEN_258; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_260 = 9'h104 == io_sel ? io_ins_260 : _GEN_259; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_261 = 9'h105 == io_sel ? io_ins_261 : _GEN_260; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_262 = 9'h106 == io_sel ? io_ins_262 : _GEN_261; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_263 = 9'h107 == io_sel ? io_ins_263 : _GEN_262; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_264 = 9'h108 == io_sel ? io_ins_264 : _GEN_263; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_265 = 9'h109 == io_sel ? io_ins_265 : _GEN_264; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_266 = 9'h10a == io_sel ? io_ins_266 : _GEN_265; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_267 = 9'h10b == io_sel ? io_ins_267 : _GEN_266; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_268 = 9'h10c == io_sel ? io_ins_268 : _GEN_267; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_269 = 9'h10d == io_sel ? io_ins_269 : _GEN_268; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_270 = 9'h10e == io_sel ? io_ins_270 : _GEN_269; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_271 = 9'h10f == io_sel ? io_ins_271 : _GEN_270; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_272 = 9'h110 == io_sel ? io_ins_272 : _GEN_271; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_273 = 9'h111 == io_sel ? io_ins_273 : _GEN_272; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_274 = 9'h112 == io_sel ? io_ins_274 : _GEN_273; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_275 = 9'h113 == io_sel ? io_ins_275 : _GEN_274; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_276 = 9'h114 == io_sel ? io_ins_276 : _GEN_275; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_277 = 9'h115 == io_sel ? io_ins_277 : _GEN_276; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_278 = 9'h116 == io_sel ? io_ins_278 : _GEN_277; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_279 = 9'h117 == io_sel ? io_ins_279 : _GEN_278; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_280 = 9'h118 == io_sel ? io_ins_280 : _GEN_279; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_281 = 9'h119 == io_sel ? io_ins_281 : _GEN_280; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_282 = 9'h11a == io_sel ? io_ins_282 : _GEN_281; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_283 = 9'h11b == io_sel ? io_ins_283 : _GEN_282; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_284 = 9'h11c == io_sel ? io_ins_284 : _GEN_283; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_285 = 9'h11d == io_sel ? io_ins_285 : _GEN_284; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_286 = 9'h11e == io_sel ? io_ins_286 : _GEN_285; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_287 = 9'h11f == io_sel ? io_ins_287 : _GEN_286; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_288 = 9'h120 == io_sel ? io_ins_288 : _GEN_287; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_289 = 9'h121 == io_sel ? io_ins_289 : _GEN_288; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_290 = 9'h122 == io_sel ? io_ins_290 : _GEN_289; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_291 = 9'h123 == io_sel ? io_ins_291 : _GEN_290; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_292 = 9'h124 == io_sel ? io_ins_292 : _GEN_291; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_293 = 9'h125 == io_sel ? io_ins_293 : _GEN_292; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_294 = 9'h126 == io_sel ? io_ins_294 : _GEN_293; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_295 = 9'h127 == io_sel ? io_ins_295 : _GEN_294; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_296 = 9'h128 == io_sel ? io_ins_296 : _GEN_295; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_297 = 9'h129 == io_sel ? io_ins_297 : _GEN_296; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_298 = 9'h12a == io_sel ? io_ins_298 : _GEN_297; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_299 = 9'h12b == io_sel ? io_ins_299 : _GEN_298; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_300 = 9'h12c == io_sel ? io_ins_300 : _GEN_299; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_301 = 9'h12d == io_sel ? io_ins_301 : _GEN_300; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_302 = 9'h12e == io_sel ? io_ins_302 : _GEN_301; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_303 = 9'h12f == io_sel ? io_ins_303 : _GEN_302; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_304 = 9'h130 == io_sel ? io_ins_304 : _GEN_303; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_305 = 9'h131 == io_sel ? io_ins_305 : _GEN_304; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_306 = 9'h132 == io_sel ? io_ins_306 : _GEN_305; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_307 = 9'h133 == io_sel ? io_ins_307 : _GEN_306; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_308 = 9'h134 == io_sel ? io_ins_308 : _GEN_307; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_309 = 9'h135 == io_sel ? io_ins_309 : _GEN_308; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_310 = 9'h136 == io_sel ? io_ins_310 : _GEN_309; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_311 = 9'h137 == io_sel ? io_ins_311 : _GEN_310; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_312 = 9'h138 == io_sel ? io_ins_312 : _GEN_311; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_313 = 9'h139 == io_sel ? io_ins_313 : _GEN_312; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_314 = 9'h13a == io_sel ? io_ins_314 : _GEN_313; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_315 = 9'h13b == io_sel ? io_ins_315 : _GEN_314; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_316 = 9'h13c == io_sel ? io_ins_316 : _GEN_315; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_317 = 9'h13d == io_sel ? io_ins_317 : _GEN_316; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_318 = 9'h13e == io_sel ? io_ins_318 : _GEN_317; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_319 = 9'h13f == io_sel ? io_ins_319 : _GEN_318; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_320 = 9'h140 == io_sel ? io_ins_320 : _GEN_319; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_321 = 9'h141 == io_sel ? io_ins_321 : _GEN_320; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_322 = 9'h142 == io_sel ? io_ins_322 : _GEN_321; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_323 = 9'h143 == io_sel ? io_ins_323 : _GEN_322; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_324 = 9'h144 == io_sel ? io_ins_324 : _GEN_323; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_325 = 9'h145 == io_sel ? io_ins_325 : _GEN_324; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_326 = 9'h146 == io_sel ? io_ins_326 : _GEN_325; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_327 = 9'h147 == io_sel ? io_ins_327 : _GEN_326; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_328 = 9'h148 == io_sel ? io_ins_328 : _GEN_327; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_329 = 9'h149 == io_sel ? io_ins_329 : _GEN_328; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_330 = 9'h14a == io_sel ? io_ins_330 : _GEN_329; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_331 = 9'h14b == io_sel ? io_ins_331 : _GEN_330; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_332 = 9'h14c == io_sel ? io_ins_332 : _GEN_331; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_333 = 9'h14d == io_sel ? io_ins_333 : _GEN_332; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_334 = 9'h14e == io_sel ? io_ins_334 : _GEN_333; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_335 = 9'h14f == io_sel ? io_ins_335 : _GEN_334; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_336 = 9'h150 == io_sel ? io_ins_336 : _GEN_335; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_337 = 9'h151 == io_sel ? io_ins_337 : _GEN_336; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_338 = 9'h152 == io_sel ? io_ins_338 : _GEN_337; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_339 = 9'h153 == io_sel ? io_ins_339 : _GEN_338; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_340 = 9'h154 == io_sel ? io_ins_340 : _GEN_339; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_341 = 9'h155 == io_sel ? io_ins_341 : _GEN_340; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_342 = 9'h156 == io_sel ? io_ins_342 : _GEN_341; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_343 = 9'h157 == io_sel ? io_ins_343 : _GEN_342; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_344 = 9'h158 == io_sel ? io_ins_344 : _GEN_343; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_345 = 9'h159 == io_sel ? io_ins_345 : _GEN_344; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_346 = 9'h15a == io_sel ? io_ins_346 : _GEN_345; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_347 = 9'h15b == io_sel ? io_ins_347 : _GEN_346; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_348 = 9'h15c == io_sel ? io_ins_348 : _GEN_347; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_349 = 9'h15d == io_sel ? io_ins_349 : _GEN_348; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_350 = 9'h15e == io_sel ? io_ins_350 : _GEN_349; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_351 = 9'h15f == io_sel ? io_ins_351 : _GEN_350; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_352 = 9'h160 == io_sel ? io_ins_352 : _GEN_351; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_353 = 9'h161 == io_sel ? io_ins_353 : _GEN_352; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_354 = 9'h162 == io_sel ? io_ins_354 : _GEN_353; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_355 = 9'h163 == io_sel ? io_ins_355 : _GEN_354; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_356 = 9'h164 == io_sel ? io_ins_356 : _GEN_355; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_357 = 9'h165 == io_sel ? io_ins_357 : _GEN_356; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_358 = 9'h166 == io_sel ? io_ins_358 : _GEN_357; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_359 = 9'h167 == io_sel ? io_ins_359 : _GEN_358; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_360 = 9'h168 == io_sel ? io_ins_360 : _GEN_359; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_361 = 9'h169 == io_sel ? io_ins_361 : _GEN_360; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_362 = 9'h16a == io_sel ? io_ins_362 : _GEN_361; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_363 = 9'h16b == io_sel ? io_ins_363 : _GEN_362; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_364 = 9'h16c == io_sel ? io_ins_364 : _GEN_363; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_365 = 9'h16d == io_sel ? io_ins_365 : _GEN_364; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_366 = 9'h16e == io_sel ? io_ins_366 : _GEN_365; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_367 = 9'h16f == io_sel ? io_ins_367 : _GEN_366; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_368 = 9'h170 == io_sel ? io_ins_368 : _GEN_367; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_369 = 9'h171 == io_sel ? io_ins_369 : _GEN_368; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_370 = 9'h172 == io_sel ? io_ins_370 : _GEN_369; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_371 = 9'h173 == io_sel ? io_ins_371 : _GEN_370; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_372 = 9'h174 == io_sel ? io_ins_372 : _GEN_371; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_373 = 9'h175 == io_sel ? io_ins_373 : _GEN_372; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_374 = 9'h176 == io_sel ? io_ins_374 : _GEN_373; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_375 = 9'h177 == io_sel ? io_ins_375 : _GEN_374; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_376 = 9'h178 == io_sel ? io_ins_376 : _GEN_375; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_377 = 9'h179 == io_sel ? io_ins_377 : _GEN_376; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_378 = 9'h17a == io_sel ? io_ins_378 : _GEN_377; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_379 = 9'h17b == io_sel ? io_ins_379 : _GEN_378; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_380 = 9'h17c == io_sel ? io_ins_380 : _GEN_379; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_381 = 9'h17d == io_sel ? io_ins_381 : _GEN_380; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_382 = 9'h17e == io_sel ? io_ins_382 : _GEN_381; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_383 = 9'h17f == io_sel ? io_ins_383 : _GEN_382; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_384 = 9'h180 == io_sel ? io_ins_384 : _GEN_383; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_385 = 9'h181 == io_sel ? io_ins_385 : _GEN_384; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_386 = 9'h182 == io_sel ? io_ins_386 : _GEN_385; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_387 = 9'h183 == io_sel ? io_ins_387 : _GEN_386; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_388 = 9'h184 == io_sel ? io_ins_388 : _GEN_387; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_389 = 9'h185 == io_sel ? io_ins_389 : _GEN_388; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_390 = 9'h186 == io_sel ? io_ins_390 : _GEN_389; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_391 = 9'h187 == io_sel ? io_ins_391 : _GEN_390; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_392 = 9'h188 == io_sel ? io_ins_392 : _GEN_391; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_393 = 9'h189 == io_sel ? io_ins_393 : _GEN_392; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_394 = 9'h18a == io_sel ? io_ins_394 : _GEN_393; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_395 = 9'h18b == io_sel ? io_ins_395 : _GEN_394; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_396 = 9'h18c == io_sel ? io_ins_396 : _GEN_395; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_397 = 9'h18d == io_sel ? io_ins_397 : _GEN_396; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_398 = 9'h18e == io_sel ? io_ins_398 : _GEN_397; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_399 = 9'h18f == io_sel ? io_ins_399 : _GEN_398; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_400 = 9'h190 == io_sel ? io_ins_400 : _GEN_399; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_401 = 9'h191 == io_sel ? io_ins_401 : _GEN_400; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_402 = 9'h192 == io_sel ? io_ins_402 : _GEN_401; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_403 = 9'h193 == io_sel ? io_ins_403 : _GEN_402; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_404 = 9'h194 == io_sel ? io_ins_404 : _GEN_403; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_405 = 9'h195 == io_sel ? io_ins_405 : _GEN_404; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_406 = 9'h196 == io_sel ? io_ins_406 : _GEN_405; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_407 = 9'h197 == io_sel ? io_ins_407 : _GEN_406; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_408 = 9'h198 == io_sel ? io_ins_408 : _GEN_407; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_409 = 9'h199 == io_sel ? io_ins_409 : _GEN_408; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_410 = 9'h19a == io_sel ? io_ins_410 : _GEN_409; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_411 = 9'h19b == io_sel ? io_ins_411 : _GEN_410; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_412 = 9'h19c == io_sel ? io_ins_412 : _GEN_411; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_413 = 9'h19d == io_sel ? io_ins_413 : _GEN_412; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_414 = 9'h19e == io_sel ? io_ins_414 : _GEN_413; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_415 = 9'h19f == io_sel ? io_ins_415 : _GEN_414; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_416 = 9'h1a0 == io_sel ? io_ins_416 : _GEN_415; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_417 = 9'h1a1 == io_sel ? io_ins_417 : _GEN_416; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_418 = 9'h1a2 == io_sel ? io_ins_418 : _GEN_417; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_419 = 9'h1a3 == io_sel ? io_ins_419 : _GEN_418; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_420 = 9'h1a4 == io_sel ? io_ins_420 : _GEN_419; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_421 = 9'h1a5 == io_sel ? io_ins_421 : _GEN_420; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_422 = 9'h1a6 == io_sel ? io_ins_422 : _GEN_421; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_423 = 9'h1a7 == io_sel ? io_ins_423 : _GEN_422; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_424 = 9'h1a8 == io_sel ? io_ins_424 : _GEN_423; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_425 = 9'h1a9 == io_sel ? io_ins_425 : _GEN_424; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_426 = 9'h1aa == io_sel ? io_ins_426 : _GEN_425; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_427 = 9'h1ab == io_sel ? io_ins_427 : _GEN_426; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_428 = 9'h1ac == io_sel ? io_ins_428 : _GEN_427; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_429 = 9'h1ad == io_sel ? io_ins_429 : _GEN_428; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_430 = 9'h1ae == io_sel ? io_ins_430 : _GEN_429; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_431 = 9'h1af == io_sel ? io_ins_431 : _GEN_430; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_432 = 9'h1b0 == io_sel ? io_ins_432 : _GEN_431; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_433 = 9'h1b1 == io_sel ? io_ins_433 : _GEN_432; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_434 = 9'h1b2 == io_sel ? io_ins_434 : _GEN_433; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_435 = 9'h1b3 == io_sel ? io_ins_435 : _GEN_434; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_436 = 9'h1b4 == io_sel ? io_ins_436 : _GEN_435; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_437 = 9'h1b5 == io_sel ? io_ins_437 : _GEN_436; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_438 = 9'h1b6 == io_sel ? io_ins_438 : _GEN_437; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_439 = 9'h1b7 == io_sel ? io_ins_439 : _GEN_438; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_440 = 9'h1b8 == io_sel ? io_ins_440 : _GEN_439; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_441 = 9'h1b9 == io_sel ? io_ins_441 : _GEN_440; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_442 = 9'h1ba == io_sel ? io_ins_442 : _GEN_441; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_443 = 9'h1bb == io_sel ? io_ins_443 : _GEN_442; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_444 = 9'h1bc == io_sel ? io_ins_444 : _GEN_443; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_445 = 9'h1bd == io_sel ? io_ins_445 : _GEN_444; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_446 = 9'h1be == io_sel ? io_ins_446 : _GEN_445; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_447 = 9'h1bf == io_sel ? io_ins_447 : _GEN_446; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_448 = 9'h1c0 == io_sel ? io_ins_448 : _GEN_447; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_449 = 9'h1c1 == io_sel ? io_ins_449 : _GEN_448; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_450 = 9'h1c2 == io_sel ? io_ins_450 : _GEN_449; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_451 = 9'h1c3 == io_sel ? io_ins_451 : _GEN_450; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_452 = 9'h1c4 == io_sel ? io_ins_452 : _GEN_451; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_453 = 9'h1c5 == io_sel ? io_ins_453 : _GEN_452; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_454 = 9'h1c6 == io_sel ? io_ins_454 : _GEN_453; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_455 = 9'h1c7 == io_sel ? io_ins_455 : _GEN_454; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_456 = 9'h1c8 == io_sel ? io_ins_456 : _GEN_455; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_457 = 9'h1c9 == io_sel ? io_ins_457 : _GEN_456; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_458 = 9'h1ca == io_sel ? io_ins_458 : _GEN_457; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_459 = 9'h1cb == io_sel ? io_ins_459 : _GEN_458; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_460 = 9'h1cc == io_sel ? io_ins_460 : _GEN_459; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_461 = 9'h1cd == io_sel ? io_ins_461 : _GEN_460; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_462 = 9'h1ce == io_sel ? io_ins_462 : _GEN_461; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_463 = 9'h1cf == io_sel ? io_ins_463 : _GEN_462; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_464 = 9'h1d0 == io_sel ? io_ins_464 : _GEN_463; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_465 = 9'h1d1 == io_sel ? io_ins_465 : _GEN_464; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_466 = 9'h1d2 == io_sel ? io_ins_466 : _GEN_465; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_467 = 9'h1d3 == io_sel ? io_ins_467 : _GEN_466; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_468 = 9'h1d4 == io_sel ? io_ins_468 : _GEN_467; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_469 = 9'h1d5 == io_sel ? io_ins_469 : _GEN_468; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_470 = 9'h1d6 == io_sel ? io_ins_470 : _GEN_469; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_471 = 9'h1d7 == io_sel ? io_ins_471 : _GEN_470; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_472 = 9'h1d8 == io_sel ? io_ins_472 : _GEN_471; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_473 = 9'h1d9 == io_sel ? io_ins_473 : _GEN_472; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_474 = 9'h1da == io_sel ? io_ins_474 : _GEN_473; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_475 = 9'h1db == io_sel ? io_ins_475 : _GEN_474; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_476 = 9'h1dc == io_sel ? io_ins_476 : _GEN_475; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_477 = 9'h1dd == io_sel ? io_ins_477 : _GEN_476; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_478 = 9'h1de == io_sel ? io_ins_478 : _GEN_477; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_479 = 9'h1df == io_sel ? io_ins_479 : _GEN_478; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_480 = 9'h1e0 == io_sel ? io_ins_480 : _GEN_479; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_481 = 9'h1e1 == io_sel ? io_ins_481 : _GEN_480; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_482 = 9'h1e2 == io_sel ? io_ins_482 : _GEN_481; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_483 = 9'h1e3 == io_sel ? io_ins_483 : _GEN_482; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_484 = 9'h1e4 == io_sel ? io_ins_484 : _GEN_483; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_485 = 9'h1e5 == io_sel ? io_ins_485 : _GEN_484; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_486 = 9'h1e6 == io_sel ? io_ins_486 : _GEN_485; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_487 = 9'h1e7 == io_sel ? io_ins_487 : _GEN_486; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_488 = 9'h1e8 == io_sel ? io_ins_488 : _GEN_487; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_489 = 9'h1e9 == io_sel ? io_ins_489 : _GEN_488; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_490 = 9'h1ea == io_sel ? io_ins_490 : _GEN_489; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_491 = 9'h1eb == io_sel ? io_ins_491 : _GEN_490; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_492 = 9'h1ec == io_sel ? io_ins_492 : _GEN_491; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_493 = 9'h1ed == io_sel ? io_ins_493 : _GEN_492; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_494 = 9'h1ee == io_sel ? io_ins_494 : _GEN_493; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_495 = 9'h1ef == io_sel ? io_ins_495 : _GEN_494; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_496 = 9'h1f0 == io_sel ? io_ins_496 : _GEN_495; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_497 = 9'h1f1 == io_sel ? io_ins_497 : _GEN_496; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_498 = 9'h1f2 == io_sel ? io_ins_498 : _GEN_497; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_499 = 9'h1f3 == io_sel ? io_ins_499 : _GEN_498; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_500 = 9'h1f4 == io_sel ? io_ins_500 : _GEN_499; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_501 = 9'h1f5 == io_sel ? io_ins_501 : _GEN_500; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_502 = 9'h1f6 == io_sel ? io_ins_502 : _GEN_501; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_503 = 9'h1f7 == io_sel ? io_ins_503 : _GEN_502; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_504 = 9'h1f8 == io_sel ? io_ins_504 : _GEN_503; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_505 = 9'h1f9 == io_sel ? io_ins_505 : _GEN_504; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_506 = 9'h1fa == io_sel ? io_ins_506 : _GEN_505; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_507 = 9'h1fb == io_sel ? io_ins_507 : _GEN_506; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_508 = 9'h1fc == io_sel ? io_ins_508 : _GEN_507; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_509 = 9'h1fd == io_sel ? io_ins_509 : _GEN_508; // @[MuxN.scala 16:10:@35577.4]
  assign _GEN_510 = 9'h1fe == io_sel ? io_ins_510 : _GEN_509; // @[MuxN.scala 16:10:@35577.4]
  assign io_out = 9'h1ff == io_sel ? io_ins_511 : _GEN_510; // @[MuxN.scala 16:10:@35577.4]
endmodule
module RegFile( // @[:@35579.2]
  input         clock, // @[:@35580.4]
  input         reset, // @[:@35581.4]
  input  [31:0] io_raddr, // @[:@35582.4]
  input         io_wen, // @[:@35582.4]
  input  [31:0] io_waddr, // @[:@35582.4]
  input  [63:0] io_wdata, // @[:@35582.4]
  output [63:0] io_rdata, // @[:@35582.4]
  input         io_reset, // @[:@35582.4]
  output [63:0] io_argIns_0, // @[:@35582.4]
  output [63:0] io_argIns_1, // @[:@35582.4]
  output [63:0] io_argIns_2, // @[:@35582.4]
  input         io_argOuts_0_valid, // @[:@35582.4]
  input  [63:0] io_argOuts_0_bits, // @[:@35582.4]
  input         io_argOuts_1_valid, // @[:@35582.4]
  input  [63:0] io_argOuts_1_bits, // @[:@35582.4]
  input         io_argOuts_2_valid, // @[:@35582.4]
  input  [63:0] io_argOuts_2_bits, // @[:@35582.4]
  input         io_argOuts_3_valid, // @[:@35582.4]
  input  [63:0] io_argOuts_3_bits, // @[:@35582.4]
  input         io_argOuts_4_valid, // @[:@35582.4]
  input  [63:0] io_argOuts_4_bits, // @[:@35582.4]
  input         io_argOuts_5_valid, // @[:@35582.4]
  input  [63:0] io_argOuts_5_bits, // @[:@35582.4]
  input         io_argOuts_6_valid, // @[:@35582.4]
  input  [63:0] io_argOuts_6_bits, // @[:@35582.4]
  input         io_argOuts_7_valid, // @[:@35582.4]
  input  [63:0] io_argOuts_7_bits, // @[:@35582.4]
  input         io_argOuts_8_valid, // @[:@35582.4]
  input  [63:0] io_argOuts_8_bits, // @[:@35582.4]
  input         io_argOuts_9_valid, // @[:@35582.4]
  input  [63:0] io_argOuts_9_bits, // @[:@35582.4]
  input         io_argOuts_10_valid, // @[:@35582.4]
  input  [63:0] io_argOuts_10_bits // @[:@35582.4]
);
  wire  regs_0_clock; // @[RegFile.scala 66:20:@37628.4]
  wire  regs_0_reset; // @[RegFile.scala 66:20:@37628.4]
  wire [63:0] regs_0_io_in; // @[RegFile.scala 66:20:@37628.4]
  wire  regs_0_io_reset; // @[RegFile.scala 66:20:@37628.4]
  wire [63:0] regs_0_io_out; // @[RegFile.scala 66:20:@37628.4]
  wire  regs_0_io_enable; // @[RegFile.scala 66:20:@37628.4]
  wire  regs_1_clock; // @[RegFile.scala 66:20:@37640.4]
  wire  regs_1_reset; // @[RegFile.scala 66:20:@37640.4]
  wire [63:0] regs_1_io_in; // @[RegFile.scala 66:20:@37640.4]
  wire  regs_1_io_reset; // @[RegFile.scala 66:20:@37640.4]
  wire [63:0] regs_1_io_out; // @[RegFile.scala 66:20:@37640.4]
  wire  regs_1_io_enable; // @[RegFile.scala 66:20:@37640.4]
  wire  regs_2_clock; // @[RegFile.scala 66:20:@37659.4]
  wire  regs_2_reset; // @[RegFile.scala 66:20:@37659.4]
  wire [63:0] regs_2_io_in; // @[RegFile.scala 66:20:@37659.4]
  wire  regs_2_io_reset; // @[RegFile.scala 66:20:@37659.4]
  wire [63:0] regs_2_io_out; // @[RegFile.scala 66:20:@37659.4]
  wire  regs_2_io_enable; // @[RegFile.scala 66:20:@37659.4]
  wire  regs_3_clock; // @[RegFile.scala 66:20:@37671.4]
  wire  regs_3_reset; // @[RegFile.scala 66:20:@37671.4]
  wire [63:0] regs_3_io_in; // @[RegFile.scala 66:20:@37671.4]
  wire  regs_3_io_reset; // @[RegFile.scala 66:20:@37671.4]
  wire [63:0] regs_3_io_out; // @[RegFile.scala 66:20:@37671.4]
  wire  regs_3_io_enable; // @[RegFile.scala 66:20:@37671.4]
  wire  regs_4_clock; // @[RegFile.scala 66:20:@37685.4]
  wire  regs_4_reset; // @[RegFile.scala 66:20:@37685.4]
  wire [63:0] regs_4_io_in; // @[RegFile.scala 66:20:@37685.4]
  wire  regs_4_io_reset; // @[RegFile.scala 66:20:@37685.4]
  wire [63:0] regs_4_io_out; // @[RegFile.scala 66:20:@37685.4]
  wire  regs_4_io_enable; // @[RegFile.scala 66:20:@37685.4]
  wire  regs_5_clock; // @[RegFile.scala 66:20:@37699.4]
  wire  regs_5_reset; // @[RegFile.scala 66:20:@37699.4]
  wire [63:0] regs_5_io_in; // @[RegFile.scala 66:20:@37699.4]
  wire  regs_5_io_reset; // @[RegFile.scala 66:20:@37699.4]
  wire [63:0] regs_5_io_out; // @[RegFile.scala 66:20:@37699.4]
  wire  regs_5_io_enable; // @[RegFile.scala 66:20:@37699.4]
  wire  regs_6_clock; // @[RegFile.scala 66:20:@37713.4]
  wire  regs_6_reset; // @[RegFile.scala 66:20:@37713.4]
  wire [63:0] regs_6_io_in; // @[RegFile.scala 66:20:@37713.4]
  wire  regs_6_io_reset; // @[RegFile.scala 66:20:@37713.4]
  wire [63:0] regs_6_io_out; // @[RegFile.scala 66:20:@37713.4]
  wire  regs_6_io_enable; // @[RegFile.scala 66:20:@37713.4]
  wire  regs_7_clock; // @[RegFile.scala 66:20:@37727.4]
  wire  regs_7_reset; // @[RegFile.scala 66:20:@37727.4]
  wire [63:0] regs_7_io_in; // @[RegFile.scala 66:20:@37727.4]
  wire  regs_7_io_reset; // @[RegFile.scala 66:20:@37727.4]
  wire [63:0] regs_7_io_out; // @[RegFile.scala 66:20:@37727.4]
  wire  regs_7_io_enable; // @[RegFile.scala 66:20:@37727.4]
  wire  regs_8_clock; // @[RegFile.scala 66:20:@37741.4]
  wire  regs_8_reset; // @[RegFile.scala 66:20:@37741.4]
  wire [63:0] regs_8_io_in; // @[RegFile.scala 66:20:@37741.4]
  wire  regs_8_io_reset; // @[RegFile.scala 66:20:@37741.4]
  wire [63:0] regs_8_io_out; // @[RegFile.scala 66:20:@37741.4]
  wire  regs_8_io_enable; // @[RegFile.scala 66:20:@37741.4]
  wire  regs_9_clock; // @[RegFile.scala 66:20:@37755.4]
  wire  regs_9_reset; // @[RegFile.scala 66:20:@37755.4]
  wire [63:0] regs_9_io_in; // @[RegFile.scala 66:20:@37755.4]
  wire  regs_9_io_reset; // @[RegFile.scala 66:20:@37755.4]
  wire [63:0] regs_9_io_out; // @[RegFile.scala 66:20:@37755.4]
  wire  regs_9_io_enable; // @[RegFile.scala 66:20:@37755.4]
  wire  regs_10_clock; // @[RegFile.scala 66:20:@37769.4]
  wire  regs_10_reset; // @[RegFile.scala 66:20:@37769.4]
  wire [63:0] regs_10_io_in; // @[RegFile.scala 66:20:@37769.4]
  wire  regs_10_io_reset; // @[RegFile.scala 66:20:@37769.4]
  wire [63:0] regs_10_io_out; // @[RegFile.scala 66:20:@37769.4]
  wire  regs_10_io_enable; // @[RegFile.scala 66:20:@37769.4]
  wire  regs_11_clock; // @[RegFile.scala 66:20:@37783.4]
  wire  regs_11_reset; // @[RegFile.scala 66:20:@37783.4]
  wire [63:0] regs_11_io_in; // @[RegFile.scala 66:20:@37783.4]
  wire  regs_11_io_reset; // @[RegFile.scala 66:20:@37783.4]
  wire [63:0] regs_11_io_out; // @[RegFile.scala 66:20:@37783.4]
  wire  regs_11_io_enable; // @[RegFile.scala 66:20:@37783.4]
  wire  regs_12_clock; // @[RegFile.scala 66:20:@37797.4]
  wire  regs_12_reset; // @[RegFile.scala 66:20:@37797.4]
  wire [63:0] regs_12_io_in; // @[RegFile.scala 66:20:@37797.4]
  wire  regs_12_io_reset; // @[RegFile.scala 66:20:@37797.4]
  wire [63:0] regs_12_io_out; // @[RegFile.scala 66:20:@37797.4]
  wire  regs_12_io_enable; // @[RegFile.scala 66:20:@37797.4]
  wire  regs_13_clock; // @[RegFile.scala 66:20:@37811.4]
  wire  regs_13_reset; // @[RegFile.scala 66:20:@37811.4]
  wire [63:0] regs_13_io_in; // @[RegFile.scala 66:20:@37811.4]
  wire  regs_13_io_reset; // @[RegFile.scala 66:20:@37811.4]
  wire [63:0] regs_13_io_out; // @[RegFile.scala 66:20:@37811.4]
  wire  regs_13_io_enable; // @[RegFile.scala 66:20:@37811.4]
  wire  regs_14_clock; // @[RegFile.scala 66:20:@37825.4]
  wire  regs_14_reset; // @[RegFile.scala 66:20:@37825.4]
  wire [63:0] regs_14_io_in; // @[RegFile.scala 66:20:@37825.4]
  wire  regs_14_io_reset; // @[RegFile.scala 66:20:@37825.4]
  wire [63:0] regs_14_io_out; // @[RegFile.scala 66:20:@37825.4]
  wire  regs_14_io_enable; // @[RegFile.scala 66:20:@37825.4]
  wire  regs_15_clock; // @[RegFile.scala 66:20:@37839.4]
  wire  regs_15_reset; // @[RegFile.scala 66:20:@37839.4]
  wire [63:0] regs_15_io_in; // @[RegFile.scala 66:20:@37839.4]
  wire  regs_15_io_reset; // @[RegFile.scala 66:20:@37839.4]
  wire [63:0] regs_15_io_out; // @[RegFile.scala 66:20:@37839.4]
  wire  regs_15_io_enable; // @[RegFile.scala 66:20:@37839.4]
  wire  regs_16_clock; // @[RegFile.scala 66:20:@37853.4]
  wire  regs_16_reset; // @[RegFile.scala 66:20:@37853.4]
  wire [63:0] regs_16_io_in; // @[RegFile.scala 66:20:@37853.4]
  wire  regs_16_io_reset; // @[RegFile.scala 66:20:@37853.4]
  wire [63:0] regs_16_io_out; // @[RegFile.scala 66:20:@37853.4]
  wire  regs_16_io_enable; // @[RegFile.scala 66:20:@37853.4]
  wire  regs_17_clock; // @[RegFile.scala 66:20:@37867.4]
  wire  regs_17_reset; // @[RegFile.scala 66:20:@37867.4]
  wire [63:0] regs_17_io_in; // @[RegFile.scala 66:20:@37867.4]
  wire  regs_17_io_reset; // @[RegFile.scala 66:20:@37867.4]
  wire [63:0] regs_17_io_out; // @[RegFile.scala 66:20:@37867.4]
  wire  regs_17_io_enable; // @[RegFile.scala 66:20:@37867.4]
  wire  regs_18_clock; // @[RegFile.scala 66:20:@37881.4]
  wire  regs_18_reset; // @[RegFile.scala 66:20:@37881.4]
  wire [63:0] regs_18_io_in; // @[RegFile.scala 66:20:@37881.4]
  wire  regs_18_io_reset; // @[RegFile.scala 66:20:@37881.4]
  wire [63:0] regs_18_io_out; // @[RegFile.scala 66:20:@37881.4]
  wire  regs_18_io_enable; // @[RegFile.scala 66:20:@37881.4]
  wire  regs_19_clock; // @[RegFile.scala 66:20:@37895.4]
  wire  regs_19_reset; // @[RegFile.scala 66:20:@37895.4]
  wire [63:0] regs_19_io_in; // @[RegFile.scala 66:20:@37895.4]
  wire  regs_19_io_reset; // @[RegFile.scala 66:20:@37895.4]
  wire [63:0] regs_19_io_out; // @[RegFile.scala 66:20:@37895.4]
  wire  regs_19_io_enable; // @[RegFile.scala 66:20:@37895.4]
  wire  regs_20_clock; // @[RegFile.scala 66:20:@37909.4]
  wire  regs_20_reset; // @[RegFile.scala 66:20:@37909.4]
  wire [63:0] regs_20_io_in; // @[RegFile.scala 66:20:@37909.4]
  wire  regs_20_io_reset; // @[RegFile.scala 66:20:@37909.4]
  wire [63:0] regs_20_io_out; // @[RegFile.scala 66:20:@37909.4]
  wire  regs_20_io_enable; // @[RegFile.scala 66:20:@37909.4]
  wire  regs_21_clock; // @[RegFile.scala 66:20:@37923.4]
  wire  regs_21_reset; // @[RegFile.scala 66:20:@37923.4]
  wire [63:0] regs_21_io_in; // @[RegFile.scala 66:20:@37923.4]
  wire  regs_21_io_reset; // @[RegFile.scala 66:20:@37923.4]
  wire [63:0] regs_21_io_out; // @[RegFile.scala 66:20:@37923.4]
  wire  regs_21_io_enable; // @[RegFile.scala 66:20:@37923.4]
  wire  regs_22_clock; // @[RegFile.scala 66:20:@37937.4]
  wire  regs_22_reset; // @[RegFile.scala 66:20:@37937.4]
  wire [63:0] regs_22_io_in; // @[RegFile.scala 66:20:@37937.4]
  wire  regs_22_io_reset; // @[RegFile.scala 66:20:@37937.4]
  wire [63:0] regs_22_io_out; // @[RegFile.scala 66:20:@37937.4]
  wire  regs_22_io_enable; // @[RegFile.scala 66:20:@37937.4]
  wire  regs_23_clock; // @[RegFile.scala 66:20:@37951.4]
  wire  regs_23_reset; // @[RegFile.scala 66:20:@37951.4]
  wire [63:0] regs_23_io_in; // @[RegFile.scala 66:20:@37951.4]
  wire  regs_23_io_reset; // @[RegFile.scala 66:20:@37951.4]
  wire [63:0] regs_23_io_out; // @[RegFile.scala 66:20:@37951.4]
  wire  regs_23_io_enable; // @[RegFile.scala 66:20:@37951.4]
  wire  regs_24_clock; // @[RegFile.scala 66:20:@37965.4]
  wire  regs_24_reset; // @[RegFile.scala 66:20:@37965.4]
  wire [63:0] regs_24_io_in; // @[RegFile.scala 66:20:@37965.4]
  wire  regs_24_io_reset; // @[RegFile.scala 66:20:@37965.4]
  wire [63:0] regs_24_io_out; // @[RegFile.scala 66:20:@37965.4]
  wire  regs_24_io_enable; // @[RegFile.scala 66:20:@37965.4]
  wire  regs_25_clock; // @[RegFile.scala 66:20:@37979.4]
  wire  regs_25_reset; // @[RegFile.scala 66:20:@37979.4]
  wire [63:0] regs_25_io_in; // @[RegFile.scala 66:20:@37979.4]
  wire  regs_25_io_reset; // @[RegFile.scala 66:20:@37979.4]
  wire [63:0] regs_25_io_out; // @[RegFile.scala 66:20:@37979.4]
  wire  regs_25_io_enable; // @[RegFile.scala 66:20:@37979.4]
  wire  regs_26_clock; // @[RegFile.scala 66:20:@37993.4]
  wire  regs_26_reset; // @[RegFile.scala 66:20:@37993.4]
  wire [63:0] regs_26_io_in; // @[RegFile.scala 66:20:@37993.4]
  wire  regs_26_io_reset; // @[RegFile.scala 66:20:@37993.4]
  wire [63:0] regs_26_io_out; // @[RegFile.scala 66:20:@37993.4]
  wire  regs_26_io_enable; // @[RegFile.scala 66:20:@37993.4]
  wire  regs_27_clock; // @[RegFile.scala 66:20:@38007.4]
  wire  regs_27_reset; // @[RegFile.scala 66:20:@38007.4]
  wire [63:0] regs_27_io_in; // @[RegFile.scala 66:20:@38007.4]
  wire  regs_27_io_reset; // @[RegFile.scala 66:20:@38007.4]
  wire [63:0] regs_27_io_out; // @[RegFile.scala 66:20:@38007.4]
  wire  regs_27_io_enable; // @[RegFile.scala 66:20:@38007.4]
  wire  regs_28_clock; // @[RegFile.scala 66:20:@38021.4]
  wire  regs_28_reset; // @[RegFile.scala 66:20:@38021.4]
  wire [63:0] regs_28_io_in; // @[RegFile.scala 66:20:@38021.4]
  wire  regs_28_io_reset; // @[RegFile.scala 66:20:@38021.4]
  wire [63:0] regs_28_io_out; // @[RegFile.scala 66:20:@38021.4]
  wire  regs_28_io_enable; // @[RegFile.scala 66:20:@38021.4]
  wire  regs_29_clock; // @[RegFile.scala 66:20:@38035.4]
  wire  regs_29_reset; // @[RegFile.scala 66:20:@38035.4]
  wire [63:0] regs_29_io_in; // @[RegFile.scala 66:20:@38035.4]
  wire  regs_29_io_reset; // @[RegFile.scala 66:20:@38035.4]
  wire [63:0] regs_29_io_out; // @[RegFile.scala 66:20:@38035.4]
  wire  regs_29_io_enable; // @[RegFile.scala 66:20:@38035.4]
  wire  regs_30_clock; // @[RegFile.scala 66:20:@38049.4]
  wire  regs_30_reset; // @[RegFile.scala 66:20:@38049.4]
  wire [63:0] regs_30_io_in; // @[RegFile.scala 66:20:@38049.4]
  wire  regs_30_io_reset; // @[RegFile.scala 66:20:@38049.4]
  wire [63:0] regs_30_io_out; // @[RegFile.scala 66:20:@38049.4]
  wire  regs_30_io_enable; // @[RegFile.scala 66:20:@38049.4]
  wire  regs_31_clock; // @[RegFile.scala 66:20:@38063.4]
  wire  regs_31_reset; // @[RegFile.scala 66:20:@38063.4]
  wire [63:0] regs_31_io_in; // @[RegFile.scala 66:20:@38063.4]
  wire  regs_31_io_reset; // @[RegFile.scala 66:20:@38063.4]
  wire [63:0] regs_31_io_out; // @[RegFile.scala 66:20:@38063.4]
  wire  regs_31_io_enable; // @[RegFile.scala 66:20:@38063.4]
  wire  regs_32_clock; // @[RegFile.scala 66:20:@38077.4]
  wire  regs_32_reset; // @[RegFile.scala 66:20:@38077.4]
  wire [63:0] regs_32_io_in; // @[RegFile.scala 66:20:@38077.4]
  wire  regs_32_io_reset; // @[RegFile.scala 66:20:@38077.4]
  wire [63:0] regs_32_io_out; // @[RegFile.scala 66:20:@38077.4]
  wire  regs_32_io_enable; // @[RegFile.scala 66:20:@38077.4]
  wire  regs_33_clock; // @[RegFile.scala 66:20:@38091.4]
  wire  regs_33_reset; // @[RegFile.scala 66:20:@38091.4]
  wire [63:0] regs_33_io_in; // @[RegFile.scala 66:20:@38091.4]
  wire  regs_33_io_reset; // @[RegFile.scala 66:20:@38091.4]
  wire [63:0] regs_33_io_out; // @[RegFile.scala 66:20:@38091.4]
  wire  regs_33_io_enable; // @[RegFile.scala 66:20:@38091.4]
  wire  regs_34_clock; // @[RegFile.scala 66:20:@38105.4]
  wire  regs_34_reset; // @[RegFile.scala 66:20:@38105.4]
  wire [63:0] regs_34_io_in; // @[RegFile.scala 66:20:@38105.4]
  wire  regs_34_io_reset; // @[RegFile.scala 66:20:@38105.4]
  wire [63:0] regs_34_io_out; // @[RegFile.scala 66:20:@38105.4]
  wire  regs_34_io_enable; // @[RegFile.scala 66:20:@38105.4]
  wire  regs_35_clock; // @[RegFile.scala 66:20:@38119.4]
  wire  regs_35_reset; // @[RegFile.scala 66:20:@38119.4]
  wire [63:0] regs_35_io_in; // @[RegFile.scala 66:20:@38119.4]
  wire  regs_35_io_reset; // @[RegFile.scala 66:20:@38119.4]
  wire [63:0] regs_35_io_out; // @[RegFile.scala 66:20:@38119.4]
  wire  regs_35_io_enable; // @[RegFile.scala 66:20:@38119.4]
  wire  regs_36_clock; // @[RegFile.scala 66:20:@38133.4]
  wire  regs_36_reset; // @[RegFile.scala 66:20:@38133.4]
  wire [63:0] regs_36_io_in; // @[RegFile.scala 66:20:@38133.4]
  wire  regs_36_io_reset; // @[RegFile.scala 66:20:@38133.4]
  wire [63:0] regs_36_io_out; // @[RegFile.scala 66:20:@38133.4]
  wire  regs_36_io_enable; // @[RegFile.scala 66:20:@38133.4]
  wire  regs_37_clock; // @[RegFile.scala 66:20:@38147.4]
  wire  regs_37_reset; // @[RegFile.scala 66:20:@38147.4]
  wire [63:0] regs_37_io_in; // @[RegFile.scala 66:20:@38147.4]
  wire  regs_37_io_reset; // @[RegFile.scala 66:20:@38147.4]
  wire [63:0] regs_37_io_out; // @[RegFile.scala 66:20:@38147.4]
  wire  regs_37_io_enable; // @[RegFile.scala 66:20:@38147.4]
  wire  regs_38_clock; // @[RegFile.scala 66:20:@38161.4]
  wire  regs_38_reset; // @[RegFile.scala 66:20:@38161.4]
  wire [63:0] regs_38_io_in; // @[RegFile.scala 66:20:@38161.4]
  wire  regs_38_io_reset; // @[RegFile.scala 66:20:@38161.4]
  wire [63:0] regs_38_io_out; // @[RegFile.scala 66:20:@38161.4]
  wire  regs_38_io_enable; // @[RegFile.scala 66:20:@38161.4]
  wire  regs_39_clock; // @[RegFile.scala 66:20:@38175.4]
  wire  regs_39_reset; // @[RegFile.scala 66:20:@38175.4]
  wire [63:0] regs_39_io_in; // @[RegFile.scala 66:20:@38175.4]
  wire  regs_39_io_reset; // @[RegFile.scala 66:20:@38175.4]
  wire [63:0] regs_39_io_out; // @[RegFile.scala 66:20:@38175.4]
  wire  regs_39_io_enable; // @[RegFile.scala 66:20:@38175.4]
  wire  regs_40_clock; // @[RegFile.scala 66:20:@38189.4]
  wire  regs_40_reset; // @[RegFile.scala 66:20:@38189.4]
  wire [63:0] regs_40_io_in; // @[RegFile.scala 66:20:@38189.4]
  wire  regs_40_io_reset; // @[RegFile.scala 66:20:@38189.4]
  wire [63:0] regs_40_io_out; // @[RegFile.scala 66:20:@38189.4]
  wire  regs_40_io_enable; // @[RegFile.scala 66:20:@38189.4]
  wire  regs_41_clock; // @[RegFile.scala 66:20:@38203.4]
  wire  regs_41_reset; // @[RegFile.scala 66:20:@38203.4]
  wire [63:0] regs_41_io_in; // @[RegFile.scala 66:20:@38203.4]
  wire  regs_41_io_reset; // @[RegFile.scala 66:20:@38203.4]
  wire [63:0] regs_41_io_out; // @[RegFile.scala 66:20:@38203.4]
  wire  regs_41_io_enable; // @[RegFile.scala 66:20:@38203.4]
  wire  regs_42_clock; // @[RegFile.scala 66:20:@38217.4]
  wire  regs_42_reset; // @[RegFile.scala 66:20:@38217.4]
  wire [63:0] regs_42_io_in; // @[RegFile.scala 66:20:@38217.4]
  wire  regs_42_io_reset; // @[RegFile.scala 66:20:@38217.4]
  wire [63:0] regs_42_io_out; // @[RegFile.scala 66:20:@38217.4]
  wire  regs_42_io_enable; // @[RegFile.scala 66:20:@38217.4]
  wire  regs_43_clock; // @[RegFile.scala 66:20:@38231.4]
  wire  regs_43_reset; // @[RegFile.scala 66:20:@38231.4]
  wire [63:0] regs_43_io_in; // @[RegFile.scala 66:20:@38231.4]
  wire  regs_43_io_reset; // @[RegFile.scala 66:20:@38231.4]
  wire [63:0] regs_43_io_out; // @[RegFile.scala 66:20:@38231.4]
  wire  regs_43_io_enable; // @[RegFile.scala 66:20:@38231.4]
  wire  regs_44_clock; // @[RegFile.scala 66:20:@38245.4]
  wire  regs_44_reset; // @[RegFile.scala 66:20:@38245.4]
  wire [63:0] regs_44_io_in; // @[RegFile.scala 66:20:@38245.4]
  wire  regs_44_io_reset; // @[RegFile.scala 66:20:@38245.4]
  wire [63:0] regs_44_io_out; // @[RegFile.scala 66:20:@38245.4]
  wire  regs_44_io_enable; // @[RegFile.scala 66:20:@38245.4]
  wire  regs_45_clock; // @[RegFile.scala 66:20:@38259.4]
  wire  regs_45_reset; // @[RegFile.scala 66:20:@38259.4]
  wire [63:0] regs_45_io_in; // @[RegFile.scala 66:20:@38259.4]
  wire  regs_45_io_reset; // @[RegFile.scala 66:20:@38259.4]
  wire [63:0] regs_45_io_out; // @[RegFile.scala 66:20:@38259.4]
  wire  regs_45_io_enable; // @[RegFile.scala 66:20:@38259.4]
  wire  regs_46_clock; // @[RegFile.scala 66:20:@38273.4]
  wire  regs_46_reset; // @[RegFile.scala 66:20:@38273.4]
  wire [63:0] regs_46_io_in; // @[RegFile.scala 66:20:@38273.4]
  wire  regs_46_io_reset; // @[RegFile.scala 66:20:@38273.4]
  wire [63:0] regs_46_io_out; // @[RegFile.scala 66:20:@38273.4]
  wire  regs_46_io_enable; // @[RegFile.scala 66:20:@38273.4]
  wire  regs_47_clock; // @[RegFile.scala 66:20:@38287.4]
  wire  regs_47_reset; // @[RegFile.scala 66:20:@38287.4]
  wire [63:0] regs_47_io_in; // @[RegFile.scala 66:20:@38287.4]
  wire  regs_47_io_reset; // @[RegFile.scala 66:20:@38287.4]
  wire [63:0] regs_47_io_out; // @[RegFile.scala 66:20:@38287.4]
  wire  regs_47_io_enable; // @[RegFile.scala 66:20:@38287.4]
  wire  regs_48_clock; // @[RegFile.scala 66:20:@38301.4]
  wire  regs_48_reset; // @[RegFile.scala 66:20:@38301.4]
  wire [63:0] regs_48_io_in; // @[RegFile.scala 66:20:@38301.4]
  wire  regs_48_io_reset; // @[RegFile.scala 66:20:@38301.4]
  wire [63:0] regs_48_io_out; // @[RegFile.scala 66:20:@38301.4]
  wire  regs_48_io_enable; // @[RegFile.scala 66:20:@38301.4]
  wire  regs_49_clock; // @[RegFile.scala 66:20:@38315.4]
  wire  regs_49_reset; // @[RegFile.scala 66:20:@38315.4]
  wire [63:0] regs_49_io_in; // @[RegFile.scala 66:20:@38315.4]
  wire  regs_49_io_reset; // @[RegFile.scala 66:20:@38315.4]
  wire [63:0] regs_49_io_out; // @[RegFile.scala 66:20:@38315.4]
  wire  regs_49_io_enable; // @[RegFile.scala 66:20:@38315.4]
  wire  regs_50_clock; // @[RegFile.scala 66:20:@38329.4]
  wire  regs_50_reset; // @[RegFile.scala 66:20:@38329.4]
  wire [63:0] regs_50_io_in; // @[RegFile.scala 66:20:@38329.4]
  wire  regs_50_io_reset; // @[RegFile.scala 66:20:@38329.4]
  wire [63:0] regs_50_io_out; // @[RegFile.scala 66:20:@38329.4]
  wire  regs_50_io_enable; // @[RegFile.scala 66:20:@38329.4]
  wire  regs_51_clock; // @[RegFile.scala 66:20:@38343.4]
  wire  regs_51_reset; // @[RegFile.scala 66:20:@38343.4]
  wire [63:0] regs_51_io_in; // @[RegFile.scala 66:20:@38343.4]
  wire  regs_51_io_reset; // @[RegFile.scala 66:20:@38343.4]
  wire [63:0] regs_51_io_out; // @[RegFile.scala 66:20:@38343.4]
  wire  regs_51_io_enable; // @[RegFile.scala 66:20:@38343.4]
  wire  regs_52_clock; // @[RegFile.scala 66:20:@38357.4]
  wire  regs_52_reset; // @[RegFile.scala 66:20:@38357.4]
  wire [63:0] regs_52_io_in; // @[RegFile.scala 66:20:@38357.4]
  wire  regs_52_io_reset; // @[RegFile.scala 66:20:@38357.4]
  wire [63:0] regs_52_io_out; // @[RegFile.scala 66:20:@38357.4]
  wire  regs_52_io_enable; // @[RegFile.scala 66:20:@38357.4]
  wire  regs_53_clock; // @[RegFile.scala 66:20:@38371.4]
  wire  regs_53_reset; // @[RegFile.scala 66:20:@38371.4]
  wire [63:0] regs_53_io_in; // @[RegFile.scala 66:20:@38371.4]
  wire  regs_53_io_reset; // @[RegFile.scala 66:20:@38371.4]
  wire [63:0] regs_53_io_out; // @[RegFile.scala 66:20:@38371.4]
  wire  regs_53_io_enable; // @[RegFile.scala 66:20:@38371.4]
  wire  regs_54_clock; // @[RegFile.scala 66:20:@38385.4]
  wire  regs_54_reset; // @[RegFile.scala 66:20:@38385.4]
  wire [63:0] regs_54_io_in; // @[RegFile.scala 66:20:@38385.4]
  wire  regs_54_io_reset; // @[RegFile.scala 66:20:@38385.4]
  wire [63:0] regs_54_io_out; // @[RegFile.scala 66:20:@38385.4]
  wire  regs_54_io_enable; // @[RegFile.scala 66:20:@38385.4]
  wire  regs_55_clock; // @[RegFile.scala 66:20:@38399.4]
  wire  regs_55_reset; // @[RegFile.scala 66:20:@38399.4]
  wire [63:0] regs_55_io_in; // @[RegFile.scala 66:20:@38399.4]
  wire  regs_55_io_reset; // @[RegFile.scala 66:20:@38399.4]
  wire [63:0] regs_55_io_out; // @[RegFile.scala 66:20:@38399.4]
  wire  regs_55_io_enable; // @[RegFile.scala 66:20:@38399.4]
  wire  regs_56_clock; // @[RegFile.scala 66:20:@38413.4]
  wire  regs_56_reset; // @[RegFile.scala 66:20:@38413.4]
  wire [63:0] regs_56_io_in; // @[RegFile.scala 66:20:@38413.4]
  wire  regs_56_io_reset; // @[RegFile.scala 66:20:@38413.4]
  wire [63:0] regs_56_io_out; // @[RegFile.scala 66:20:@38413.4]
  wire  regs_56_io_enable; // @[RegFile.scala 66:20:@38413.4]
  wire  regs_57_clock; // @[RegFile.scala 66:20:@38427.4]
  wire  regs_57_reset; // @[RegFile.scala 66:20:@38427.4]
  wire [63:0] regs_57_io_in; // @[RegFile.scala 66:20:@38427.4]
  wire  regs_57_io_reset; // @[RegFile.scala 66:20:@38427.4]
  wire [63:0] regs_57_io_out; // @[RegFile.scala 66:20:@38427.4]
  wire  regs_57_io_enable; // @[RegFile.scala 66:20:@38427.4]
  wire  regs_58_clock; // @[RegFile.scala 66:20:@38441.4]
  wire  regs_58_reset; // @[RegFile.scala 66:20:@38441.4]
  wire [63:0] regs_58_io_in; // @[RegFile.scala 66:20:@38441.4]
  wire  regs_58_io_reset; // @[RegFile.scala 66:20:@38441.4]
  wire [63:0] regs_58_io_out; // @[RegFile.scala 66:20:@38441.4]
  wire  regs_58_io_enable; // @[RegFile.scala 66:20:@38441.4]
  wire  regs_59_clock; // @[RegFile.scala 66:20:@38455.4]
  wire  regs_59_reset; // @[RegFile.scala 66:20:@38455.4]
  wire [63:0] regs_59_io_in; // @[RegFile.scala 66:20:@38455.4]
  wire  regs_59_io_reset; // @[RegFile.scala 66:20:@38455.4]
  wire [63:0] regs_59_io_out; // @[RegFile.scala 66:20:@38455.4]
  wire  regs_59_io_enable; // @[RegFile.scala 66:20:@38455.4]
  wire  regs_60_clock; // @[RegFile.scala 66:20:@38469.4]
  wire  regs_60_reset; // @[RegFile.scala 66:20:@38469.4]
  wire [63:0] regs_60_io_in; // @[RegFile.scala 66:20:@38469.4]
  wire  regs_60_io_reset; // @[RegFile.scala 66:20:@38469.4]
  wire [63:0] regs_60_io_out; // @[RegFile.scala 66:20:@38469.4]
  wire  regs_60_io_enable; // @[RegFile.scala 66:20:@38469.4]
  wire  regs_61_clock; // @[RegFile.scala 66:20:@38483.4]
  wire  regs_61_reset; // @[RegFile.scala 66:20:@38483.4]
  wire [63:0] regs_61_io_in; // @[RegFile.scala 66:20:@38483.4]
  wire  regs_61_io_reset; // @[RegFile.scala 66:20:@38483.4]
  wire [63:0] regs_61_io_out; // @[RegFile.scala 66:20:@38483.4]
  wire  regs_61_io_enable; // @[RegFile.scala 66:20:@38483.4]
  wire  regs_62_clock; // @[RegFile.scala 66:20:@38497.4]
  wire  regs_62_reset; // @[RegFile.scala 66:20:@38497.4]
  wire [63:0] regs_62_io_in; // @[RegFile.scala 66:20:@38497.4]
  wire  regs_62_io_reset; // @[RegFile.scala 66:20:@38497.4]
  wire [63:0] regs_62_io_out; // @[RegFile.scala 66:20:@38497.4]
  wire  regs_62_io_enable; // @[RegFile.scala 66:20:@38497.4]
  wire  regs_63_clock; // @[RegFile.scala 66:20:@38511.4]
  wire  regs_63_reset; // @[RegFile.scala 66:20:@38511.4]
  wire [63:0] regs_63_io_in; // @[RegFile.scala 66:20:@38511.4]
  wire  regs_63_io_reset; // @[RegFile.scala 66:20:@38511.4]
  wire [63:0] regs_63_io_out; // @[RegFile.scala 66:20:@38511.4]
  wire  regs_63_io_enable; // @[RegFile.scala 66:20:@38511.4]
  wire  regs_64_clock; // @[RegFile.scala 66:20:@38525.4]
  wire  regs_64_reset; // @[RegFile.scala 66:20:@38525.4]
  wire [63:0] regs_64_io_in; // @[RegFile.scala 66:20:@38525.4]
  wire  regs_64_io_reset; // @[RegFile.scala 66:20:@38525.4]
  wire [63:0] regs_64_io_out; // @[RegFile.scala 66:20:@38525.4]
  wire  regs_64_io_enable; // @[RegFile.scala 66:20:@38525.4]
  wire  regs_65_clock; // @[RegFile.scala 66:20:@38539.4]
  wire  regs_65_reset; // @[RegFile.scala 66:20:@38539.4]
  wire [63:0] regs_65_io_in; // @[RegFile.scala 66:20:@38539.4]
  wire  regs_65_io_reset; // @[RegFile.scala 66:20:@38539.4]
  wire [63:0] regs_65_io_out; // @[RegFile.scala 66:20:@38539.4]
  wire  regs_65_io_enable; // @[RegFile.scala 66:20:@38539.4]
  wire  regs_66_clock; // @[RegFile.scala 66:20:@38553.4]
  wire  regs_66_reset; // @[RegFile.scala 66:20:@38553.4]
  wire [63:0] regs_66_io_in; // @[RegFile.scala 66:20:@38553.4]
  wire  regs_66_io_reset; // @[RegFile.scala 66:20:@38553.4]
  wire [63:0] regs_66_io_out; // @[RegFile.scala 66:20:@38553.4]
  wire  regs_66_io_enable; // @[RegFile.scala 66:20:@38553.4]
  wire  regs_67_clock; // @[RegFile.scala 66:20:@38567.4]
  wire  regs_67_reset; // @[RegFile.scala 66:20:@38567.4]
  wire [63:0] regs_67_io_in; // @[RegFile.scala 66:20:@38567.4]
  wire  regs_67_io_reset; // @[RegFile.scala 66:20:@38567.4]
  wire [63:0] regs_67_io_out; // @[RegFile.scala 66:20:@38567.4]
  wire  regs_67_io_enable; // @[RegFile.scala 66:20:@38567.4]
  wire  regs_68_clock; // @[RegFile.scala 66:20:@38581.4]
  wire  regs_68_reset; // @[RegFile.scala 66:20:@38581.4]
  wire [63:0] regs_68_io_in; // @[RegFile.scala 66:20:@38581.4]
  wire  regs_68_io_reset; // @[RegFile.scala 66:20:@38581.4]
  wire [63:0] regs_68_io_out; // @[RegFile.scala 66:20:@38581.4]
  wire  regs_68_io_enable; // @[RegFile.scala 66:20:@38581.4]
  wire  regs_69_clock; // @[RegFile.scala 66:20:@38595.4]
  wire  regs_69_reset; // @[RegFile.scala 66:20:@38595.4]
  wire [63:0] regs_69_io_in; // @[RegFile.scala 66:20:@38595.4]
  wire  regs_69_io_reset; // @[RegFile.scala 66:20:@38595.4]
  wire [63:0] regs_69_io_out; // @[RegFile.scala 66:20:@38595.4]
  wire  regs_69_io_enable; // @[RegFile.scala 66:20:@38595.4]
  wire  regs_70_clock; // @[RegFile.scala 66:20:@38609.4]
  wire  regs_70_reset; // @[RegFile.scala 66:20:@38609.4]
  wire [63:0] regs_70_io_in; // @[RegFile.scala 66:20:@38609.4]
  wire  regs_70_io_reset; // @[RegFile.scala 66:20:@38609.4]
  wire [63:0] regs_70_io_out; // @[RegFile.scala 66:20:@38609.4]
  wire  regs_70_io_enable; // @[RegFile.scala 66:20:@38609.4]
  wire  regs_71_clock; // @[RegFile.scala 66:20:@38623.4]
  wire  regs_71_reset; // @[RegFile.scala 66:20:@38623.4]
  wire [63:0] regs_71_io_in; // @[RegFile.scala 66:20:@38623.4]
  wire  regs_71_io_reset; // @[RegFile.scala 66:20:@38623.4]
  wire [63:0] regs_71_io_out; // @[RegFile.scala 66:20:@38623.4]
  wire  regs_71_io_enable; // @[RegFile.scala 66:20:@38623.4]
  wire  regs_72_clock; // @[RegFile.scala 66:20:@38637.4]
  wire  regs_72_reset; // @[RegFile.scala 66:20:@38637.4]
  wire [63:0] regs_72_io_in; // @[RegFile.scala 66:20:@38637.4]
  wire  regs_72_io_reset; // @[RegFile.scala 66:20:@38637.4]
  wire [63:0] regs_72_io_out; // @[RegFile.scala 66:20:@38637.4]
  wire  regs_72_io_enable; // @[RegFile.scala 66:20:@38637.4]
  wire  regs_73_clock; // @[RegFile.scala 66:20:@38651.4]
  wire  regs_73_reset; // @[RegFile.scala 66:20:@38651.4]
  wire [63:0] regs_73_io_in; // @[RegFile.scala 66:20:@38651.4]
  wire  regs_73_io_reset; // @[RegFile.scala 66:20:@38651.4]
  wire [63:0] regs_73_io_out; // @[RegFile.scala 66:20:@38651.4]
  wire  regs_73_io_enable; // @[RegFile.scala 66:20:@38651.4]
  wire  regs_74_clock; // @[RegFile.scala 66:20:@38665.4]
  wire  regs_74_reset; // @[RegFile.scala 66:20:@38665.4]
  wire [63:0] regs_74_io_in; // @[RegFile.scala 66:20:@38665.4]
  wire  regs_74_io_reset; // @[RegFile.scala 66:20:@38665.4]
  wire [63:0] regs_74_io_out; // @[RegFile.scala 66:20:@38665.4]
  wire  regs_74_io_enable; // @[RegFile.scala 66:20:@38665.4]
  wire  regs_75_clock; // @[RegFile.scala 66:20:@38679.4]
  wire  regs_75_reset; // @[RegFile.scala 66:20:@38679.4]
  wire [63:0] regs_75_io_in; // @[RegFile.scala 66:20:@38679.4]
  wire  regs_75_io_reset; // @[RegFile.scala 66:20:@38679.4]
  wire [63:0] regs_75_io_out; // @[RegFile.scala 66:20:@38679.4]
  wire  regs_75_io_enable; // @[RegFile.scala 66:20:@38679.4]
  wire  regs_76_clock; // @[RegFile.scala 66:20:@38693.4]
  wire  regs_76_reset; // @[RegFile.scala 66:20:@38693.4]
  wire [63:0] regs_76_io_in; // @[RegFile.scala 66:20:@38693.4]
  wire  regs_76_io_reset; // @[RegFile.scala 66:20:@38693.4]
  wire [63:0] regs_76_io_out; // @[RegFile.scala 66:20:@38693.4]
  wire  regs_76_io_enable; // @[RegFile.scala 66:20:@38693.4]
  wire  regs_77_clock; // @[RegFile.scala 66:20:@38707.4]
  wire  regs_77_reset; // @[RegFile.scala 66:20:@38707.4]
  wire [63:0] regs_77_io_in; // @[RegFile.scala 66:20:@38707.4]
  wire  regs_77_io_reset; // @[RegFile.scala 66:20:@38707.4]
  wire [63:0] regs_77_io_out; // @[RegFile.scala 66:20:@38707.4]
  wire  regs_77_io_enable; // @[RegFile.scala 66:20:@38707.4]
  wire  regs_78_clock; // @[RegFile.scala 66:20:@38721.4]
  wire  regs_78_reset; // @[RegFile.scala 66:20:@38721.4]
  wire [63:0] regs_78_io_in; // @[RegFile.scala 66:20:@38721.4]
  wire  regs_78_io_reset; // @[RegFile.scala 66:20:@38721.4]
  wire [63:0] regs_78_io_out; // @[RegFile.scala 66:20:@38721.4]
  wire  regs_78_io_enable; // @[RegFile.scala 66:20:@38721.4]
  wire  regs_79_clock; // @[RegFile.scala 66:20:@38735.4]
  wire  regs_79_reset; // @[RegFile.scala 66:20:@38735.4]
  wire [63:0] regs_79_io_in; // @[RegFile.scala 66:20:@38735.4]
  wire  regs_79_io_reset; // @[RegFile.scala 66:20:@38735.4]
  wire [63:0] regs_79_io_out; // @[RegFile.scala 66:20:@38735.4]
  wire  regs_79_io_enable; // @[RegFile.scala 66:20:@38735.4]
  wire  regs_80_clock; // @[RegFile.scala 66:20:@38749.4]
  wire  regs_80_reset; // @[RegFile.scala 66:20:@38749.4]
  wire [63:0] regs_80_io_in; // @[RegFile.scala 66:20:@38749.4]
  wire  regs_80_io_reset; // @[RegFile.scala 66:20:@38749.4]
  wire [63:0] regs_80_io_out; // @[RegFile.scala 66:20:@38749.4]
  wire  regs_80_io_enable; // @[RegFile.scala 66:20:@38749.4]
  wire  regs_81_clock; // @[RegFile.scala 66:20:@38763.4]
  wire  regs_81_reset; // @[RegFile.scala 66:20:@38763.4]
  wire [63:0] regs_81_io_in; // @[RegFile.scala 66:20:@38763.4]
  wire  regs_81_io_reset; // @[RegFile.scala 66:20:@38763.4]
  wire [63:0] regs_81_io_out; // @[RegFile.scala 66:20:@38763.4]
  wire  regs_81_io_enable; // @[RegFile.scala 66:20:@38763.4]
  wire  regs_82_clock; // @[RegFile.scala 66:20:@38777.4]
  wire  regs_82_reset; // @[RegFile.scala 66:20:@38777.4]
  wire [63:0] regs_82_io_in; // @[RegFile.scala 66:20:@38777.4]
  wire  regs_82_io_reset; // @[RegFile.scala 66:20:@38777.4]
  wire [63:0] regs_82_io_out; // @[RegFile.scala 66:20:@38777.4]
  wire  regs_82_io_enable; // @[RegFile.scala 66:20:@38777.4]
  wire  regs_83_clock; // @[RegFile.scala 66:20:@38791.4]
  wire  regs_83_reset; // @[RegFile.scala 66:20:@38791.4]
  wire [63:0] regs_83_io_in; // @[RegFile.scala 66:20:@38791.4]
  wire  regs_83_io_reset; // @[RegFile.scala 66:20:@38791.4]
  wire [63:0] regs_83_io_out; // @[RegFile.scala 66:20:@38791.4]
  wire  regs_83_io_enable; // @[RegFile.scala 66:20:@38791.4]
  wire  regs_84_clock; // @[RegFile.scala 66:20:@38805.4]
  wire  regs_84_reset; // @[RegFile.scala 66:20:@38805.4]
  wire [63:0] regs_84_io_in; // @[RegFile.scala 66:20:@38805.4]
  wire  regs_84_io_reset; // @[RegFile.scala 66:20:@38805.4]
  wire [63:0] regs_84_io_out; // @[RegFile.scala 66:20:@38805.4]
  wire  regs_84_io_enable; // @[RegFile.scala 66:20:@38805.4]
  wire  regs_85_clock; // @[RegFile.scala 66:20:@38819.4]
  wire  regs_85_reset; // @[RegFile.scala 66:20:@38819.4]
  wire [63:0] regs_85_io_in; // @[RegFile.scala 66:20:@38819.4]
  wire  regs_85_io_reset; // @[RegFile.scala 66:20:@38819.4]
  wire [63:0] regs_85_io_out; // @[RegFile.scala 66:20:@38819.4]
  wire  regs_85_io_enable; // @[RegFile.scala 66:20:@38819.4]
  wire  regs_86_clock; // @[RegFile.scala 66:20:@38833.4]
  wire  regs_86_reset; // @[RegFile.scala 66:20:@38833.4]
  wire [63:0] regs_86_io_in; // @[RegFile.scala 66:20:@38833.4]
  wire  regs_86_io_reset; // @[RegFile.scala 66:20:@38833.4]
  wire [63:0] regs_86_io_out; // @[RegFile.scala 66:20:@38833.4]
  wire  regs_86_io_enable; // @[RegFile.scala 66:20:@38833.4]
  wire  regs_87_clock; // @[RegFile.scala 66:20:@38847.4]
  wire  regs_87_reset; // @[RegFile.scala 66:20:@38847.4]
  wire [63:0] regs_87_io_in; // @[RegFile.scala 66:20:@38847.4]
  wire  regs_87_io_reset; // @[RegFile.scala 66:20:@38847.4]
  wire [63:0] regs_87_io_out; // @[RegFile.scala 66:20:@38847.4]
  wire  regs_87_io_enable; // @[RegFile.scala 66:20:@38847.4]
  wire  regs_88_clock; // @[RegFile.scala 66:20:@38861.4]
  wire  regs_88_reset; // @[RegFile.scala 66:20:@38861.4]
  wire [63:0] regs_88_io_in; // @[RegFile.scala 66:20:@38861.4]
  wire  regs_88_io_reset; // @[RegFile.scala 66:20:@38861.4]
  wire [63:0] regs_88_io_out; // @[RegFile.scala 66:20:@38861.4]
  wire  regs_88_io_enable; // @[RegFile.scala 66:20:@38861.4]
  wire  regs_89_clock; // @[RegFile.scala 66:20:@38875.4]
  wire  regs_89_reset; // @[RegFile.scala 66:20:@38875.4]
  wire [63:0] regs_89_io_in; // @[RegFile.scala 66:20:@38875.4]
  wire  regs_89_io_reset; // @[RegFile.scala 66:20:@38875.4]
  wire [63:0] regs_89_io_out; // @[RegFile.scala 66:20:@38875.4]
  wire  regs_89_io_enable; // @[RegFile.scala 66:20:@38875.4]
  wire  regs_90_clock; // @[RegFile.scala 66:20:@38889.4]
  wire  regs_90_reset; // @[RegFile.scala 66:20:@38889.4]
  wire [63:0] regs_90_io_in; // @[RegFile.scala 66:20:@38889.4]
  wire  regs_90_io_reset; // @[RegFile.scala 66:20:@38889.4]
  wire [63:0] regs_90_io_out; // @[RegFile.scala 66:20:@38889.4]
  wire  regs_90_io_enable; // @[RegFile.scala 66:20:@38889.4]
  wire  regs_91_clock; // @[RegFile.scala 66:20:@38903.4]
  wire  regs_91_reset; // @[RegFile.scala 66:20:@38903.4]
  wire [63:0] regs_91_io_in; // @[RegFile.scala 66:20:@38903.4]
  wire  regs_91_io_reset; // @[RegFile.scala 66:20:@38903.4]
  wire [63:0] regs_91_io_out; // @[RegFile.scala 66:20:@38903.4]
  wire  regs_91_io_enable; // @[RegFile.scala 66:20:@38903.4]
  wire  regs_92_clock; // @[RegFile.scala 66:20:@38917.4]
  wire  regs_92_reset; // @[RegFile.scala 66:20:@38917.4]
  wire [63:0] regs_92_io_in; // @[RegFile.scala 66:20:@38917.4]
  wire  regs_92_io_reset; // @[RegFile.scala 66:20:@38917.4]
  wire [63:0] regs_92_io_out; // @[RegFile.scala 66:20:@38917.4]
  wire  regs_92_io_enable; // @[RegFile.scala 66:20:@38917.4]
  wire  regs_93_clock; // @[RegFile.scala 66:20:@38931.4]
  wire  regs_93_reset; // @[RegFile.scala 66:20:@38931.4]
  wire [63:0] regs_93_io_in; // @[RegFile.scala 66:20:@38931.4]
  wire  regs_93_io_reset; // @[RegFile.scala 66:20:@38931.4]
  wire [63:0] regs_93_io_out; // @[RegFile.scala 66:20:@38931.4]
  wire  regs_93_io_enable; // @[RegFile.scala 66:20:@38931.4]
  wire  regs_94_clock; // @[RegFile.scala 66:20:@38945.4]
  wire  regs_94_reset; // @[RegFile.scala 66:20:@38945.4]
  wire [63:0] regs_94_io_in; // @[RegFile.scala 66:20:@38945.4]
  wire  regs_94_io_reset; // @[RegFile.scala 66:20:@38945.4]
  wire [63:0] regs_94_io_out; // @[RegFile.scala 66:20:@38945.4]
  wire  regs_94_io_enable; // @[RegFile.scala 66:20:@38945.4]
  wire  regs_95_clock; // @[RegFile.scala 66:20:@38959.4]
  wire  regs_95_reset; // @[RegFile.scala 66:20:@38959.4]
  wire [63:0] regs_95_io_in; // @[RegFile.scala 66:20:@38959.4]
  wire  regs_95_io_reset; // @[RegFile.scala 66:20:@38959.4]
  wire [63:0] regs_95_io_out; // @[RegFile.scala 66:20:@38959.4]
  wire  regs_95_io_enable; // @[RegFile.scala 66:20:@38959.4]
  wire  regs_96_clock; // @[RegFile.scala 66:20:@38973.4]
  wire  regs_96_reset; // @[RegFile.scala 66:20:@38973.4]
  wire [63:0] regs_96_io_in; // @[RegFile.scala 66:20:@38973.4]
  wire  regs_96_io_reset; // @[RegFile.scala 66:20:@38973.4]
  wire [63:0] regs_96_io_out; // @[RegFile.scala 66:20:@38973.4]
  wire  regs_96_io_enable; // @[RegFile.scala 66:20:@38973.4]
  wire  regs_97_clock; // @[RegFile.scala 66:20:@38987.4]
  wire  regs_97_reset; // @[RegFile.scala 66:20:@38987.4]
  wire [63:0] regs_97_io_in; // @[RegFile.scala 66:20:@38987.4]
  wire  regs_97_io_reset; // @[RegFile.scala 66:20:@38987.4]
  wire [63:0] regs_97_io_out; // @[RegFile.scala 66:20:@38987.4]
  wire  regs_97_io_enable; // @[RegFile.scala 66:20:@38987.4]
  wire  regs_98_clock; // @[RegFile.scala 66:20:@39001.4]
  wire  regs_98_reset; // @[RegFile.scala 66:20:@39001.4]
  wire [63:0] regs_98_io_in; // @[RegFile.scala 66:20:@39001.4]
  wire  regs_98_io_reset; // @[RegFile.scala 66:20:@39001.4]
  wire [63:0] regs_98_io_out; // @[RegFile.scala 66:20:@39001.4]
  wire  regs_98_io_enable; // @[RegFile.scala 66:20:@39001.4]
  wire  regs_99_clock; // @[RegFile.scala 66:20:@39015.4]
  wire  regs_99_reset; // @[RegFile.scala 66:20:@39015.4]
  wire [63:0] regs_99_io_in; // @[RegFile.scala 66:20:@39015.4]
  wire  regs_99_io_reset; // @[RegFile.scala 66:20:@39015.4]
  wire [63:0] regs_99_io_out; // @[RegFile.scala 66:20:@39015.4]
  wire  regs_99_io_enable; // @[RegFile.scala 66:20:@39015.4]
  wire  regs_100_clock; // @[RegFile.scala 66:20:@39029.4]
  wire  regs_100_reset; // @[RegFile.scala 66:20:@39029.4]
  wire [63:0] regs_100_io_in; // @[RegFile.scala 66:20:@39029.4]
  wire  regs_100_io_reset; // @[RegFile.scala 66:20:@39029.4]
  wire [63:0] regs_100_io_out; // @[RegFile.scala 66:20:@39029.4]
  wire  regs_100_io_enable; // @[RegFile.scala 66:20:@39029.4]
  wire  regs_101_clock; // @[RegFile.scala 66:20:@39043.4]
  wire  regs_101_reset; // @[RegFile.scala 66:20:@39043.4]
  wire [63:0] regs_101_io_in; // @[RegFile.scala 66:20:@39043.4]
  wire  regs_101_io_reset; // @[RegFile.scala 66:20:@39043.4]
  wire [63:0] regs_101_io_out; // @[RegFile.scala 66:20:@39043.4]
  wire  regs_101_io_enable; // @[RegFile.scala 66:20:@39043.4]
  wire  regs_102_clock; // @[RegFile.scala 66:20:@39057.4]
  wire  regs_102_reset; // @[RegFile.scala 66:20:@39057.4]
  wire [63:0] regs_102_io_in; // @[RegFile.scala 66:20:@39057.4]
  wire  regs_102_io_reset; // @[RegFile.scala 66:20:@39057.4]
  wire [63:0] regs_102_io_out; // @[RegFile.scala 66:20:@39057.4]
  wire  regs_102_io_enable; // @[RegFile.scala 66:20:@39057.4]
  wire  regs_103_clock; // @[RegFile.scala 66:20:@39071.4]
  wire  regs_103_reset; // @[RegFile.scala 66:20:@39071.4]
  wire [63:0] regs_103_io_in; // @[RegFile.scala 66:20:@39071.4]
  wire  regs_103_io_reset; // @[RegFile.scala 66:20:@39071.4]
  wire [63:0] regs_103_io_out; // @[RegFile.scala 66:20:@39071.4]
  wire  regs_103_io_enable; // @[RegFile.scala 66:20:@39071.4]
  wire  regs_104_clock; // @[RegFile.scala 66:20:@39085.4]
  wire  regs_104_reset; // @[RegFile.scala 66:20:@39085.4]
  wire [63:0] regs_104_io_in; // @[RegFile.scala 66:20:@39085.4]
  wire  regs_104_io_reset; // @[RegFile.scala 66:20:@39085.4]
  wire [63:0] regs_104_io_out; // @[RegFile.scala 66:20:@39085.4]
  wire  regs_104_io_enable; // @[RegFile.scala 66:20:@39085.4]
  wire  regs_105_clock; // @[RegFile.scala 66:20:@39099.4]
  wire  regs_105_reset; // @[RegFile.scala 66:20:@39099.4]
  wire [63:0] regs_105_io_in; // @[RegFile.scala 66:20:@39099.4]
  wire  regs_105_io_reset; // @[RegFile.scala 66:20:@39099.4]
  wire [63:0] regs_105_io_out; // @[RegFile.scala 66:20:@39099.4]
  wire  regs_105_io_enable; // @[RegFile.scala 66:20:@39099.4]
  wire  regs_106_clock; // @[RegFile.scala 66:20:@39113.4]
  wire  regs_106_reset; // @[RegFile.scala 66:20:@39113.4]
  wire [63:0] regs_106_io_in; // @[RegFile.scala 66:20:@39113.4]
  wire  regs_106_io_reset; // @[RegFile.scala 66:20:@39113.4]
  wire [63:0] regs_106_io_out; // @[RegFile.scala 66:20:@39113.4]
  wire  regs_106_io_enable; // @[RegFile.scala 66:20:@39113.4]
  wire  regs_107_clock; // @[RegFile.scala 66:20:@39127.4]
  wire  regs_107_reset; // @[RegFile.scala 66:20:@39127.4]
  wire [63:0] regs_107_io_in; // @[RegFile.scala 66:20:@39127.4]
  wire  regs_107_io_reset; // @[RegFile.scala 66:20:@39127.4]
  wire [63:0] regs_107_io_out; // @[RegFile.scala 66:20:@39127.4]
  wire  regs_107_io_enable; // @[RegFile.scala 66:20:@39127.4]
  wire  regs_108_clock; // @[RegFile.scala 66:20:@39141.4]
  wire  regs_108_reset; // @[RegFile.scala 66:20:@39141.4]
  wire [63:0] regs_108_io_in; // @[RegFile.scala 66:20:@39141.4]
  wire  regs_108_io_reset; // @[RegFile.scala 66:20:@39141.4]
  wire [63:0] regs_108_io_out; // @[RegFile.scala 66:20:@39141.4]
  wire  regs_108_io_enable; // @[RegFile.scala 66:20:@39141.4]
  wire  regs_109_clock; // @[RegFile.scala 66:20:@39155.4]
  wire  regs_109_reset; // @[RegFile.scala 66:20:@39155.4]
  wire [63:0] regs_109_io_in; // @[RegFile.scala 66:20:@39155.4]
  wire  regs_109_io_reset; // @[RegFile.scala 66:20:@39155.4]
  wire [63:0] regs_109_io_out; // @[RegFile.scala 66:20:@39155.4]
  wire  regs_109_io_enable; // @[RegFile.scala 66:20:@39155.4]
  wire  regs_110_clock; // @[RegFile.scala 66:20:@39169.4]
  wire  regs_110_reset; // @[RegFile.scala 66:20:@39169.4]
  wire [63:0] regs_110_io_in; // @[RegFile.scala 66:20:@39169.4]
  wire  regs_110_io_reset; // @[RegFile.scala 66:20:@39169.4]
  wire [63:0] regs_110_io_out; // @[RegFile.scala 66:20:@39169.4]
  wire  regs_110_io_enable; // @[RegFile.scala 66:20:@39169.4]
  wire  regs_111_clock; // @[RegFile.scala 66:20:@39183.4]
  wire  regs_111_reset; // @[RegFile.scala 66:20:@39183.4]
  wire [63:0] regs_111_io_in; // @[RegFile.scala 66:20:@39183.4]
  wire  regs_111_io_reset; // @[RegFile.scala 66:20:@39183.4]
  wire [63:0] regs_111_io_out; // @[RegFile.scala 66:20:@39183.4]
  wire  regs_111_io_enable; // @[RegFile.scala 66:20:@39183.4]
  wire  regs_112_clock; // @[RegFile.scala 66:20:@39197.4]
  wire  regs_112_reset; // @[RegFile.scala 66:20:@39197.4]
  wire [63:0] regs_112_io_in; // @[RegFile.scala 66:20:@39197.4]
  wire  regs_112_io_reset; // @[RegFile.scala 66:20:@39197.4]
  wire [63:0] regs_112_io_out; // @[RegFile.scala 66:20:@39197.4]
  wire  regs_112_io_enable; // @[RegFile.scala 66:20:@39197.4]
  wire  regs_113_clock; // @[RegFile.scala 66:20:@39211.4]
  wire  regs_113_reset; // @[RegFile.scala 66:20:@39211.4]
  wire [63:0] regs_113_io_in; // @[RegFile.scala 66:20:@39211.4]
  wire  regs_113_io_reset; // @[RegFile.scala 66:20:@39211.4]
  wire [63:0] regs_113_io_out; // @[RegFile.scala 66:20:@39211.4]
  wire  regs_113_io_enable; // @[RegFile.scala 66:20:@39211.4]
  wire  regs_114_clock; // @[RegFile.scala 66:20:@39225.4]
  wire  regs_114_reset; // @[RegFile.scala 66:20:@39225.4]
  wire [63:0] regs_114_io_in; // @[RegFile.scala 66:20:@39225.4]
  wire  regs_114_io_reset; // @[RegFile.scala 66:20:@39225.4]
  wire [63:0] regs_114_io_out; // @[RegFile.scala 66:20:@39225.4]
  wire  regs_114_io_enable; // @[RegFile.scala 66:20:@39225.4]
  wire  regs_115_clock; // @[RegFile.scala 66:20:@39239.4]
  wire  regs_115_reset; // @[RegFile.scala 66:20:@39239.4]
  wire [63:0] regs_115_io_in; // @[RegFile.scala 66:20:@39239.4]
  wire  regs_115_io_reset; // @[RegFile.scala 66:20:@39239.4]
  wire [63:0] regs_115_io_out; // @[RegFile.scala 66:20:@39239.4]
  wire  regs_115_io_enable; // @[RegFile.scala 66:20:@39239.4]
  wire  regs_116_clock; // @[RegFile.scala 66:20:@39253.4]
  wire  regs_116_reset; // @[RegFile.scala 66:20:@39253.4]
  wire [63:0] regs_116_io_in; // @[RegFile.scala 66:20:@39253.4]
  wire  regs_116_io_reset; // @[RegFile.scala 66:20:@39253.4]
  wire [63:0] regs_116_io_out; // @[RegFile.scala 66:20:@39253.4]
  wire  regs_116_io_enable; // @[RegFile.scala 66:20:@39253.4]
  wire  regs_117_clock; // @[RegFile.scala 66:20:@39267.4]
  wire  regs_117_reset; // @[RegFile.scala 66:20:@39267.4]
  wire [63:0] regs_117_io_in; // @[RegFile.scala 66:20:@39267.4]
  wire  regs_117_io_reset; // @[RegFile.scala 66:20:@39267.4]
  wire [63:0] regs_117_io_out; // @[RegFile.scala 66:20:@39267.4]
  wire  regs_117_io_enable; // @[RegFile.scala 66:20:@39267.4]
  wire  regs_118_clock; // @[RegFile.scala 66:20:@39281.4]
  wire  regs_118_reset; // @[RegFile.scala 66:20:@39281.4]
  wire [63:0] regs_118_io_in; // @[RegFile.scala 66:20:@39281.4]
  wire  regs_118_io_reset; // @[RegFile.scala 66:20:@39281.4]
  wire [63:0] regs_118_io_out; // @[RegFile.scala 66:20:@39281.4]
  wire  regs_118_io_enable; // @[RegFile.scala 66:20:@39281.4]
  wire  regs_119_clock; // @[RegFile.scala 66:20:@39295.4]
  wire  regs_119_reset; // @[RegFile.scala 66:20:@39295.4]
  wire [63:0] regs_119_io_in; // @[RegFile.scala 66:20:@39295.4]
  wire  regs_119_io_reset; // @[RegFile.scala 66:20:@39295.4]
  wire [63:0] regs_119_io_out; // @[RegFile.scala 66:20:@39295.4]
  wire  regs_119_io_enable; // @[RegFile.scala 66:20:@39295.4]
  wire  regs_120_clock; // @[RegFile.scala 66:20:@39309.4]
  wire  regs_120_reset; // @[RegFile.scala 66:20:@39309.4]
  wire [63:0] regs_120_io_in; // @[RegFile.scala 66:20:@39309.4]
  wire  regs_120_io_reset; // @[RegFile.scala 66:20:@39309.4]
  wire [63:0] regs_120_io_out; // @[RegFile.scala 66:20:@39309.4]
  wire  regs_120_io_enable; // @[RegFile.scala 66:20:@39309.4]
  wire  regs_121_clock; // @[RegFile.scala 66:20:@39323.4]
  wire  regs_121_reset; // @[RegFile.scala 66:20:@39323.4]
  wire [63:0] regs_121_io_in; // @[RegFile.scala 66:20:@39323.4]
  wire  regs_121_io_reset; // @[RegFile.scala 66:20:@39323.4]
  wire [63:0] regs_121_io_out; // @[RegFile.scala 66:20:@39323.4]
  wire  regs_121_io_enable; // @[RegFile.scala 66:20:@39323.4]
  wire  regs_122_clock; // @[RegFile.scala 66:20:@39337.4]
  wire  regs_122_reset; // @[RegFile.scala 66:20:@39337.4]
  wire [63:0] regs_122_io_in; // @[RegFile.scala 66:20:@39337.4]
  wire  regs_122_io_reset; // @[RegFile.scala 66:20:@39337.4]
  wire [63:0] regs_122_io_out; // @[RegFile.scala 66:20:@39337.4]
  wire  regs_122_io_enable; // @[RegFile.scala 66:20:@39337.4]
  wire  regs_123_clock; // @[RegFile.scala 66:20:@39351.4]
  wire  regs_123_reset; // @[RegFile.scala 66:20:@39351.4]
  wire [63:0] regs_123_io_in; // @[RegFile.scala 66:20:@39351.4]
  wire  regs_123_io_reset; // @[RegFile.scala 66:20:@39351.4]
  wire [63:0] regs_123_io_out; // @[RegFile.scala 66:20:@39351.4]
  wire  regs_123_io_enable; // @[RegFile.scala 66:20:@39351.4]
  wire  regs_124_clock; // @[RegFile.scala 66:20:@39365.4]
  wire  regs_124_reset; // @[RegFile.scala 66:20:@39365.4]
  wire [63:0] regs_124_io_in; // @[RegFile.scala 66:20:@39365.4]
  wire  regs_124_io_reset; // @[RegFile.scala 66:20:@39365.4]
  wire [63:0] regs_124_io_out; // @[RegFile.scala 66:20:@39365.4]
  wire  regs_124_io_enable; // @[RegFile.scala 66:20:@39365.4]
  wire  regs_125_clock; // @[RegFile.scala 66:20:@39379.4]
  wire  regs_125_reset; // @[RegFile.scala 66:20:@39379.4]
  wire [63:0] regs_125_io_in; // @[RegFile.scala 66:20:@39379.4]
  wire  regs_125_io_reset; // @[RegFile.scala 66:20:@39379.4]
  wire [63:0] regs_125_io_out; // @[RegFile.scala 66:20:@39379.4]
  wire  regs_125_io_enable; // @[RegFile.scala 66:20:@39379.4]
  wire  regs_126_clock; // @[RegFile.scala 66:20:@39393.4]
  wire  regs_126_reset; // @[RegFile.scala 66:20:@39393.4]
  wire [63:0] regs_126_io_in; // @[RegFile.scala 66:20:@39393.4]
  wire  regs_126_io_reset; // @[RegFile.scala 66:20:@39393.4]
  wire [63:0] regs_126_io_out; // @[RegFile.scala 66:20:@39393.4]
  wire  regs_126_io_enable; // @[RegFile.scala 66:20:@39393.4]
  wire  regs_127_clock; // @[RegFile.scala 66:20:@39407.4]
  wire  regs_127_reset; // @[RegFile.scala 66:20:@39407.4]
  wire [63:0] regs_127_io_in; // @[RegFile.scala 66:20:@39407.4]
  wire  regs_127_io_reset; // @[RegFile.scala 66:20:@39407.4]
  wire [63:0] regs_127_io_out; // @[RegFile.scala 66:20:@39407.4]
  wire  regs_127_io_enable; // @[RegFile.scala 66:20:@39407.4]
  wire  regs_128_clock; // @[RegFile.scala 66:20:@39421.4]
  wire  regs_128_reset; // @[RegFile.scala 66:20:@39421.4]
  wire [63:0] regs_128_io_in; // @[RegFile.scala 66:20:@39421.4]
  wire  regs_128_io_reset; // @[RegFile.scala 66:20:@39421.4]
  wire [63:0] regs_128_io_out; // @[RegFile.scala 66:20:@39421.4]
  wire  regs_128_io_enable; // @[RegFile.scala 66:20:@39421.4]
  wire  regs_129_clock; // @[RegFile.scala 66:20:@39435.4]
  wire  regs_129_reset; // @[RegFile.scala 66:20:@39435.4]
  wire [63:0] regs_129_io_in; // @[RegFile.scala 66:20:@39435.4]
  wire  regs_129_io_reset; // @[RegFile.scala 66:20:@39435.4]
  wire [63:0] regs_129_io_out; // @[RegFile.scala 66:20:@39435.4]
  wire  regs_129_io_enable; // @[RegFile.scala 66:20:@39435.4]
  wire  regs_130_clock; // @[RegFile.scala 66:20:@39449.4]
  wire  regs_130_reset; // @[RegFile.scala 66:20:@39449.4]
  wire [63:0] regs_130_io_in; // @[RegFile.scala 66:20:@39449.4]
  wire  regs_130_io_reset; // @[RegFile.scala 66:20:@39449.4]
  wire [63:0] regs_130_io_out; // @[RegFile.scala 66:20:@39449.4]
  wire  regs_130_io_enable; // @[RegFile.scala 66:20:@39449.4]
  wire  regs_131_clock; // @[RegFile.scala 66:20:@39463.4]
  wire  regs_131_reset; // @[RegFile.scala 66:20:@39463.4]
  wire [63:0] regs_131_io_in; // @[RegFile.scala 66:20:@39463.4]
  wire  regs_131_io_reset; // @[RegFile.scala 66:20:@39463.4]
  wire [63:0] regs_131_io_out; // @[RegFile.scala 66:20:@39463.4]
  wire  regs_131_io_enable; // @[RegFile.scala 66:20:@39463.4]
  wire  regs_132_clock; // @[RegFile.scala 66:20:@39477.4]
  wire  regs_132_reset; // @[RegFile.scala 66:20:@39477.4]
  wire [63:0] regs_132_io_in; // @[RegFile.scala 66:20:@39477.4]
  wire  regs_132_io_reset; // @[RegFile.scala 66:20:@39477.4]
  wire [63:0] regs_132_io_out; // @[RegFile.scala 66:20:@39477.4]
  wire  regs_132_io_enable; // @[RegFile.scala 66:20:@39477.4]
  wire  regs_133_clock; // @[RegFile.scala 66:20:@39491.4]
  wire  regs_133_reset; // @[RegFile.scala 66:20:@39491.4]
  wire [63:0] regs_133_io_in; // @[RegFile.scala 66:20:@39491.4]
  wire  regs_133_io_reset; // @[RegFile.scala 66:20:@39491.4]
  wire [63:0] regs_133_io_out; // @[RegFile.scala 66:20:@39491.4]
  wire  regs_133_io_enable; // @[RegFile.scala 66:20:@39491.4]
  wire  regs_134_clock; // @[RegFile.scala 66:20:@39505.4]
  wire  regs_134_reset; // @[RegFile.scala 66:20:@39505.4]
  wire [63:0] regs_134_io_in; // @[RegFile.scala 66:20:@39505.4]
  wire  regs_134_io_reset; // @[RegFile.scala 66:20:@39505.4]
  wire [63:0] regs_134_io_out; // @[RegFile.scala 66:20:@39505.4]
  wire  regs_134_io_enable; // @[RegFile.scala 66:20:@39505.4]
  wire  regs_135_clock; // @[RegFile.scala 66:20:@39519.4]
  wire  regs_135_reset; // @[RegFile.scala 66:20:@39519.4]
  wire [63:0] regs_135_io_in; // @[RegFile.scala 66:20:@39519.4]
  wire  regs_135_io_reset; // @[RegFile.scala 66:20:@39519.4]
  wire [63:0] regs_135_io_out; // @[RegFile.scala 66:20:@39519.4]
  wire  regs_135_io_enable; // @[RegFile.scala 66:20:@39519.4]
  wire  regs_136_clock; // @[RegFile.scala 66:20:@39533.4]
  wire  regs_136_reset; // @[RegFile.scala 66:20:@39533.4]
  wire [63:0] regs_136_io_in; // @[RegFile.scala 66:20:@39533.4]
  wire  regs_136_io_reset; // @[RegFile.scala 66:20:@39533.4]
  wire [63:0] regs_136_io_out; // @[RegFile.scala 66:20:@39533.4]
  wire  regs_136_io_enable; // @[RegFile.scala 66:20:@39533.4]
  wire  regs_137_clock; // @[RegFile.scala 66:20:@39547.4]
  wire  regs_137_reset; // @[RegFile.scala 66:20:@39547.4]
  wire [63:0] regs_137_io_in; // @[RegFile.scala 66:20:@39547.4]
  wire  regs_137_io_reset; // @[RegFile.scala 66:20:@39547.4]
  wire [63:0] regs_137_io_out; // @[RegFile.scala 66:20:@39547.4]
  wire  regs_137_io_enable; // @[RegFile.scala 66:20:@39547.4]
  wire  regs_138_clock; // @[RegFile.scala 66:20:@39561.4]
  wire  regs_138_reset; // @[RegFile.scala 66:20:@39561.4]
  wire [63:0] regs_138_io_in; // @[RegFile.scala 66:20:@39561.4]
  wire  regs_138_io_reset; // @[RegFile.scala 66:20:@39561.4]
  wire [63:0] regs_138_io_out; // @[RegFile.scala 66:20:@39561.4]
  wire  regs_138_io_enable; // @[RegFile.scala 66:20:@39561.4]
  wire  regs_139_clock; // @[RegFile.scala 66:20:@39575.4]
  wire  regs_139_reset; // @[RegFile.scala 66:20:@39575.4]
  wire [63:0] regs_139_io_in; // @[RegFile.scala 66:20:@39575.4]
  wire  regs_139_io_reset; // @[RegFile.scala 66:20:@39575.4]
  wire [63:0] regs_139_io_out; // @[RegFile.scala 66:20:@39575.4]
  wire  regs_139_io_enable; // @[RegFile.scala 66:20:@39575.4]
  wire  regs_140_clock; // @[RegFile.scala 66:20:@39589.4]
  wire  regs_140_reset; // @[RegFile.scala 66:20:@39589.4]
  wire [63:0] regs_140_io_in; // @[RegFile.scala 66:20:@39589.4]
  wire  regs_140_io_reset; // @[RegFile.scala 66:20:@39589.4]
  wire [63:0] regs_140_io_out; // @[RegFile.scala 66:20:@39589.4]
  wire  regs_140_io_enable; // @[RegFile.scala 66:20:@39589.4]
  wire  regs_141_clock; // @[RegFile.scala 66:20:@39603.4]
  wire  regs_141_reset; // @[RegFile.scala 66:20:@39603.4]
  wire [63:0] regs_141_io_in; // @[RegFile.scala 66:20:@39603.4]
  wire  regs_141_io_reset; // @[RegFile.scala 66:20:@39603.4]
  wire [63:0] regs_141_io_out; // @[RegFile.scala 66:20:@39603.4]
  wire  regs_141_io_enable; // @[RegFile.scala 66:20:@39603.4]
  wire  regs_142_clock; // @[RegFile.scala 66:20:@39617.4]
  wire  regs_142_reset; // @[RegFile.scala 66:20:@39617.4]
  wire [63:0] regs_142_io_in; // @[RegFile.scala 66:20:@39617.4]
  wire  regs_142_io_reset; // @[RegFile.scala 66:20:@39617.4]
  wire [63:0] regs_142_io_out; // @[RegFile.scala 66:20:@39617.4]
  wire  regs_142_io_enable; // @[RegFile.scala 66:20:@39617.4]
  wire  regs_143_clock; // @[RegFile.scala 66:20:@39631.4]
  wire  regs_143_reset; // @[RegFile.scala 66:20:@39631.4]
  wire [63:0] regs_143_io_in; // @[RegFile.scala 66:20:@39631.4]
  wire  regs_143_io_reset; // @[RegFile.scala 66:20:@39631.4]
  wire [63:0] regs_143_io_out; // @[RegFile.scala 66:20:@39631.4]
  wire  regs_143_io_enable; // @[RegFile.scala 66:20:@39631.4]
  wire  regs_144_clock; // @[RegFile.scala 66:20:@39645.4]
  wire  regs_144_reset; // @[RegFile.scala 66:20:@39645.4]
  wire [63:0] regs_144_io_in; // @[RegFile.scala 66:20:@39645.4]
  wire  regs_144_io_reset; // @[RegFile.scala 66:20:@39645.4]
  wire [63:0] regs_144_io_out; // @[RegFile.scala 66:20:@39645.4]
  wire  regs_144_io_enable; // @[RegFile.scala 66:20:@39645.4]
  wire  regs_145_clock; // @[RegFile.scala 66:20:@39659.4]
  wire  regs_145_reset; // @[RegFile.scala 66:20:@39659.4]
  wire [63:0] regs_145_io_in; // @[RegFile.scala 66:20:@39659.4]
  wire  regs_145_io_reset; // @[RegFile.scala 66:20:@39659.4]
  wire [63:0] regs_145_io_out; // @[RegFile.scala 66:20:@39659.4]
  wire  regs_145_io_enable; // @[RegFile.scala 66:20:@39659.4]
  wire  regs_146_clock; // @[RegFile.scala 66:20:@39673.4]
  wire  regs_146_reset; // @[RegFile.scala 66:20:@39673.4]
  wire [63:0] regs_146_io_in; // @[RegFile.scala 66:20:@39673.4]
  wire  regs_146_io_reset; // @[RegFile.scala 66:20:@39673.4]
  wire [63:0] regs_146_io_out; // @[RegFile.scala 66:20:@39673.4]
  wire  regs_146_io_enable; // @[RegFile.scala 66:20:@39673.4]
  wire  regs_147_clock; // @[RegFile.scala 66:20:@39687.4]
  wire  regs_147_reset; // @[RegFile.scala 66:20:@39687.4]
  wire [63:0] regs_147_io_in; // @[RegFile.scala 66:20:@39687.4]
  wire  regs_147_io_reset; // @[RegFile.scala 66:20:@39687.4]
  wire [63:0] regs_147_io_out; // @[RegFile.scala 66:20:@39687.4]
  wire  regs_147_io_enable; // @[RegFile.scala 66:20:@39687.4]
  wire  regs_148_clock; // @[RegFile.scala 66:20:@39701.4]
  wire  regs_148_reset; // @[RegFile.scala 66:20:@39701.4]
  wire [63:0] regs_148_io_in; // @[RegFile.scala 66:20:@39701.4]
  wire  regs_148_io_reset; // @[RegFile.scala 66:20:@39701.4]
  wire [63:0] regs_148_io_out; // @[RegFile.scala 66:20:@39701.4]
  wire  regs_148_io_enable; // @[RegFile.scala 66:20:@39701.4]
  wire  regs_149_clock; // @[RegFile.scala 66:20:@39715.4]
  wire  regs_149_reset; // @[RegFile.scala 66:20:@39715.4]
  wire [63:0] regs_149_io_in; // @[RegFile.scala 66:20:@39715.4]
  wire  regs_149_io_reset; // @[RegFile.scala 66:20:@39715.4]
  wire [63:0] regs_149_io_out; // @[RegFile.scala 66:20:@39715.4]
  wire  regs_149_io_enable; // @[RegFile.scala 66:20:@39715.4]
  wire  regs_150_clock; // @[RegFile.scala 66:20:@39729.4]
  wire  regs_150_reset; // @[RegFile.scala 66:20:@39729.4]
  wire [63:0] regs_150_io_in; // @[RegFile.scala 66:20:@39729.4]
  wire  regs_150_io_reset; // @[RegFile.scala 66:20:@39729.4]
  wire [63:0] regs_150_io_out; // @[RegFile.scala 66:20:@39729.4]
  wire  regs_150_io_enable; // @[RegFile.scala 66:20:@39729.4]
  wire  regs_151_clock; // @[RegFile.scala 66:20:@39743.4]
  wire  regs_151_reset; // @[RegFile.scala 66:20:@39743.4]
  wire [63:0] regs_151_io_in; // @[RegFile.scala 66:20:@39743.4]
  wire  regs_151_io_reset; // @[RegFile.scala 66:20:@39743.4]
  wire [63:0] regs_151_io_out; // @[RegFile.scala 66:20:@39743.4]
  wire  regs_151_io_enable; // @[RegFile.scala 66:20:@39743.4]
  wire  regs_152_clock; // @[RegFile.scala 66:20:@39757.4]
  wire  regs_152_reset; // @[RegFile.scala 66:20:@39757.4]
  wire [63:0] regs_152_io_in; // @[RegFile.scala 66:20:@39757.4]
  wire  regs_152_io_reset; // @[RegFile.scala 66:20:@39757.4]
  wire [63:0] regs_152_io_out; // @[RegFile.scala 66:20:@39757.4]
  wire  regs_152_io_enable; // @[RegFile.scala 66:20:@39757.4]
  wire  regs_153_clock; // @[RegFile.scala 66:20:@39771.4]
  wire  regs_153_reset; // @[RegFile.scala 66:20:@39771.4]
  wire [63:0] regs_153_io_in; // @[RegFile.scala 66:20:@39771.4]
  wire  regs_153_io_reset; // @[RegFile.scala 66:20:@39771.4]
  wire [63:0] regs_153_io_out; // @[RegFile.scala 66:20:@39771.4]
  wire  regs_153_io_enable; // @[RegFile.scala 66:20:@39771.4]
  wire  regs_154_clock; // @[RegFile.scala 66:20:@39785.4]
  wire  regs_154_reset; // @[RegFile.scala 66:20:@39785.4]
  wire [63:0] regs_154_io_in; // @[RegFile.scala 66:20:@39785.4]
  wire  regs_154_io_reset; // @[RegFile.scala 66:20:@39785.4]
  wire [63:0] regs_154_io_out; // @[RegFile.scala 66:20:@39785.4]
  wire  regs_154_io_enable; // @[RegFile.scala 66:20:@39785.4]
  wire  regs_155_clock; // @[RegFile.scala 66:20:@39799.4]
  wire  regs_155_reset; // @[RegFile.scala 66:20:@39799.4]
  wire [63:0] regs_155_io_in; // @[RegFile.scala 66:20:@39799.4]
  wire  regs_155_io_reset; // @[RegFile.scala 66:20:@39799.4]
  wire [63:0] regs_155_io_out; // @[RegFile.scala 66:20:@39799.4]
  wire  regs_155_io_enable; // @[RegFile.scala 66:20:@39799.4]
  wire  regs_156_clock; // @[RegFile.scala 66:20:@39813.4]
  wire  regs_156_reset; // @[RegFile.scala 66:20:@39813.4]
  wire [63:0] regs_156_io_in; // @[RegFile.scala 66:20:@39813.4]
  wire  regs_156_io_reset; // @[RegFile.scala 66:20:@39813.4]
  wire [63:0] regs_156_io_out; // @[RegFile.scala 66:20:@39813.4]
  wire  regs_156_io_enable; // @[RegFile.scala 66:20:@39813.4]
  wire  regs_157_clock; // @[RegFile.scala 66:20:@39827.4]
  wire  regs_157_reset; // @[RegFile.scala 66:20:@39827.4]
  wire [63:0] regs_157_io_in; // @[RegFile.scala 66:20:@39827.4]
  wire  regs_157_io_reset; // @[RegFile.scala 66:20:@39827.4]
  wire [63:0] regs_157_io_out; // @[RegFile.scala 66:20:@39827.4]
  wire  regs_157_io_enable; // @[RegFile.scala 66:20:@39827.4]
  wire  regs_158_clock; // @[RegFile.scala 66:20:@39841.4]
  wire  regs_158_reset; // @[RegFile.scala 66:20:@39841.4]
  wire [63:0] regs_158_io_in; // @[RegFile.scala 66:20:@39841.4]
  wire  regs_158_io_reset; // @[RegFile.scala 66:20:@39841.4]
  wire [63:0] regs_158_io_out; // @[RegFile.scala 66:20:@39841.4]
  wire  regs_158_io_enable; // @[RegFile.scala 66:20:@39841.4]
  wire  regs_159_clock; // @[RegFile.scala 66:20:@39855.4]
  wire  regs_159_reset; // @[RegFile.scala 66:20:@39855.4]
  wire [63:0] regs_159_io_in; // @[RegFile.scala 66:20:@39855.4]
  wire  regs_159_io_reset; // @[RegFile.scala 66:20:@39855.4]
  wire [63:0] regs_159_io_out; // @[RegFile.scala 66:20:@39855.4]
  wire  regs_159_io_enable; // @[RegFile.scala 66:20:@39855.4]
  wire  regs_160_clock; // @[RegFile.scala 66:20:@39869.4]
  wire  regs_160_reset; // @[RegFile.scala 66:20:@39869.4]
  wire [63:0] regs_160_io_in; // @[RegFile.scala 66:20:@39869.4]
  wire  regs_160_io_reset; // @[RegFile.scala 66:20:@39869.4]
  wire [63:0] regs_160_io_out; // @[RegFile.scala 66:20:@39869.4]
  wire  regs_160_io_enable; // @[RegFile.scala 66:20:@39869.4]
  wire  regs_161_clock; // @[RegFile.scala 66:20:@39883.4]
  wire  regs_161_reset; // @[RegFile.scala 66:20:@39883.4]
  wire [63:0] regs_161_io_in; // @[RegFile.scala 66:20:@39883.4]
  wire  regs_161_io_reset; // @[RegFile.scala 66:20:@39883.4]
  wire [63:0] regs_161_io_out; // @[RegFile.scala 66:20:@39883.4]
  wire  regs_161_io_enable; // @[RegFile.scala 66:20:@39883.4]
  wire  regs_162_clock; // @[RegFile.scala 66:20:@39897.4]
  wire  regs_162_reset; // @[RegFile.scala 66:20:@39897.4]
  wire [63:0] regs_162_io_in; // @[RegFile.scala 66:20:@39897.4]
  wire  regs_162_io_reset; // @[RegFile.scala 66:20:@39897.4]
  wire [63:0] regs_162_io_out; // @[RegFile.scala 66:20:@39897.4]
  wire  regs_162_io_enable; // @[RegFile.scala 66:20:@39897.4]
  wire  regs_163_clock; // @[RegFile.scala 66:20:@39911.4]
  wire  regs_163_reset; // @[RegFile.scala 66:20:@39911.4]
  wire [63:0] regs_163_io_in; // @[RegFile.scala 66:20:@39911.4]
  wire  regs_163_io_reset; // @[RegFile.scala 66:20:@39911.4]
  wire [63:0] regs_163_io_out; // @[RegFile.scala 66:20:@39911.4]
  wire  regs_163_io_enable; // @[RegFile.scala 66:20:@39911.4]
  wire  regs_164_clock; // @[RegFile.scala 66:20:@39925.4]
  wire  regs_164_reset; // @[RegFile.scala 66:20:@39925.4]
  wire [63:0] regs_164_io_in; // @[RegFile.scala 66:20:@39925.4]
  wire  regs_164_io_reset; // @[RegFile.scala 66:20:@39925.4]
  wire [63:0] regs_164_io_out; // @[RegFile.scala 66:20:@39925.4]
  wire  regs_164_io_enable; // @[RegFile.scala 66:20:@39925.4]
  wire  regs_165_clock; // @[RegFile.scala 66:20:@39939.4]
  wire  regs_165_reset; // @[RegFile.scala 66:20:@39939.4]
  wire [63:0] regs_165_io_in; // @[RegFile.scala 66:20:@39939.4]
  wire  regs_165_io_reset; // @[RegFile.scala 66:20:@39939.4]
  wire [63:0] regs_165_io_out; // @[RegFile.scala 66:20:@39939.4]
  wire  regs_165_io_enable; // @[RegFile.scala 66:20:@39939.4]
  wire  regs_166_clock; // @[RegFile.scala 66:20:@39953.4]
  wire  regs_166_reset; // @[RegFile.scala 66:20:@39953.4]
  wire [63:0] regs_166_io_in; // @[RegFile.scala 66:20:@39953.4]
  wire  regs_166_io_reset; // @[RegFile.scala 66:20:@39953.4]
  wire [63:0] regs_166_io_out; // @[RegFile.scala 66:20:@39953.4]
  wire  regs_166_io_enable; // @[RegFile.scala 66:20:@39953.4]
  wire  regs_167_clock; // @[RegFile.scala 66:20:@39967.4]
  wire  regs_167_reset; // @[RegFile.scala 66:20:@39967.4]
  wire [63:0] regs_167_io_in; // @[RegFile.scala 66:20:@39967.4]
  wire  regs_167_io_reset; // @[RegFile.scala 66:20:@39967.4]
  wire [63:0] regs_167_io_out; // @[RegFile.scala 66:20:@39967.4]
  wire  regs_167_io_enable; // @[RegFile.scala 66:20:@39967.4]
  wire  regs_168_clock; // @[RegFile.scala 66:20:@39981.4]
  wire  regs_168_reset; // @[RegFile.scala 66:20:@39981.4]
  wire [63:0] regs_168_io_in; // @[RegFile.scala 66:20:@39981.4]
  wire  regs_168_io_reset; // @[RegFile.scala 66:20:@39981.4]
  wire [63:0] regs_168_io_out; // @[RegFile.scala 66:20:@39981.4]
  wire  regs_168_io_enable; // @[RegFile.scala 66:20:@39981.4]
  wire  regs_169_clock; // @[RegFile.scala 66:20:@39995.4]
  wire  regs_169_reset; // @[RegFile.scala 66:20:@39995.4]
  wire [63:0] regs_169_io_in; // @[RegFile.scala 66:20:@39995.4]
  wire  regs_169_io_reset; // @[RegFile.scala 66:20:@39995.4]
  wire [63:0] regs_169_io_out; // @[RegFile.scala 66:20:@39995.4]
  wire  regs_169_io_enable; // @[RegFile.scala 66:20:@39995.4]
  wire  regs_170_clock; // @[RegFile.scala 66:20:@40009.4]
  wire  regs_170_reset; // @[RegFile.scala 66:20:@40009.4]
  wire [63:0] regs_170_io_in; // @[RegFile.scala 66:20:@40009.4]
  wire  regs_170_io_reset; // @[RegFile.scala 66:20:@40009.4]
  wire [63:0] regs_170_io_out; // @[RegFile.scala 66:20:@40009.4]
  wire  regs_170_io_enable; // @[RegFile.scala 66:20:@40009.4]
  wire  regs_171_clock; // @[RegFile.scala 66:20:@40023.4]
  wire  regs_171_reset; // @[RegFile.scala 66:20:@40023.4]
  wire [63:0] regs_171_io_in; // @[RegFile.scala 66:20:@40023.4]
  wire  regs_171_io_reset; // @[RegFile.scala 66:20:@40023.4]
  wire [63:0] regs_171_io_out; // @[RegFile.scala 66:20:@40023.4]
  wire  regs_171_io_enable; // @[RegFile.scala 66:20:@40023.4]
  wire  regs_172_clock; // @[RegFile.scala 66:20:@40037.4]
  wire  regs_172_reset; // @[RegFile.scala 66:20:@40037.4]
  wire [63:0] regs_172_io_in; // @[RegFile.scala 66:20:@40037.4]
  wire  regs_172_io_reset; // @[RegFile.scala 66:20:@40037.4]
  wire [63:0] regs_172_io_out; // @[RegFile.scala 66:20:@40037.4]
  wire  regs_172_io_enable; // @[RegFile.scala 66:20:@40037.4]
  wire  regs_173_clock; // @[RegFile.scala 66:20:@40051.4]
  wire  regs_173_reset; // @[RegFile.scala 66:20:@40051.4]
  wire [63:0] regs_173_io_in; // @[RegFile.scala 66:20:@40051.4]
  wire  regs_173_io_reset; // @[RegFile.scala 66:20:@40051.4]
  wire [63:0] regs_173_io_out; // @[RegFile.scala 66:20:@40051.4]
  wire  regs_173_io_enable; // @[RegFile.scala 66:20:@40051.4]
  wire  regs_174_clock; // @[RegFile.scala 66:20:@40065.4]
  wire  regs_174_reset; // @[RegFile.scala 66:20:@40065.4]
  wire [63:0] regs_174_io_in; // @[RegFile.scala 66:20:@40065.4]
  wire  regs_174_io_reset; // @[RegFile.scala 66:20:@40065.4]
  wire [63:0] regs_174_io_out; // @[RegFile.scala 66:20:@40065.4]
  wire  regs_174_io_enable; // @[RegFile.scala 66:20:@40065.4]
  wire  regs_175_clock; // @[RegFile.scala 66:20:@40079.4]
  wire  regs_175_reset; // @[RegFile.scala 66:20:@40079.4]
  wire [63:0] regs_175_io_in; // @[RegFile.scala 66:20:@40079.4]
  wire  regs_175_io_reset; // @[RegFile.scala 66:20:@40079.4]
  wire [63:0] regs_175_io_out; // @[RegFile.scala 66:20:@40079.4]
  wire  regs_175_io_enable; // @[RegFile.scala 66:20:@40079.4]
  wire  regs_176_clock; // @[RegFile.scala 66:20:@40093.4]
  wire  regs_176_reset; // @[RegFile.scala 66:20:@40093.4]
  wire [63:0] regs_176_io_in; // @[RegFile.scala 66:20:@40093.4]
  wire  regs_176_io_reset; // @[RegFile.scala 66:20:@40093.4]
  wire [63:0] regs_176_io_out; // @[RegFile.scala 66:20:@40093.4]
  wire  regs_176_io_enable; // @[RegFile.scala 66:20:@40093.4]
  wire  regs_177_clock; // @[RegFile.scala 66:20:@40107.4]
  wire  regs_177_reset; // @[RegFile.scala 66:20:@40107.4]
  wire [63:0] regs_177_io_in; // @[RegFile.scala 66:20:@40107.4]
  wire  regs_177_io_reset; // @[RegFile.scala 66:20:@40107.4]
  wire [63:0] regs_177_io_out; // @[RegFile.scala 66:20:@40107.4]
  wire  regs_177_io_enable; // @[RegFile.scala 66:20:@40107.4]
  wire  regs_178_clock; // @[RegFile.scala 66:20:@40121.4]
  wire  regs_178_reset; // @[RegFile.scala 66:20:@40121.4]
  wire [63:0] regs_178_io_in; // @[RegFile.scala 66:20:@40121.4]
  wire  regs_178_io_reset; // @[RegFile.scala 66:20:@40121.4]
  wire [63:0] regs_178_io_out; // @[RegFile.scala 66:20:@40121.4]
  wire  regs_178_io_enable; // @[RegFile.scala 66:20:@40121.4]
  wire  regs_179_clock; // @[RegFile.scala 66:20:@40135.4]
  wire  regs_179_reset; // @[RegFile.scala 66:20:@40135.4]
  wire [63:0] regs_179_io_in; // @[RegFile.scala 66:20:@40135.4]
  wire  regs_179_io_reset; // @[RegFile.scala 66:20:@40135.4]
  wire [63:0] regs_179_io_out; // @[RegFile.scala 66:20:@40135.4]
  wire  regs_179_io_enable; // @[RegFile.scala 66:20:@40135.4]
  wire  regs_180_clock; // @[RegFile.scala 66:20:@40149.4]
  wire  regs_180_reset; // @[RegFile.scala 66:20:@40149.4]
  wire [63:0] regs_180_io_in; // @[RegFile.scala 66:20:@40149.4]
  wire  regs_180_io_reset; // @[RegFile.scala 66:20:@40149.4]
  wire [63:0] regs_180_io_out; // @[RegFile.scala 66:20:@40149.4]
  wire  regs_180_io_enable; // @[RegFile.scala 66:20:@40149.4]
  wire  regs_181_clock; // @[RegFile.scala 66:20:@40163.4]
  wire  regs_181_reset; // @[RegFile.scala 66:20:@40163.4]
  wire [63:0] regs_181_io_in; // @[RegFile.scala 66:20:@40163.4]
  wire  regs_181_io_reset; // @[RegFile.scala 66:20:@40163.4]
  wire [63:0] regs_181_io_out; // @[RegFile.scala 66:20:@40163.4]
  wire  regs_181_io_enable; // @[RegFile.scala 66:20:@40163.4]
  wire  regs_182_clock; // @[RegFile.scala 66:20:@40177.4]
  wire  regs_182_reset; // @[RegFile.scala 66:20:@40177.4]
  wire [63:0] regs_182_io_in; // @[RegFile.scala 66:20:@40177.4]
  wire  regs_182_io_reset; // @[RegFile.scala 66:20:@40177.4]
  wire [63:0] regs_182_io_out; // @[RegFile.scala 66:20:@40177.4]
  wire  regs_182_io_enable; // @[RegFile.scala 66:20:@40177.4]
  wire  regs_183_clock; // @[RegFile.scala 66:20:@40191.4]
  wire  regs_183_reset; // @[RegFile.scala 66:20:@40191.4]
  wire [63:0] regs_183_io_in; // @[RegFile.scala 66:20:@40191.4]
  wire  regs_183_io_reset; // @[RegFile.scala 66:20:@40191.4]
  wire [63:0] regs_183_io_out; // @[RegFile.scala 66:20:@40191.4]
  wire  regs_183_io_enable; // @[RegFile.scala 66:20:@40191.4]
  wire  regs_184_clock; // @[RegFile.scala 66:20:@40205.4]
  wire  regs_184_reset; // @[RegFile.scala 66:20:@40205.4]
  wire [63:0] regs_184_io_in; // @[RegFile.scala 66:20:@40205.4]
  wire  regs_184_io_reset; // @[RegFile.scala 66:20:@40205.4]
  wire [63:0] regs_184_io_out; // @[RegFile.scala 66:20:@40205.4]
  wire  regs_184_io_enable; // @[RegFile.scala 66:20:@40205.4]
  wire  regs_185_clock; // @[RegFile.scala 66:20:@40219.4]
  wire  regs_185_reset; // @[RegFile.scala 66:20:@40219.4]
  wire [63:0] regs_185_io_in; // @[RegFile.scala 66:20:@40219.4]
  wire  regs_185_io_reset; // @[RegFile.scala 66:20:@40219.4]
  wire [63:0] regs_185_io_out; // @[RegFile.scala 66:20:@40219.4]
  wire  regs_185_io_enable; // @[RegFile.scala 66:20:@40219.4]
  wire  regs_186_clock; // @[RegFile.scala 66:20:@40233.4]
  wire  regs_186_reset; // @[RegFile.scala 66:20:@40233.4]
  wire [63:0] regs_186_io_in; // @[RegFile.scala 66:20:@40233.4]
  wire  regs_186_io_reset; // @[RegFile.scala 66:20:@40233.4]
  wire [63:0] regs_186_io_out; // @[RegFile.scala 66:20:@40233.4]
  wire  regs_186_io_enable; // @[RegFile.scala 66:20:@40233.4]
  wire  regs_187_clock; // @[RegFile.scala 66:20:@40247.4]
  wire  regs_187_reset; // @[RegFile.scala 66:20:@40247.4]
  wire [63:0] regs_187_io_in; // @[RegFile.scala 66:20:@40247.4]
  wire  regs_187_io_reset; // @[RegFile.scala 66:20:@40247.4]
  wire [63:0] regs_187_io_out; // @[RegFile.scala 66:20:@40247.4]
  wire  regs_187_io_enable; // @[RegFile.scala 66:20:@40247.4]
  wire  regs_188_clock; // @[RegFile.scala 66:20:@40261.4]
  wire  regs_188_reset; // @[RegFile.scala 66:20:@40261.4]
  wire [63:0] regs_188_io_in; // @[RegFile.scala 66:20:@40261.4]
  wire  regs_188_io_reset; // @[RegFile.scala 66:20:@40261.4]
  wire [63:0] regs_188_io_out; // @[RegFile.scala 66:20:@40261.4]
  wire  regs_188_io_enable; // @[RegFile.scala 66:20:@40261.4]
  wire  regs_189_clock; // @[RegFile.scala 66:20:@40275.4]
  wire  regs_189_reset; // @[RegFile.scala 66:20:@40275.4]
  wire [63:0] regs_189_io_in; // @[RegFile.scala 66:20:@40275.4]
  wire  regs_189_io_reset; // @[RegFile.scala 66:20:@40275.4]
  wire [63:0] regs_189_io_out; // @[RegFile.scala 66:20:@40275.4]
  wire  regs_189_io_enable; // @[RegFile.scala 66:20:@40275.4]
  wire  regs_190_clock; // @[RegFile.scala 66:20:@40289.4]
  wire  regs_190_reset; // @[RegFile.scala 66:20:@40289.4]
  wire [63:0] regs_190_io_in; // @[RegFile.scala 66:20:@40289.4]
  wire  regs_190_io_reset; // @[RegFile.scala 66:20:@40289.4]
  wire [63:0] regs_190_io_out; // @[RegFile.scala 66:20:@40289.4]
  wire  regs_190_io_enable; // @[RegFile.scala 66:20:@40289.4]
  wire  regs_191_clock; // @[RegFile.scala 66:20:@40303.4]
  wire  regs_191_reset; // @[RegFile.scala 66:20:@40303.4]
  wire [63:0] regs_191_io_in; // @[RegFile.scala 66:20:@40303.4]
  wire  regs_191_io_reset; // @[RegFile.scala 66:20:@40303.4]
  wire [63:0] regs_191_io_out; // @[RegFile.scala 66:20:@40303.4]
  wire  regs_191_io_enable; // @[RegFile.scala 66:20:@40303.4]
  wire  regs_192_clock; // @[RegFile.scala 66:20:@40317.4]
  wire  regs_192_reset; // @[RegFile.scala 66:20:@40317.4]
  wire [63:0] regs_192_io_in; // @[RegFile.scala 66:20:@40317.4]
  wire  regs_192_io_reset; // @[RegFile.scala 66:20:@40317.4]
  wire [63:0] regs_192_io_out; // @[RegFile.scala 66:20:@40317.4]
  wire  regs_192_io_enable; // @[RegFile.scala 66:20:@40317.4]
  wire  regs_193_clock; // @[RegFile.scala 66:20:@40331.4]
  wire  regs_193_reset; // @[RegFile.scala 66:20:@40331.4]
  wire [63:0] regs_193_io_in; // @[RegFile.scala 66:20:@40331.4]
  wire  regs_193_io_reset; // @[RegFile.scala 66:20:@40331.4]
  wire [63:0] regs_193_io_out; // @[RegFile.scala 66:20:@40331.4]
  wire  regs_193_io_enable; // @[RegFile.scala 66:20:@40331.4]
  wire  regs_194_clock; // @[RegFile.scala 66:20:@40345.4]
  wire  regs_194_reset; // @[RegFile.scala 66:20:@40345.4]
  wire [63:0] regs_194_io_in; // @[RegFile.scala 66:20:@40345.4]
  wire  regs_194_io_reset; // @[RegFile.scala 66:20:@40345.4]
  wire [63:0] regs_194_io_out; // @[RegFile.scala 66:20:@40345.4]
  wire  regs_194_io_enable; // @[RegFile.scala 66:20:@40345.4]
  wire  regs_195_clock; // @[RegFile.scala 66:20:@40359.4]
  wire  regs_195_reset; // @[RegFile.scala 66:20:@40359.4]
  wire [63:0] regs_195_io_in; // @[RegFile.scala 66:20:@40359.4]
  wire  regs_195_io_reset; // @[RegFile.scala 66:20:@40359.4]
  wire [63:0] regs_195_io_out; // @[RegFile.scala 66:20:@40359.4]
  wire  regs_195_io_enable; // @[RegFile.scala 66:20:@40359.4]
  wire  regs_196_clock; // @[RegFile.scala 66:20:@40373.4]
  wire  regs_196_reset; // @[RegFile.scala 66:20:@40373.4]
  wire [63:0] regs_196_io_in; // @[RegFile.scala 66:20:@40373.4]
  wire  regs_196_io_reset; // @[RegFile.scala 66:20:@40373.4]
  wire [63:0] regs_196_io_out; // @[RegFile.scala 66:20:@40373.4]
  wire  regs_196_io_enable; // @[RegFile.scala 66:20:@40373.4]
  wire  regs_197_clock; // @[RegFile.scala 66:20:@40387.4]
  wire  regs_197_reset; // @[RegFile.scala 66:20:@40387.4]
  wire [63:0] regs_197_io_in; // @[RegFile.scala 66:20:@40387.4]
  wire  regs_197_io_reset; // @[RegFile.scala 66:20:@40387.4]
  wire [63:0] regs_197_io_out; // @[RegFile.scala 66:20:@40387.4]
  wire  regs_197_io_enable; // @[RegFile.scala 66:20:@40387.4]
  wire  regs_198_clock; // @[RegFile.scala 66:20:@40401.4]
  wire  regs_198_reset; // @[RegFile.scala 66:20:@40401.4]
  wire [63:0] regs_198_io_in; // @[RegFile.scala 66:20:@40401.4]
  wire  regs_198_io_reset; // @[RegFile.scala 66:20:@40401.4]
  wire [63:0] regs_198_io_out; // @[RegFile.scala 66:20:@40401.4]
  wire  regs_198_io_enable; // @[RegFile.scala 66:20:@40401.4]
  wire  regs_199_clock; // @[RegFile.scala 66:20:@40415.4]
  wire  regs_199_reset; // @[RegFile.scala 66:20:@40415.4]
  wire [63:0] regs_199_io_in; // @[RegFile.scala 66:20:@40415.4]
  wire  regs_199_io_reset; // @[RegFile.scala 66:20:@40415.4]
  wire [63:0] regs_199_io_out; // @[RegFile.scala 66:20:@40415.4]
  wire  regs_199_io_enable; // @[RegFile.scala 66:20:@40415.4]
  wire  regs_200_clock; // @[RegFile.scala 66:20:@40429.4]
  wire  regs_200_reset; // @[RegFile.scala 66:20:@40429.4]
  wire [63:0] regs_200_io_in; // @[RegFile.scala 66:20:@40429.4]
  wire  regs_200_io_reset; // @[RegFile.scala 66:20:@40429.4]
  wire [63:0] regs_200_io_out; // @[RegFile.scala 66:20:@40429.4]
  wire  regs_200_io_enable; // @[RegFile.scala 66:20:@40429.4]
  wire  regs_201_clock; // @[RegFile.scala 66:20:@40443.4]
  wire  regs_201_reset; // @[RegFile.scala 66:20:@40443.4]
  wire [63:0] regs_201_io_in; // @[RegFile.scala 66:20:@40443.4]
  wire  regs_201_io_reset; // @[RegFile.scala 66:20:@40443.4]
  wire [63:0] regs_201_io_out; // @[RegFile.scala 66:20:@40443.4]
  wire  regs_201_io_enable; // @[RegFile.scala 66:20:@40443.4]
  wire  regs_202_clock; // @[RegFile.scala 66:20:@40457.4]
  wire  regs_202_reset; // @[RegFile.scala 66:20:@40457.4]
  wire [63:0] regs_202_io_in; // @[RegFile.scala 66:20:@40457.4]
  wire  regs_202_io_reset; // @[RegFile.scala 66:20:@40457.4]
  wire [63:0] regs_202_io_out; // @[RegFile.scala 66:20:@40457.4]
  wire  regs_202_io_enable; // @[RegFile.scala 66:20:@40457.4]
  wire  regs_203_clock; // @[RegFile.scala 66:20:@40471.4]
  wire  regs_203_reset; // @[RegFile.scala 66:20:@40471.4]
  wire [63:0] regs_203_io_in; // @[RegFile.scala 66:20:@40471.4]
  wire  regs_203_io_reset; // @[RegFile.scala 66:20:@40471.4]
  wire [63:0] regs_203_io_out; // @[RegFile.scala 66:20:@40471.4]
  wire  regs_203_io_enable; // @[RegFile.scala 66:20:@40471.4]
  wire  regs_204_clock; // @[RegFile.scala 66:20:@40485.4]
  wire  regs_204_reset; // @[RegFile.scala 66:20:@40485.4]
  wire [63:0] regs_204_io_in; // @[RegFile.scala 66:20:@40485.4]
  wire  regs_204_io_reset; // @[RegFile.scala 66:20:@40485.4]
  wire [63:0] regs_204_io_out; // @[RegFile.scala 66:20:@40485.4]
  wire  regs_204_io_enable; // @[RegFile.scala 66:20:@40485.4]
  wire  regs_205_clock; // @[RegFile.scala 66:20:@40499.4]
  wire  regs_205_reset; // @[RegFile.scala 66:20:@40499.4]
  wire [63:0] regs_205_io_in; // @[RegFile.scala 66:20:@40499.4]
  wire  regs_205_io_reset; // @[RegFile.scala 66:20:@40499.4]
  wire [63:0] regs_205_io_out; // @[RegFile.scala 66:20:@40499.4]
  wire  regs_205_io_enable; // @[RegFile.scala 66:20:@40499.4]
  wire  regs_206_clock; // @[RegFile.scala 66:20:@40513.4]
  wire  regs_206_reset; // @[RegFile.scala 66:20:@40513.4]
  wire [63:0] regs_206_io_in; // @[RegFile.scala 66:20:@40513.4]
  wire  regs_206_io_reset; // @[RegFile.scala 66:20:@40513.4]
  wire [63:0] regs_206_io_out; // @[RegFile.scala 66:20:@40513.4]
  wire  regs_206_io_enable; // @[RegFile.scala 66:20:@40513.4]
  wire  regs_207_clock; // @[RegFile.scala 66:20:@40527.4]
  wire  regs_207_reset; // @[RegFile.scala 66:20:@40527.4]
  wire [63:0] regs_207_io_in; // @[RegFile.scala 66:20:@40527.4]
  wire  regs_207_io_reset; // @[RegFile.scala 66:20:@40527.4]
  wire [63:0] regs_207_io_out; // @[RegFile.scala 66:20:@40527.4]
  wire  regs_207_io_enable; // @[RegFile.scala 66:20:@40527.4]
  wire  regs_208_clock; // @[RegFile.scala 66:20:@40541.4]
  wire  regs_208_reset; // @[RegFile.scala 66:20:@40541.4]
  wire [63:0] regs_208_io_in; // @[RegFile.scala 66:20:@40541.4]
  wire  regs_208_io_reset; // @[RegFile.scala 66:20:@40541.4]
  wire [63:0] regs_208_io_out; // @[RegFile.scala 66:20:@40541.4]
  wire  regs_208_io_enable; // @[RegFile.scala 66:20:@40541.4]
  wire  regs_209_clock; // @[RegFile.scala 66:20:@40555.4]
  wire  regs_209_reset; // @[RegFile.scala 66:20:@40555.4]
  wire [63:0] regs_209_io_in; // @[RegFile.scala 66:20:@40555.4]
  wire  regs_209_io_reset; // @[RegFile.scala 66:20:@40555.4]
  wire [63:0] regs_209_io_out; // @[RegFile.scala 66:20:@40555.4]
  wire  regs_209_io_enable; // @[RegFile.scala 66:20:@40555.4]
  wire  regs_210_clock; // @[RegFile.scala 66:20:@40569.4]
  wire  regs_210_reset; // @[RegFile.scala 66:20:@40569.4]
  wire [63:0] regs_210_io_in; // @[RegFile.scala 66:20:@40569.4]
  wire  regs_210_io_reset; // @[RegFile.scala 66:20:@40569.4]
  wire [63:0] regs_210_io_out; // @[RegFile.scala 66:20:@40569.4]
  wire  regs_210_io_enable; // @[RegFile.scala 66:20:@40569.4]
  wire  regs_211_clock; // @[RegFile.scala 66:20:@40583.4]
  wire  regs_211_reset; // @[RegFile.scala 66:20:@40583.4]
  wire [63:0] regs_211_io_in; // @[RegFile.scala 66:20:@40583.4]
  wire  regs_211_io_reset; // @[RegFile.scala 66:20:@40583.4]
  wire [63:0] regs_211_io_out; // @[RegFile.scala 66:20:@40583.4]
  wire  regs_211_io_enable; // @[RegFile.scala 66:20:@40583.4]
  wire  regs_212_clock; // @[RegFile.scala 66:20:@40597.4]
  wire  regs_212_reset; // @[RegFile.scala 66:20:@40597.4]
  wire [63:0] regs_212_io_in; // @[RegFile.scala 66:20:@40597.4]
  wire  regs_212_io_reset; // @[RegFile.scala 66:20:@40597.4]
  wire [63:0] regs_212_io_out; // @[RegFile.scala 66:20:@40597.4]
  wire  regs_212_io_enable; // @[RegFile.scala 66:20:@40597.4]
  wire  regs_213_clock; // @[RegFile.scala 66:20:@40611.4]
  wire  regs_213_reset; // @[RegFile.scala 66:20:@40611.4]
  wire [63:0] regs_213_io_in; // @[RegFile.scala 66:20:@40611.4]
  wire  regs_213_io_reset; // @[RegFile.scala 66:20:@40611.4]
  wire [63:0] regs_213_io_out; // @[RegFile.scala 66:20:@40611.4]
  wire  regs_213_io_enable; // @[RegFile.scala 66:20:@40611.4]
  wire  regs_214_clock; // @[RegFile.scala 66:20:@40625.4]
  wire  regs_214_reset; // @[RegFile.scala 66:20:@40625.4]
  wire [63:0] regs_214_io_in; // @[RegFile.scala 66:20:@40625.4]
  wire  regs_214_io_reset; // @[RegFile.scala 66:20:@40625.4]
  wire [63:0] regs_214_io_out; // @[RegFile.scala 66:20:@40625.4]
  wire  regs_214_io_enable; // @[RegFile.scala 66:20:@40625.4]
  wire  regs_215_clock; // @[RegFile.scala 66:20:@40639.4]
  wire  regs_215_reset; // @[RegFile.scala 66:20:@40639.4]
  wire [63:0] regs_215_io_in; // @[RegFile.scala 66:20:@40639.4]
  wire  regs_215_io_reset; // @[RegFile.scala 66:20:@40639.4]
  wire [63:0] regs_215_io_out; // @[RegFile.scala 66:20:@40639.4]
  wire  regs_215_io_enable; // @[RegFile.scala 66:20:@40639.4]
  wire  regs_216_clock; // @[RegFile.scala 66:20:@40653.4]
  wire  regs_216_reset; // @[RegFile.scala 66:20:@40653.4]
  wire [63:0] regs_216_io_in; // @[RegFile.scala 66:20:@40653.4]
  wire  regs_216_io_reset; // @[RegFile.scala 66:20:@40653.4]
  wire [63:0] regs_216_io_out; // @[RegFile.scala 66:20:@40653.4]
  wire  regs_216_io_enable; // @[RegFile.scala 66:20:@40653.4]
  wire  regs_217_clock; // @[RegFile.scala 66:20:@40667.4]
  wire  regs_217_reset; // @[RegFile.scala 66:20:@40667.4]
  wire [63:0] regs_217_io_in; // @[RegFile.scala 66:20:@40667.4]
  wire  regs_217_io_reset; // @[RegFile.scala 66:20:@40667.4]
  wire [63:0] regs_217_io_out; // @[RegFile.scala 66:20:@40667.4]
  wire  regs_217_io_enable; // @[RegFile.scala 66:20:@40667.4]
  wire  regs_218_clock; // @[RegFile.scala 66:20:@40681.4]
  wire  regs_218_reset; // @[RegFile.scala 66:20:@40681.4]
  wire [63:0] regs_218_io_in; // @[RegFile.scala 66:20:@40681.4]
  wire  regs_218_io_reset; // @[RegFile.scala 66:20:@40681.4]
  wire [63:0] regs_218_io_out; // @[RegFile.scala 66:20:@40681.4]
  wire  regs_218_io_enable; // @[RegFile.scala 66:20:@40681.4]
  wire  regs_219_clock; // @[RegFile.scala 66:20:@40695.4]
  wire  regs_219_reset; // @[RegFile.scala 66:20:@40695.4]
  wire [63:0] regs_219_io_in; // @[RegFile.scala 66:20:@40695.4]
  wire  regs_219_io_reset; // @[RegFile.scala 66:20:@40695.4]
  wire [63:0] regs_219_io_out; // @[RegFile.scala 66:20:@40695.4]
  wire  regs_219_io_enable; // @[RegFile.scala 66:20:@40695.4]
  wire  regs_220_clock; // @[RegFile.scala 66:20:@40709.4]
  wire  regs_220_reset; // @[RegFile.scala 66:20:@40709.4]
  wire [63:0] regs_220_io_in; // @[RegFile.scala 66:20:@40709.4]
  wire  regs_220_io_reset; // @[RegFile.scala 66:20:@40709.4]
  wire [63:0] regs_220_io_out; // @[RegFile.scala 66:20:@40709.4]
  wire  regs_220_io_enable; // @[RegFile.scala 66:20:@40709.4]
  wire  regs_221_clock; // @[RegFile.scala 66:20:@40723.4]
  wire  regs_221_reset; // @[RegFile.scala 66:20:@40723.4]
  wire [63:0] regs_221_io_in; // @[RegFile.scala 66:20:@40723.4]
  wire  regs_221_io_reset; // @[RegFile.scala 66:20:@40723.4]
  wire [63:0] regs_221_io_out; // @[RegFile.scala 66:20:@40723.4]
  wire  regs_221_io_enable; // @[RegFile.scala 66:20:@40723.4]
  wire  regs_222_clock; // @[RegFile.scala 66:20:@40737.4]
  wire  regs_222_reset; // @[RegFile.scala 66:20:@40737.4]
  wire [63:0] regs_222_io_in; // @[RegFile.scala 66:20:@40737.4]
  wire  regs_222_io_reset; // @[RegFile.scala 66:20:@40737.4]
  wire [63:0] regs_222_io_out; // @[RegFile.scala 66:20:@40737.4]
  wire  regs_222_io_enable; // @[RegFile.scala 66:20:@40737.4]
  wire  regs_223_clock; // @[RegFile.scala 66:20:@40751.4]
  wire  regs_223_reset; // @[RegFile.scala 66:20:@40751.4]
  wire [63:0] regs_223_io_in; // @[RegFile.scala 66:20:@40751.4]
  wire  regs_223_io_reset; // @[RegFile.scala 66:20:@40751.4]
  wire [63:0] regs_223_io_out; // @[RegFile.scala 66:20:@40751.4]
  wire  regs_223_io_enable; // @[RegFile.scala 66:20:@40751.4]
  wire  regs_224_clock; // @[RegFile.scala 66:20:@40765.4]
  wire  regs_224_reset; // @[RegFile.scala 66:20:@40765.4]
  wire [63:0] regs_224_io_in; // @[RegFile.scala 66:20:@40765.4]
  wire  regs_224_io_reset; // @[RegFile.scala 66:20:@40765.4]
  wire [63:0] regs_224_io_out; // @[RegFile.scala 66:20:@40765.4]
  wire  regs_224_io_enable; // @[RegFile.scala 66:20:@40765.4]
  wire  regs_225_clock; // @[RegFile.scala 66:20:@40779.4]
  wire  regs_225_reset; // @[RegFile.scala 66:20:@40779.4]
  wire [63:0] regs_225_io_in; // @[RegFile.scala 66:20:@40779.4]
  wire  regs_225_io_reset; // @[RegFile.scala 66:20:@40779.4]
  wire [63:0] regs_225_io_out; // @[RegFile.scala 66:20:@40779.4]
  wire  regs_225_io_enable; // @[RegFile.scala 66:20:@40779.4]
  wire  regs_226_clock; // @[RegFile.scala 66:20:@40793.4]
  wire  regs_226_reset; // @[RegFile.scala 66:20:@40793.4]
  wire [63:0] regs_226_io_in; // @[RegFile.scala 66:20:@40793.4]
  wire  regs_226_io_reset; // @[RegFile.scala 66:20:@40793.4]
  wire [63:0] regs_226_io_out; // @[RegFile.scala 66:20:@40793.4]
  wire  regs_226_io_enable; // @[RegFile.scala 66:20:@40793.4]
  wire  regs_227_clock; // @[RegFile.scala 66:20:@40807.4]
  wire  regs_227_reset; // @[RegFile.scala 66:20:@40807.4]
  wire [63:0] regs_227_io_in; // @[RegFile.scala 66:20:@40807.4]
  wire  regs_227_io_reset; // @[RegFile.scala 66:20:@40807.4]
  wire [63:0] regs_227_io_out; // @[RegFile.scala 66:20:@40807.4]
  wire  regs_227_io_enable; // @[RegFile.scala 66:20:@40807.4]
  wire  regs_228_clock; // @[RegFile.scala 66:20:@40821.4]
  wire  regs_228_reset; // @[RegFile.scala 66:20:@40821.4]
  wire [63:0] regs_228_io_in; // @[RegFile.scala 66:20:@40821.4]
  wire  regs_228_io_reset; // @[RegFile.scala 66:20:@40821.4]
  wire [63:0] regs_228_io_out; // @[RegFile.scala 66:20:@40821.4]
  wire  regs_228_io_enable; // @[RegFile.scala 66:20:@40821.4]
  wire  regs_229_clock; // @[RegFile.scala 66:20:@40835.4]
  wire  regs_229_reset; // @[RegFile.scala 66:20:@40835.4]
  wire [63:0] regs_229_io_in; // @[RegFile.scala 66:20:@40835.4]
  wire  regs_229_io_reset; // @[RegFile.scala 66:20:@40835.4]
  wire [63:0] regs_229_io_out; // @[RegFile.scala 66:20:@40835.4]
  wire  regs_229_io_enable; // @[RegFile.scala 66:20:@40835.4]
  wire  regs_230_clock; // @[RegFile.scala 66:20:@40849.4]
  wire  regs_230_reset; // @[RegFile.scala 66:20:@40849.4]
  wire [63:0] regs_230_io_in; // @[RegFile.scala 66:20:@40849.4]
  wire  regs_230_io_reset; // @[RegFile.scala 66:20:@40849.4]
  wire [63:0] regs_230_io_out; // @[RegFile.scala 66:20:@40849.4]
  wire  regs_230_io_enable; // @[RegFile.scala 66:20:@40849.4]
  wire  regs_231_clock; // @[RegFile.scala 66:20:@40863.4]
  wire  regs_231_reset; // @[RegFile.scala 66:20:@40863.4]
  wire [63:0] regs_231_io_in; // @[RegFile.scala 66:20:@40863.4]
  wire  regs_231_io_reset; // @[RegFile.scala 66:20:@40863.4]
  wire [63:0] regs_231_io_out; // @[RegFile.scala 66:20:@40863.4]
  wire  regs_231_io_enable; // @[RegFile.scala 66:20:@40863.4]
  wire  regs_232_clock; // @[RegFile.scala 66:20:@40877.4]
  wire  regs_232_reset; // @[RegFile.scala 66:20:@40877.4]
  wire [63:0] regs_232_io_in; // @[RegFile.scala 66:20:@40877.4]
  wire  regs_232_io_reset; // @[RegFile.scala 66:20:@40877.4]
  wire [63:0] regs_232_io_out; // @[RegFile.scala 66:20:@40877.4]
  wire  regs_232_io_enable; // @[RegFile.scala 66:20:@40877.4]
  wire  regs_233_clock; // @[RegFile.scala 66:20:@40891.4]
  wire  regs_233_reset; // @[RegFile.scala 66:20:@40891.4]
  wire [63:0] regs_233_io_in; // @[RegFile.scala 66:20:@40891.4]
  wire  regs_233_io_reset; // @[RegFile.scala 66:20:@40891.4]
  wire [63:0] regs_233_io_out; // @[RegFile.scala 66:20:@40891.4]
  wire  regs_233_io_enable; // @[RegFile.scala 66:20:@40891.4]
  wire  regs_234_clock; // @[RegFile.scala 66:20:@40905.4]
  wire  regs_234_reset; // @[RegFile.scala 66:20:@40905.4]
  wire [63:0] regs_234_io_in; // @[RegFile.scala 66:20:@40905.4]
  wire  regs_234_io_reset; // @[RegFile.scala 66:20:@40905.4]
  wire [63:0] regs_234_io_out; // @[RegFile.scala 66:20:@40905.4]
  wire  regs_234_io_enable; // @[RegFile.scala 66:20:@40905.4]
  wire  regs_235_clock; // @[RegFile.scala 66:20:@40919.4]
  wire  regs_235_reset; // @[RegFile.scala 66:20:@40919.4]
  wire [63:0] regs_235_io_in; // @[RegFile.scala 66:20:@40919.4]
  wire  regs_235_io_reset; // @[RegFile.scala 66:20:@40919.4]
  wire [63:0] regs_235_io_out; // @[RegFile.scala 66:20:@40919.4]
  wire  regs_235_io_enable; // @[RegFile.scala 66:20:@40919.4]
  wire  regs_236_clock; // @[RegFile.scala 66:20:@40933.4]
  wire  regs_236_reset; // @[RegFile.scala 66:20:@40933.4]
  wire [63:0] regs_236_io_in; // @[RegFile.scala 66:20:@40933.4]
  wire  regs_236_io_reset; // @[RegFile.scala 66:20:@40933.4]
  wire [63:0] regs_236_io_out; // @[RegFile.scala 66:20:@40933.4]
  wire  regs_236_io_enable; // @[RegFile.scala 66:20:@40933.4]
  wire  regs_237_clock; // @[RegFile.scala 66:20:@40947.4]
  wire  regs_237_reset; // @[RegFile.scala 66:20:@40947.4]
  wire [63:0] regs_237_io_in; // @[RegFile.scala 66:20:@40947.4]
  wire  regs_237_io_reset; // @[RegFile.scala 66:20:@40947.4]
  wire [63:0] regs_237_io_out; // @[RegFile.scala 66:20:@40947.4]
  wire  regs_237_io_enable; // @[RegFile.scala 66:20:@40947.4]
  wire  regs_238_clock; // @[RegFile.scala 66:20:@40961.4]
  wire  regs_238_reset; // @[RegFile.scala 66:20:@40961.4]
  wire [63:0] regs_238_io_in; // @[RegFile.scala 66:20:@40961.4]
  wire  regs_238_io_reset; // @[RegFile.scala 66:20:@40961.4]
  wire [63:0] regs_238_io_out; // @[RegFile.scala 66:20:@40961.4]
  wire  regs_238_io_enable; // @[RegFile.scala 66:20:@40961.4]
  wire  regs_239_clock; // @[RegFile.scala 66:20:@40975.4]
  wire  regs_239_reset; // @[RegFile.scala 66:20:@40975.4]
  wire [63:0] regs_239_io_in; // @[RegFile.scala 66:20:@40975.4]
  wire  regs_239_io_reset; // @[RegFile.scala 66:20:@40975.4]
  wire [63:0] regs_239_io_out; // @[RegFile.scala 66:20:@40975.4]
  wire  regs_239_io_enable; // @[RegFile.scala 66:20:@40975.4]
  wire  regs_240_clock; // @[RegFile.scala 66:20:@40989.4]
  wire  regs_240_reset; // @[RegFile.scala 66:20:@40989.4]
  wire [63:0] regs_240_io_in; // @[RegFile.scala 66:20:@40989.4]
  wire  regs_240_io_reset; // @[RegFile.scala 66:20:@40989.4]
  wire [63:0] regs_240_io_out; // @[RegFile.scala 66:20:@40989.4]
  wire  regs_240_io_enable; // @[RegFile.scala 66:20:@40989.4]
  wire  regs_241_clock; // @[RegFile.scala 66:20:@41003.4]
  wire  regs_241_reset; // @[RegFile.scala 66:20:@41003.4]
  wire [63:0] regs_241_io_in; // @[RegFile.scala 66:20:@41003.4]
  wire  regs_241_io_reset; // @[RegFile.scala 66:20:@41003.4]
  wire [63:0] regs_241_io_out; // @[RegFile.scala 66:20:@41003.4]
  wire  regs_241_io_enable; // @[RegFile.scala 66:20:@41003.4]
  wire  regs_242_clock; // @[RegFile.scala 66:20:@41017.4]
  wire  regs_242_reset; // @[RegFile.scala 66:20:@41017.4]
  wire [63:0] regs_242_io_in; // @[RegFile.scala 66:20:@41017.4]
  wire  regs_242_io_reset; // @[RegFile.scala 66:20:@41017.4]
  wire [63:0] regs_242_io_out; // @[RegFile.scala 66:20:@41017.4]
  wire  regs_242_io_enable; // @[RegFile.scala 66:20:@41017.4]
  wire  regs_243_clock; // @[RegFile.scala 66:20:@41031.4]
  wire  regs_243_reset; // @[RegFile.scala 66:20:@41031.4]
  wire [63:0] regs_243_io_in; // @[RegFile.scala 66:20:@41031.4]
  wire  regs_243_io_reset; // @[RegFile.scala 66:20:@41031.4]
  wire [63:0] regs_243_io_out; // @[RegFile.scala 66:20:@41031.4]
  wire  regs_243_io_enable; // @[RegFile.scala 66:20:@41031.4]
  wire  regs_244_clock; // @[RegFile.scala 66:20:@41045.4]
  wire  regs_244_reset; // @[RegFile.scala 66:20:@41045.4]
  wire [63:0] regs_244_io_in; // @[RegFile.scala 66:20:@41045.4]
  wire  regs_244_io_reset; // @[RegFile.scala 66:20:@41045.4]
  wire [63:0] regs_244_io_out; // @[RegFile.scala 66:20:@41045.4]
  wire  regs_244_io_enable; // @[RegFile.scala 66:20:@41045.4]
  wire  regs_245_clock; // @[RegFile.scala 66:20:@41059.4]
  wire  regs_245_reset; // @[RegFile.scala 66:20:@41059.4]
  wire [63:0] regs_245_io_in; // @[RegFile.scala 66:20:@41059.4]
  wire  regs_245_io_reset; // @[RegFile.scala 66:20:@41059.4]
  wire [63:0] regs_245_io_out; // @[RegFile.scala 66:20:@41059.4]
  wire  regs_245_io_enable; // @[RegFile.scala 66:20:@41059.4]
  wire  regs_246_clock; // @[RegFile.scala 66:20:@41073.4]
  wire  regs_246_reset; // @[RegFile.scala 66:20:@41073.4]
  wire [63:0] regs_246_io_in; // @[RegFile.scala 66:20:@41073.4]
  wire  regs_246_io_reset; // @[RegFile.scala 66:20:@41073.4]
  wire [63:0] regs_246_io_out; // @[RegFile.scala 66:20:@41073.4]
  wire  regs_246_io_enable; // @[RegFile.scala 66:20:@41073.4]
  wire  regs_247_clock; // @[RegFile.scala 66:20:@41087.4]
  wire  regs_247_reset; // @[RegFile.scala 66:20:@41087.4]
  wire [63:0] regs_247_io_in; // @[RegFile.scala 66:20:@41087.4]
  wire  regs_247_io_reset; // @[RegFile.scala 66:20:@41087.4]
  wire [63:0] regs_247_io_out; // @[RegFile.scala 66:20:@41087.4]
  wire  regs_247_io_enable; // @[RegFile.scala 66:20:@41087.4]
  wire  regs_248_clock; // @[RegFile.scala 66:20:@41101.4]
  wire  regs_248_reset; // @[RegFile.scala 66:20:@41101.4]
  wire [63:0] regs_248_io_in; // @[RegFile.scala 66:20:@41101.4]
  wire  regs_248_io_reset; // @[RegFile.scala 66:20:@41101.4]
  wire [63:0] regs_248_io_out; // @[RegFile.scala 66:20:@41101.4]
  wire  regs_248_io_enable; // @[RegFile.scala 66:20:@41101.4]
  wire  regs_249_clock; // @[RegFile.scala 66:20:@41115.4]
  wire  regs_249_reset; // @[RegFile.scala 66:20:@41115.4]
  wire [63:0] regs_249_io_in; // @[RegFile.scala 66:20:@41115.4]
  wire  regs_249_io_reset; // @[RegFile.scala 66:20:@41115.4]
  wire [63:0] regs_249_io_out; // @[RegFile.scala 66:20:@41115.4]
  wire  regs_249_io_enable; // @[RegFile.scala 66:20:@41115.4]
  wire  regs_250_clock; // @[RegFile.scala 66:20:@41129.4]
  wire  regs_250_reset; // @[RegFile.scala 66:20:@41129.4]
  wire [63:0] regs_250_io_in; // @[RegFile.scala 66:20:@41129.4]
  wire  regs_250_io_reset; // @[RegFile.scala 66:20:@41129.4]
  wire [63:0] regs_250_io_out; // @[RegFile.scala 66:20:@41129.4]
  wire  regs_250_io_enable; // @[RegFile.scala 66:20:@41129.4]
  wire  regs_251_clock; // @[RegFile.scala 66:20:@41143.4]
  wire  regs_251_reset; // @[RegFile.scala 66:20:@41143.4]
  wire [63:0] regs_251_io_in; // @[RegFile.scala 66:20:@41143.4]
  wire  regs_251_io_reset; // @[RegFile.scala 66:20:@41143.4]
  wire [63:0] regs_251_io_out; // @[RegFile.scala 66:20:@41143.4]
  wire  regs_251_io_enable; // @[RegFile.scala 66:20:@41143.4]
  wire  regs_252_clock; // @[RegFile.scala 66:20:@41157.4]
  wire  regs_252_reset; // @[RegFile.scala 66:20:@41157.4]
  wire [63:0] regs_252_io_in; // @[RegFile.scala 66:20:@41157.4]
  wire  regs_252_io_reset; // @[RegFile.scala 66:20:@41157.4]
  wire [63:0] regs_252_io_out; // @[RegFile.scala 66:20:@41157.4]
  wire  regs_252_io_enable; // @[RegFile.scala 66:20:@41157.4]
  wire  regs_253_clock; // @[RegFile.scala 66:20:@41171.4]
  wire  regs_253_reset; // @[RegFile.scala 66:20:@41171.4]
  wire [63:0] regs_253_io_in; // @[RegFile.scala 66:20:@41171.4]
  wire  regs_253_io_reset; // @[RegFile.scala 66:20:@41171.4]
  wire [63:0] regs_253_io_out; // @[RegFile.scala 66:20:@41171.4]
  wire  regs_253_io_enable; // @[RegFile.scala 66:20:@41171.4]
  wire  regs_254_clock; // @[RegFile.scala 66:20:@41185.4]
  wire  regs_254_reset; // @[RegFile.scala 66:20:@41185.4]
  wire [63:0] regs_254_io_in; // @[RegFile.scala 66:20:@41185.4]
  wire  regs_254_io_reset; // @[RegFile.scala 66:20:@41185.4]
  wire [63:0] regs_254_io_out; // @[RegFile.scala 66:20:@41185.4]
  wire  regs_254_io_enable; // @[RegFile.scala 66:20:@41185.4]
  wire  regs_255_clock; // @[RegFile.scala 66:20:@41199.4]
  wire  regs_255_reset; // @[RegFile.scala 66:20:@41199.4]
  wire [63:0] regs_255_io_in; // @[RegFile.scala 66:20:@41199.4]
  wire  regs_255_io_reset; // @[RegFile.scala 66:20:@41199.4]
  wire [63:0] regs_255_io_out; // @[RegFile.scala 66:20:@41199.4]
  wire  regs_255_io_enable; // @[RegFile.scala 66:20:@41199.4]
  wire  regs_256_clock; // @[RegFile.scala 66:20:@41213.4]
  wire  regs_256_reset; // @[RegFile.scala 66:20:@41213.4]
  wire [63:0] regs_256_io_in; // @[RegFile.scala 66:20:@41213.4]
  wire  regs_256_io_reset; // @[RegFile.scala 66:20:@41213.4]
  wire [63:0] regs_256_io_out; // @[RegFile.scala 66:20:@41213.4]
  wire  regs_256_io_enable; // @[RegFile.scala 66:20:@41213.4]
  wire  regs_257_clock; // @[RegFile.scala 66:20:@41227.4]
  wire  regs_257_reset; // @[RegFile.scala 66:20:@41227.4]
  wire [63:0] regs_257_io_in; // @[RegFile.scala 66:20:@41227.4]
  wire  regs_257_io_reset; // @[RegFile.scala 66:20:@41227.4]
  wire [63:0] regs_257_io_out; // @[RegFile.scala 66:20:@41227.4]
  wire  regs_257_io_enable; // @[RegFile.scala 66:20:@41227.4]
  wire  regs_258_clock; // @[RegFile.scala 66:20:@41241.4]
  wire  regs_258_reset; // @[RegFile.scala 66:20:@41241.4]
  wire [63:0] regs_258_io_in; // @[RegFile.scala 66:20:@41241.4]
  wire  regs_258_io_reset; // @[RegFile.scala 66:20:@41241.4]
  wire [63:0] regs_258_io_out; // @[RegFile.scala 66:20:@41241.4]
  wire  regs_258_io_enable; // @[RegFile.scala 66:20:@41241.4]
  wire  regs_259_clock; // @[RegFile.scala 66:20:@41255.4]
  wire  regs_259_reset; // @[RegFile.scala 66:20:@41255.4]
  wire [63:0] regs_259_io_in; // @[RegFile.scala 66:20:@41255.4]
  wire  regs_259_io_reset; // @[RegFile.scala 66:20:@41255.4]
  wire [63:0] regs_259_io_out; // @[RegFile.scala 66:20:@41255.4]
  wire  regs_259_io_enable; // @[RegFile.scala 66:20:@41255.4]
  wire  regs_260_clock; // @[RegFile.scala 66:20:@41269.4]
  wire  regs_260_reset; // @[RegFile.scala 66:20:@41269.4]
  wire [63:0] regs_260_io_in; // @[RegFile.scala 66:20:@41269.4]
  wire  regs_260_io_reset; // @[RegFile.scala 66:20:@41269.4]
  wire [63:0] regs_260_io_out; // @[RegFile.scala 66:20:@41269.4]
  wire  regs_260_io_enable; // @[RegFile.scala 66:20:@41269.4]
  wire  regs_261_clock; // @[RegFile.scala 66:20:@41283.4]
  wire  regs_261_reset; // @[RegFile.scala 66:20:@41283.4]
  wire [63:0] regs_261_io_in; // @[RegFile.scala 66:20:@41283.4]
  wire  regs_261_io_reset; // @[RegFile.scala 66:20:@41283.4]
  wire [63:0] regs_261_io_out; // @[RegFile.scala 66:20:@41283.4]
  wire  regs_261_io_enable; // @[RegFile.scala 66:20:@41283.4]
  wire  regs_262_clock; // @[RegFile.scala 66:20:@41297.4]
  wire  regs_262_reset; // @[RegFile.scala 66:20:@41297.4]
  wire [63:0] regs_262_io_in; // @[RegFile.scala 66:20:@41297.4]
  wire  regs_262_io_reset; // @[RegFile.scala 66:20:@41297.4]
  wire [63:0] regs_262_io_out; // @[RegFile.scala 66:20:@41297.4]
  wire  regs_262_io_enable; // @[RegFile.scala 66:20:@41297.4]
  wire  regs_263_clock; // @[RegFile.scala 66:20:@41311.4]
  wire  regs_263_reset; // @[RegFile.scala 66:20:@41311.4]
  wire [63:0] regs_263_io_in; // @[RegFile.scala 66:20:@41311.4]
  wire  regs_263_io_reset; // @[RegFile.scala 66:20:@41311.4]
  wire [63:0] regs_263_io_out; // @[RegFile.scala 66:20:@41311.4]
  wire  regs_263_io_enable; // @[RegFile.scala 66:20:@41311.4]
  wire  regs_264_clock; // @[RegFile.scala 66:20:@41325.4]
  wire  regs_264_reset; // @[RegFile.scala 66:20:@41325.4]
  wire [63:0] regs_264_io_in; // @[RegFile.scala 66:20:@41325.4]
  wire  regs_264_io_reset; // @[RegFile.scala 66:20:@41325.4]
  wire [63:0] regs_264_io_out; // @[RegFile.scala 66:20:@41325.4]
  wire  regs_264_io_enable; // @[RegFile.scala 66:20:@41325.4]
  wire  regs_265_clock; // @[RegFile.scala 66:20:@41339.4]
  wire  regs_265_reset; // @[RegFile.scala 66:20:@41339.4]
  wire [63:0] regs_265_io_in; // @[RegFile.scala 66:20:@41339.4]
  wire  regs_265_io_reset; // @[RegFile.scala 66:20:@41339.4]
  wire [63:0] regs_265_io_out; // @[RegFile.scala 66:20:@41339.4]
  wire  regs_265_io_enable; // @[RegFile.scala 66:20:@41339.4]
  wire  regs_266_clock; // @[RegFile.scala 66:20:@41353.4]
  wire  regs_266_reset; // @[RegFile.scala 66:20:@41353.4]
  wire [63:0] regs_266_io_in; // @[RegFile.scala 66:20:@41353.4]
  wire  regs_266_io_reset; // @[RegFile.scala 66:20:@41353.4]
  wire [63:0] regs_266_io_out; // @[RegFile.scala 66:20:@41353.4]
  wire  regs_266_io_enable; // @[RegFile.scala 66:20:@41353.4]
  wire  regs_267_clock; // @[RegFile.scala 66:20:@41367.4]
  wire  regs_267_reset; // @[RegFile.scala 66:20:@41367.4]
  wire [63:0] regs_267_io_in; // @[RegFile.scala 66:20:@41367.4]
  wire  regs_267_io_reset; // @[RegFile.scala 66:20:@41367.4]
  wire [63:0] regs_267_io_out; // @[RegFile.scala 66:20:@41367.4]
  wire  regs_267_io_enable; // @[RegFile.scala 66:20:@41367.4]
  wire  regs_268_clock; // @[RegFile.scala 66:20:@41381.4]
  wire  regs_268_reset; // @[RegFile.scala 66:20:@41381.4]
  wire [63:0] regs_268_io_in; // @[RegFile.scala 66:20:@41381.4]
  wire  regs_268_io_reset; // @[RegFile.scala 66:20:@41381.4]
  wire [63:0] regs_268_io_out; // @[RegFile.scala 66:20:@41381.4]
  wire  regs_268_io_enable; // @[RegFile.scala 66:20:@41381.4]
  wire  regs_269_clock; // @[RegFile.scala 66:20:@41395.4]
  wire  regs_269_reset; // @[RegFile.scala 66:20:@41395.4]
  wire [63:0] regs_269_io_in; // @[RegFile.scala 66:20:@41395.4]
  wire  regs_269_io_reset; // @[RegFile.scala 66:20:@41395.4]
  wire [63:0] regs_269_io_out; // @[RegFile.scala 66:20:@41395.4]
  wire  regs_269_io_enable; // @[RegFile.scala 66:20:@41395.4]
  wire  regs_270_clock; // @[RegFile.scala 66:20:@41409.4]
  wire  regs_270_reset; // @[RegFile.scala 66:20:@41409.4]
  wire [63:0] regs_270_io_in; // @[RegFile.scala 66:20:@41409.4]
  wire  regs_270_io_reset; // @[RegFile.scala 66:20:@41409.4]
  wire [63:0] regs_270_io_out; // @[RegFile.scala 66:20:@41409.4]
  wire  regs_270_io_enable; // @[RegFile.scala 66:20:@41409.4]
  wire  regs_271_clock; // @[RegFile.scala 66:20:@41423.4]
  wire  regs_271_reset; // @[RegFile.scala 66:20:@41423.4]
  wire [63:0] regs_271_io_in; // @[RegFile.scala 66:20:@41423.4]
  wire  regs_271_io_reset; // @[RegFile.scala 66:20:@41423.4]
  wire [63:0] regs_271_io_out; // @[RegFile.scala 66:20:@41423.4]
  wire  regs_271_io_enable; // @[RegFile.scala 66:20:@41423.4]
  wire  regs_272_clock; // @[RegFile.scala 66:20:@41437.4]
  wire  regs_272_reset; // @[RegFile.scala 66:20:@41437.4]
  wire [63:0] regs_272_io_in; // @[RegFile.scala 66:20:@41437.4]
  wire  regs_272_io_reset; // @[RegFile.scala 66:20:@41437.4]
  wire [63:0] regs_272_io_out; // @[RegFile.scala 66:20:@41437.4]
  wire  regs_272_io_enable; // @[RegFile.scala 66:20:@41437.4]
  wire  regs_273_clock; // @[RegFile.scala 66:20:@41451.4]
  wire  regs_273_reset; // @[RegFile.scala 66:20:@41451.4]
  wire [63:0] regs_273_io_in; // @[RegFile.scala 66:20:@41451.4]
  wire  regs_273_io_reset; // @[RegFile.scala 66:20:@41451.4]
  wire [63:0] regs_273_io_out; // @[RegFile.scala 66:20:@41451.4]
  wire  regs_273_io_enable; // @[RegFile.scala 66:20:@41451.4]
  wire  regs_274_clock; // @[RegFile.scala 66:20:@41465.4]
  wire  regs_274_reset; // @[RegFile.scala 66:20:@41465.4]
  wire [63:0] regs_274_io_in; // @[RegFile.scala 66:20:@41465.4]
  wire  regs_274_io_reset; // @[RegFile.scala 66:20:@41465.4]
  wire [63:0] regs_274_io_out; // @[RegFile.scala 66:20:@41465.4]
  wire  regs_274_io_enable; // @[RegFile.scala 66:20:@41465.4]
  wire  regs_275_clock; // @[RegFile.scala 66:20:@41479.4]
  wire  regs_275_reset; // @[RegFile.scala 66:20:@41479.4]
  wire [63:0] regs_275_io_in; // @[RegFile.scala 66:20:@41479.4]
  wire  regs_275_io_reset; // @[RegFile.scala 66:20:@41479.4]
  wire [63:0] regs_275_io_out; // @[RegFile.scala 66:20:@41479.4]
  wire  regs_275_io_enable; // @[RegFile.scala 66:20:@41479.4]
  wire  regs_276_clock; // @[RegFile.scala 66:20:@41493.4]
  wire  regs_276_reset; // @[RegFile.scala 66:20:@41493.4]
  wire [63:0] regs_276_io_in; // @[RegFile.scala 66:20:@41493.4]
  wire  regs_276_io_reset; // @[RegFile.scala 66:20:@41493.4]
  wire [63:0] regs_276_io_out; // @[RegFile.scala 66:20:@41493.4]
  wire  regs_276_io_enable; // @[RegFile.scala 66:20:@41493.4]
  wire  regs_277_clock; // @[RegFile.scala 66:20:@41507.4]
  wire  regs_277_reset; // @[RegFile.scala 66:20:@41507.4]
  wire [63:0] regs_277_io_in; // @[RegFile.scala 66:20:@41507.4]
  wire  regs_277_io_reset; // @[RegFile.scala 66:20:@41507.4]
  wire [63:0] regs_277_io_out; // @[RegFile.scala 66:20:@41507.4]
  wire  regs_277_io_enable; // @[RegFile.scala 66:20:@41507.4]
  wire  regs_278_clock; // @[RegFile.scala 66:20:@41521.4]
  wire  regs_278_reset; // @[RegFile.scala 66:20:@41521.4]
  wire [63:0] regs_278_io_in; // @[RegFile.scala 66:20:@41521.4]
  wire  regs_278_io_reset; // @[RegFile.scala 66:20:@41521.4]
  wire [63:0] regs_278_io_out; // @[RegFile.scala 66:20:@41521.4]
  wire  regs_278_io_enable; // @[RegFile.scala 66:20:@41521.4]
  wire  regs_279_clock; // @[RegFile.scala 66:20:@41535.4]
  wire  regs_279_reset; // @[RegFile.scala 66:20:@41535.4]
  wire [63:0] regs_279_io_in; // @[RegFile.scala 66:20:@41535.4]
  wire  regs_279_io_reset; // @[RegFile.scala 66:20:@41535.4]
  wire [63:0] regs_279_io_out; // @[RegFile.scala 66:20:@41535.4]
  wire  regs_279_io_enable; // @[RegFile.scala 66:20:@41535.4]
  wire  regs_280_clock; // @[RegFile.scala 66:20:@41549.4]
  wire  regs_280_reset; // @[RegFile.scala 66:20:@41549.4]
  wire [63:0] regs_280_io_in; // @[RegFile.scala 66:20:@41549.4]
  wire  regs_280_io_reset; // @[RegFile.scala 66:20:@41549.4]
  wire [63:0] regs_280_io_out; // @[RegFile.scala 66:20:@41549.4]
  wire  regs_280_io_enable; // @[RegFile.scala 66:20:@41549.4]
  wire  regs_281_clock; // @[RegFile.scala 66:20:@41563.4]
  wire  regs_281_reset; // @[RegFile.scala 66:20:@41563.4]
  wire [63:0] regs_281_io_in; // @[RegFile.scala 66:20:@41563.4]
  wire  regs_281_io_reset; // @[RegFile.scala 66:20:@41563.4]
  wire [63:0] regs_281_io_out; // @[RegFile.scala 66:20:@41563.4]
  wire  regs_281_io_enable; // @[RegFile.scala 66:20:@41563.4]
  wire  regs_282_clock; // @[RegFile.scala 66:20:@41577.4]
  wire  regs_282_reset; // @[RegFile.scala 66:20:@41577.4]
  wire [63:0] regs_282_io_in; // @[RegFile.scala 66:20:@41577.4]
  wire  regs_282_io_reset; // @[RegFile.scala 66:20:@41577.4]
  wire [63:0] regs_282_io_out; // @[RegFile.scala 66:20:@41577.4]
  wire  regs_282_io_enable; // @[RegFile.scala 66:20:@41577.4]
  wire  regs_283_clock; // @[RegFile.scala 66:20:@41591.4]
  wire  regs_283_reset; // @[RegFile.scala 66:20:@41591.4]
  wire [63:0] regs_283_io_in; // @[RegFile.scala 66:20:@41591.4]
  wire  regs_283_io_reset; // @[RegFile.scala 66:20:@41591.4]
  wire [63:0] regs_283_io_out; // @[RegFile.scala 66:20:@41591.4]
  wire  regs_283_io_enable; // @[RegFile.scala 66:20:@41591.4]
  wire  regs_284_clock; // @[RegFile.scala 66:20:@41605.4]
  wire  regs_284_reset; // @[RegFile.scala 66:20:@41605.4]
  wire [63:0] regs_284_io_in; // @[RegFile.scala 66:20:@41605.4]
  wire  regs_284_io_reset; // @[RegFile.scala 66:20:@41605.4]
  wire [63:0] regs_284_io_out; // @[RegFile.scala 66:20:@41605.4]
  wire  regs_284_io_enable; // @[RegFile.scala 66:20:@41605.4]
  wire  regs_285_clock; // @[RegFile.scala 66:20:@41619.4]
  wire  regs_285_reset; // @[RegFile.scala 66:20:@41619.4]
  wire [63:0] regs_285_io_in; // @[RegFile.scala 66:20:@41619.4]
  wire  regs_285_io_reset; // @[RegFile.scala 66:20:@41619.4]
  wire [63:0] regs_285_io_out; // @[RegFile.scala 66:20:@41619.4]
  wire  regs_285_io_enable; // @[RegFile.scala 66:20:@41619.4]
  wire  regs_286_clock; // @[RegFile.scala 66:20:@41633.4]
  wire  regs_286_reset; // @[RegFile.scala 66:20:@41633.4]
  wire [63:0] regs_286_io_in; // @[RegFile.scala 66:20:@41633.4]
  wire  regs_286_io_reset; // @[RegFile.scala 66:20:@41633.4]
  wire [63:0] regs_286_io_out; // @[RegFile.scala 66:20:@41633.4]
  wire  regs_286_io_enable; // @[RegFile.scala 66:20:@41633.4]
  wire  regs_287_clock; // @[RegFile.scala 66:20:@41647.4]
  wire  regs_287_reset; // @[RegFile.scala 66:20:@41647.4]
  wire [63:0] regs_287_io_in; // @[RegFile.scala 66:20:@41647.4]
  wire  regs_287_io_reset; // @[RegFile.scala 66:20:@41647.4]
  wire [63:0] regs_287_io_out; // @[RegFile.scala 66:20:@41647.4]
  wire  regs_287_io_enable; // @[RegFile.scala 66:20:@41647.4]
  wire  regs_288_clock; // @[RegFile.scala 66:20:@41661.4]
  wire  regs_288_reset; // @[RegFile.scala 66:20:@41661.4]
  wire [63:0] regs_288_io_in; // @[RegFile.scala 66:20:@41661.4]
  wire  regs_288_io_reset; // @[RegFile.scala 66:20:@41661.4]
  wire [63:0] regs_288_io_out; // @[RegFile.scala 66:20:@41661.4]
  wire  regs_288_io_enable; // @[RegFile.scala 66:20:@41661.4]
  wire  regs_289_clock; // @[RegFile.scala 66:20:@41675.4]
  wire  regs_289_reset; // @[RegFile.scala 66:20:@41675.4]
  wire [63:0] regs_289_io_in; // @[RegFile.scala 66:20:@41675.4]
  wire  regs_289_io_reset; // @[RegFile.scala 66:20:@41675.4]
  wire [63:0] regs_289_io_out; // @[RegFile.scala 66:20:@41675.4]
  wire  regs_289_io_enable; // @[RegFile.scala 66:20:@41675.4]
  wire  regs_290_clock; // @[RegFile.scala 66:20:@41689.4]
  wire  regs_290_reset; // @[RegFile.scala 66:20:@41689.4]
  wire [63:0] regs_290_io_in; // @[RegFile.scala 66:20:@41689.4]
  wire  regs_290_io_reset; // @[RegFile.scala 66:20:@41689.4]
  wire [63:0] regs_290_io_out; // @[RegFile.scala 66:20:@41689.4]
  wire  regs_290_io_enable; // @[RegFile.scala 66:20:@41689.4]
  wire  regs_291_clock; // @[RegFile.scala 66:20:@41703.4]
  wire  regs_291_reset; // @[RegFile.scala 66:20:@41703.4]
  wire [63:0] regs_291_io_in; // @[RegFile.scala 66:20:@41703.4]
  wire  regs_291_io_reset; // @[RegFile.scala 66:20:@41703.4]
  wire [63:0] regs_291_io_out; // @[RegFile.scala 66:20:@41703.4]
  wire  regs_291_io_enable; // @[RegFile.scala 66:20:@41703.4]
  wire  regs_292_clock; // @[RegFile.scala 66:20:@41717.4]
  wire  regs_292_reset; // @[RegFile.scala 66:20:@41717.4]
  wire [63:0] regs_292_io_in; // @[RegFile.scala 66:20:@41717.4]
  wire  regs_292_io_reset; // @[RegFile.scala 66:20:@41717.4]
  wire [63:0] regs_292_io_out; // @[RegFile.scala 66:20:@41717.4]
  wire  regs_292_io_enable; // @[RegFile.scala 66:20:@41717.4]
  wire  regs_293_clock; // @[RegFile.scala 66:20:@41731.4]
  wire  regs_293_reset; // @[RegFile.scala 66:20:@41731.4]
  wire [63:0] regs_293_io_in; // @[RegFile.scala 66:20:@41731.4]
  wire  regs_293_io_reset; // @[RegFile.scala 66:20:@41731.4]
  wire [63:0] regs_293_io_out; // @[RegFile.scala 66:20:@41731.4]
  wire  regs_293_io_enable; // @[RegFile.scala 66:20:@41731.4]
  wire  regs_294_clock; // @[RegFile.scala 66:20:@41745.4]
  wire  regs_294_reset; // @[RegFile.scala 66:20:@41745.4]
  wire [63:0] regs_294_io_in; // @[RegFile.scala 66:20:@41745.4]
  wire  regs_294_io_reset; // @[RegFile.scala 66:20:@41745.4]
  wire [63:0] regs_294_io_out; // @[RegFile.scala 66:20:@41745.4]
  wire  regs_294_io_enable; // @[RegFile.scala 66:20:@41745.4]
  wire  regs_295_clock; // @[RegFile.scala 66:20:@41759.4]
  wire  regs_295_reset; // @[RegFile.scala 66:20:@41759.4]
  wire [63:0] regs_295_io_in; // @[RegFile.scala 66:20:@41759.4]
  wire  regs_295_io_reset; // @[RegFile.scala 66:20:@41759.4]
  wire [63:0] regs_295_io_out; // @[RegFile.scala 66:20:@41759.4]
  wire  regs_295_io_enable; // @[RegFile.scala 66:20:@41759.4]
  wire  regs_296_clock; // @[RegFile.scala 66:20:@41773.4]
  wire  regs_296_reset; // @[RegFile.scala 66:20:@41773.4]
  wire [63:0] regs_296_io_in; // @[RegFile.scala 66:20:@41773.4]
  wire  regs_296_io_reset; // @[RegFile.scala 66:20:@41773.4]
  wire [63:0] regs_296_io_out; // @[RegFile.scala 66:20:@41773.4]
  wire  regs_296_io_enable; // @[RegFile.scala 66:20:@41773.4]
  wire  regs_297_clock; // @[RegFile.scala 66:20:@41787.4]
  wire  regs_297_reset; // @[RegFile.scala 66:20:@41787.4]
  wire [63:0] regs_297_io_in; // @[RegFile.scala 66:20:@41787.4]
  wire  regs_297_io_reset; // @[RegFile.scala 66:20:@41787.4]
  wire [63:0] regs_297_io_out; // @[RegFile.scala 66:20:@41787.4]
  wire  regs_297_io_enable; // @[RegFile.scala 66:20:@41787.4]
  wire  regs_298_clock; // @[RegFile.scala 66:20:@41801.4]
  wire  regs_298_reset; // @[RegFile.scala 66:20:@41801.4]
  wire [63:0] regs_298_io_in; // @[RegFile.scala 66:20:@41801.4]
  wire  regs_298_io_reset; // @[RegFile.scala 66:20:@41801.4]
  wire [63:0] regs_298_io_out; // @[RegFile.scala 66:20:@41801.4]
  wire  regs_298_io_enable; // @[RegFile.scala 66:20:@41801.4]
  wire  regs_299_clock; // @[RegFile.scala 66:20:@41815.4]
  wire  regs_299_reset; // @[RegFile.scala 66:20:@41815.4]
  wire [63:0] regs_299_io_in; // @[RegFile.scala 66:20:@41815.4]
  wire  regs_299_io_reset; // @[RegFile.scala 66:20:@41815.4]
  wire [63:0] regs_299_io_out; // @[RegFile.scala 66:20:@41815.4]
  wire  regs_299_io_enable; // @[RegFile.scala 66:20:@41815.4]
  wire  regs_300_clock; // @[RegFile.scala 66:20:@41829.4]
  wire  regs_300_reset; // @[RegFile.scala 66:20:@41829.4]
  wire [63:0] regs_300_io_in; // @[RegFile.scala 66:20:@41829.4]
  wire  regs_300_io_reset; // @[RegFile.scala 66:20:@41829.4]
  wire [63:0] regs_300_io_out; // @[RegFile.scala 66:20:@41829.4]
  wire  regs_300_io_enable; // @[RegFile.scala 66:20:@41829.4]
  wire  regs_301_clock; // @[RegFile.scala 66:20:@41843.4]
  wire  regs_301_reset; // @[RegFile.scala 66:20:@41843.4]
  wire [63:0] regs_301_io_in; // @[RegFile.scala 66:20:@41843.4]
  wire  regs_301_io_reset; // @[RegFile.scala 66:20:@41843.4]
  wire [63:0] regs_301_io_out; // @[RegFile.scala 66:20:@41843.4]
  wire  regs_301_io_enable; // @[RegFile.scala 66:20:@41843.4]
  wire  regs_302_clock; // @[RegFile.scala 66:20:@41857.4]
  wire  regs_302_reset; // @[RegFile.scala 66:20:@41857.4]
  wire [63:0] regs_302_io_in; // @[RegFile.scala 66:20:@41857.4]
  wire  regs_302_io_reset; // @[RegFile.scala 66:20:@41857.4]
  wire [63:0] regs_302_io_out; // @[RegFile.scala 66:20:@41857.4]
  wire  regs_302_io_enable; // @[RegFile.scala 66:20:@41857.4]
  wire  regs_303_clock; // @[RegFile.scala 66:20:@41871.4]
  wire  regs_303_reset; // @[RegFile.scala 66:20:@41871.4]
  wire [63:0] regs_303_io_in; // @[RegFile.scala 66:20:@41871.4]
  wire  regs_303_io_reset; // @[RegFile.scala 66:20:@41871.4]
  wire [63:0] regs_303_io_out; // @[RegFile.scala 66:20:@41871.4]
  wire  regs_303_io_enable; // @[RegFile.scala 66:20:@41871.4]
  wire  regs_304_clock; // @[RegFile.scala 66:20:@41885.4]
  wire  regs_304_reset; // @[RegFile.scala 66:20:@41885.4]
  wire [63:0] regs_304_io_in; // @[RegFile.scala 66:20:@41885.4]
  wire  regs_304_io_reset; // @[RegFile.scala 66:20:@41885.4]
  wire [63:0] regs_304_io_out; // @[RegFile.scala 66:20:@41885.4]
  wire  regs_304_io_enable; // @[RegFile.scala 66:20:@41885.4]
  wire  regs_305_clock; // @[RegFile.scala 66:20:@41899.4]
  wire  regs_305_reset; // @[RegFile.scala 66:20:@41899.4]
  wire [63:0] regs_305_io_in; // @[RegFile.scala 66:20:@41899.4]
  wire  regs_305_io_reset; // @[RegFile.scala 66:20:@41899.4]
  wire [63:0] regs_305_io_out; // @[RegFile.scala 66:20:@41899.4]
  wire  regs_305_io_enable; // @[RegFile.scala 66:20:@41899.4]
  wire  regs_306_clock; // @[RegFile.scala 66:20:@41913.4]
  wire  regs_306_reset; // @[RegFile.scala 66:20:@41913.4]
  wire [63:0] regs_306_io_in; // @[RegFile.scala 66:20:@41913.4]
  wire  regs_306_io_reset; // @[RegFile.scala 66:20:@41913.4]
  wire [63:0] regs_306_io_out; // @[RegFile.scala 66:20:@41913.4]
  wire  regs_306_io_enable; // @[RegFile.scala 66:20:@41913.4]
  wire  regs_307_clock; // @[RegFile.scala 66:20:@41927.4]
  wire  regs_307_reset; // @[RegFile.scala 66:20:@41927.4]
  wire [63:0] regs_307_io_in; // @[RegFile.scala 66:20:@41927.4]
  wire  regs_307_io_reset; // @[RegFile.scala 66:20:@41927.4]
  wire [63:0] regs_307_io_out; // @[RegFile.scala 66:20:@41927.4]
  wire  regs_307_io_enable; // @[RegFile.scala 66:20:@41927.4]
  wire  regs_308_clock; // @[RegFile.scala 66:20:@41941.4]
  wire  regs_308_reset; // @[RegFile.scala 66:20:@41941.4]
  wire [63:0] regs_308_io_in; // @[RegFile.scala 66:20:@41941.4]
  wire  regs_308_io_reset; // @[RegFile.scala 66:20:@41941.4]
  wire [63:0] regs_308_io_out; // @[RegFile.scala 66:20:@41941.4]
  wire  regs_308_io_enable; // @[RegFile.scala 66:20:@41941.4]
  wire  regs_309_clock; // @[RegFile.scala 66:20:@41955.4]
  wire  regs_309_reset; // @[RegFile.scala 66:20:@41955.4]
  wire [63:0] regs_309_io_in; // @[RegFile.scala 66:20:@41955.4]
  wire  regs_309_io_reset; // @[RegFile.scala 66:20:@41955.4]
  wire [63:0] regs_309_io_out; // @[RegFile.scala 66:20:@41955.4]
  wire  regs_309_io_enable; // @[RegFile.scala 66:20:@41955.4]
  wire  regs_310_clock; // @[RegFile.scala 66:20:@41969.4]
  wire  regs_310_reset; // @[RegFile.scala 66:20:@41969.4]
  wire [63:0] regs_310_io_in; // @[RegFile.scala 66:20:@41969.4]
  wire  regs_310_io_reset; // @[RegFile.scala 66:20:@41969.4]
  wire [63:0] regs_310_io_out; // @[RegFile.scala 66:20:@41969.4]
  wire  regs_310_io_enable; // @[RegFile.scala 66:20:@41969.4]
  wire  regs_311_clock; // @[RegFile.scala 66:20:@41983.4]
  wire  regs_311_reset; // @[RegFile.scala 66:20:@41983.4]
  wire [63:0] regs_311_io_in; // @[RegFile.scala 66:20:@41983.4]
  wire  regs_311_io_reset; // @[RegFile.scala 66:20:@41983.4]
  wire [63:0] regs_311_io_out; // @[RegFile.scala 66:20:@41983.4]
  wire  regs_311_io_enable; // @[RegFile.scala 66:20:@41983.4]
  wire  regs_312_clock; // @[RegFile.scala 66:20:@41997.4]
  wire  regs_312_reset; // @[RegFile.scala 66:20:@41997.4]
  wire [63:0] regs_312_io_in; // @[RegFile.scala 66:20:@41997.4]
  wire  regs_312_io_reset; // @[RegFile.scala 66:20:@41997.4]
  wire [63:0] regs_312_io_out; // @[RegFile.scala 66:20:@41997.4]
  wire  regs_312_io_enable; // @[RegFile.scala 66:20:@41997.4]
  wire  regs_313_clock; // @[RegFile.scala 66:20:@42011.4]
  wire  regs_313_reset; // @[RegFile.scala 66:20:@42011.4]
  wire [63:0] regs_313_io_in; // @[RegFile.scala 66:20:@42011.4]
  wire  regs_313_io_reset; // @[RegFile.scala 66:20:@42011.4]
  wire [63:0] regs_313_io_out; // @[RegFile.scala 66:20:@42011.4]
  wire  regs_313_io_enable; // @[RegFile.scala 66:20:@42011.4]
  wire  regs_314_clock; // @[RegFile.scala 66:20:@42025.4]
  wire  regs_314_reset; // @[RegFile.scala 66:20:@42025.4]
  wire [63:0] regs_314_io_in; // @[RegFile.scala 66:20:@42025.4]
  wire  regs_314_io_reset; // @[RegFile.scala 66:20:@42025.4]
  wire [63:0] regs_314_io_out; // @[RegFile.scala 66:20:@42025.4]
  wire  regs_314_io_enable; // @[RegFile.scala 66:20:@42025.4]
  wire  regs_315_clock; // @[RegFile.scala 66:20:@42039.4]
  wire  regs_315_reset; // @[RegFile.scala 66:20:@42039.4]
  wire [63:0] regs_315_io_in; // @[RegFile.scala 66:20:@42039.4]
  wire  regs_315_io_reset; // @[RegFile.scala 66:20:@42039.4]
  wire [63:0] regs_315_io_out; // @[RegFile.scala 66:20:@42039.4]
  wire  regs_315_io_enable; // @[RegFile.scala 66:20:@42039.4]
  wire  regs_316_clock; // @[RegFile.scala 66:20:@42053.4]
  wire  regs_316_reset; // @[RegFile.scala 66:20:@42053.4]
  wire [63:0] regs_316_io_in; // @[RegFile.scala 66:20:@42053.4]
  wire  regs_316_io_reset; // @[RegFile.scala 66:20:@42053.4]
  wire [63:0] regs_316_io_out; // @[RegFile.scala 66:20:@42053.4]
  wire  regs_316_io_enable; // @[RegFile.scala 66:20:@42053.4]
  wire  regs_317_clock; // @[RegFile.scala 66:20:@42067.4]
  wire  regs_317_reset; // @[RegFile.scala 66:20:@42067.4]
  wire [63:0] regs_317_io_in; // @[RegFile.scala 66:20:@42067.4]
  wire  regs_317_io_reset; // @[RegFile.scala 66:20:@42067.4]
  wire [63:0] regs_317_io_out; // @[RegFile.scala 66:20:@42067.4]
  wire  regs_317_io_enable; // @[RegFile.scala 66:20:@42067.4]
  wire  regs_318_clock; // @[RegFile.scala 66:20:@42081.4]
  wire  regs_318_reset; // @[RegFile.scala 66:20:@42081.4]
  wire [63:0] regs_318_io_in; // @[RegFile.scala 66:20:@42081.4]
  wire  regs_318_io_reset; // @[RegFile.scala 66:20:@42081.4]
  wire [63:0] regs_318_io_out; // @[RegFile.scala 66:20:@42081.4]
  wire  regs_318_io_enable; // @[RegFile.scala 66:20:@42081.4]
  wire  regs_319_clock; // @[RegFile.scala 66:20:@42095.4]
  wire  regs_319_reset; // @[RegFile.scala 66:20:@42095.4]
  wire [63:0] regs_319_io_in; // @[RegFile.scala 66:20:@42095.4]
  wire  regs_319_io_reset; // @[RegFile.scala 66:20:@42095.4]
  wire [63:0] regs_319_io_out; // @[RegFile.scala 66:20:@42095.4]
  wire  regs_319_io_enable; // @[RegFile.scala 66:20:@42095.4]
  wire  regs_320_clock; // @[RegFile.scala 66:20:@42109.4]
  wire  regs_320_reset; // @[RegFile.scala 66:20:@42109.4]
  wire [63:0] regs_320_io_in; // @[RegFile.scala 66:20:@42109.4]
  wire  regs_320_io_reset; // @[RegFile.scala 66:20:@42109.4]
  wire [63:0] regs_320_io_out; // @[RegFile.scala 66:20:@42109.4]
  wire  regs_320_io_enable; // @[RegFile.scala 66:20:@42109.4]
  wire  regs_321_clock; // @[RegFile.scala 66:20:@42123.4]
  wire  regs_321_reset; // @[RegFile.scala 66:20:@42123.4]
  wire [63:0] regs_321_io_in; // @[RegFile.scala 66:20:@42123.4]
  wire  regs_321_io_reset; // @[RegFile.scala 66:20:@42123.4]
  wire [63:0] regs_321_io_out; // @[RegFile.scala 66:20:@42123.4]
  wire  regs_321_io_enable; // @[RegFile.scala 66:20:@42123.4]
  wire  regs_322_clock; // @[RegFile.scala 66:20:@42137.4]
  wire  regs_322_reset; // @[RegFile.scala 66:20:@42137.4]
  wire [63:0] regs_322_io_in; // @[RegFile.scala 66:20:@42137.4]
  wire  regs_322_io_reset; // @[RegFile.scala 66:20:@42137.4]
  wire [63:0] regs_322_io_out; // @[RegFile.scala 66:20:@42137.4]
  wire  regs_322_io_enable; // @[RegFile.scala 66:20:@42137.4]
  wire  regs_323_clock; // @[RegFile.scala 66:20:@42151.4]
  wire  regs_323_reset; // @[RegFile.scala 66:20:@42151.4]
  wire [63:0] regs_323_io_in; // @[RegFile.scala 66:20:@42151.4]
  wire  regs_323_io_reset; // @[RegFile.scala 66:20:@42151.4]
  wire [63:0] regs_323_io_out; // @[RegFile.scala 66:20:@42151.4]
  wire  regs_323_io_enable; // @[RegFile.scala 66:20:@42151.4]
  wire  regs_324_clock; // @[RegFile.scala 66:20:@42165.4]
  wire  regs_324_reset; // @[RegFile.scala 66:20:@42165.4]
  wire [63:0] regs_324_io_in; // @[RegFile.scala 66:20:@42165.4]
  wire  regs_324_io_reset; // @[RegFile.scala 66:20:@42165.4]
  wire [63:0] regs_324_io_out; // @[RegFile.scala 66:20:@42165.4]
  wire  regs_324_io_enable; // @[RegFile.scala 66:20:@42165.4]
  wire  regs_325_clock; // @[RegFile.scala 66:20:@42179.4]
  wire  regs_325_reset; // @[RegFile.scala 66:20:@42179.4]
  wire [63:0] regs_325_io_in; // @[RegFile.scala 66:20:@42179.4]
  wire  regs_325_io_reset; // @[RegFile.scala 66:20:@42179.4]
  wire [63:0] regs_325_io_out; // @[RegFile.scala 66:20:@42179.4]
  wire  regs_325_io_enable; // @[RegFile.scala 66:20:@42179.4]
  wire  regs_326_clock; // @[RegFile.scala 66:20:@42193.4]
  wire  regs_326_reset; // @[RegFile.scala 66:20:@42193.4]
  wire [63:0] regs_326_io_in; // @[RegFile.scala 66:20:@42193.4]
  wire  regs_326_io_reset; // @[RegFile.scala 66:20:@42193.4]
  wire [63:0] regs_326_io_out; // @[RegFile.scala 66:20:@42193.4]
  wire  regs_326_io_enable; // @[RegFile.scala 66:20:@42193.4]
  wire  regs_327_clock; // @[RegFile.scala 66:20:@42207.4]
  wire  regs_327_reset; // @[RegFile.scala 66:20:@42207.4]
  wire [63:0] regs_327_io_in; // @[RegFile.scala 66:20:@42207.4]
  wire  regs_327_io_reset; // @[RegFile.scala 66:20:@42207.4]
  wire [63:0] regs_327_io_out; // @[RegFile.scala 66:20:@42207.4]
  wire  regs_327_io_enable; // @[RegFile.scala 66:20:@42207.4]
  wire  regs_328_clock; // @[RegFile.scala 66:20:@42221.4]
  wire  regs_328_reset; // @[RegFile.scala 66:20:@42221.4]
  wire [63:0] regs_328_io_in; // @[RegFile.scala 66:20:@42221.4]
  wire  regs_328_io_reset; // @[RegFile.scala 66:20:@42221.4]
  wire [63:0] regs_328_io_out; // @[RegFile.scala 66:20:@42221.4]
  wire  regs_328_io_enable; // @[RegFile.scala 66:20:@42221.4]
  wire  regs_329_clock; // @[RegFile.scala 66:20:@42235.4]
  wire  regs_329_reset; // @[RegFile.scala 66:20:@42235.4]
  wire [63:0] regs_329_io_in; // @[RegFile.scala 66:20:@42235.4]
  wire  regs_329_io_reset; // @[RegFile.scala 66:20:@42235.4]
  wire [63:0] regs_329_io_out; // @[RegFile.scala 66:20:@42235.4]
  wire  regs_329_io_enable; // @[RegFile.scala 66:20:@42235.4]
  wire  regs_330_clock; // @[RegFile.scala 66:20:@42249.4]
  wire  regs_330_reset; // @[RegFile.scala 66:20:@42249.4]
  wire [63:0] regs_330_io_in; // @[RegFile.scala 66:20:@42249.4]
  wire  regs_330_io_reset; // @[RegFile.scala 66:20:@42249.4]
  wire [63:0] regs_330_io_out; // @[RegFile.scala 66:20:@42249.4]
  wire  regs_330_io_enable; // @[RegFile.scala 66:20:@42249.4]
  wire  regs_331_clock; // @[RegFile.scala 66:20:@42263.4]
  wire  regs_331_reset; // @[RegFile.scala 66:20:@42263.4]
  wire [63:0] regs_331_io_in; // @[RegFile.scala 66:20:@42263.4]
  wire  regs_331_io_reset; // @[RegFile.scala 66:20:@42263.4]
  wire [63:0] regs_331_io_out; // @[RegFile.scala 66:20:@42263.4]
  wire  regs_331_io_enable; // @[RegFile.scala 66:20:@42263.4]
  wire  regs_332_clock; // @[RegFile.scala 66:20:@42277.4]
  wire  regs_332_reset; // @[RegFile.scala 66:20:@42277.4]
  wire [63:0] regs_332_io_in; // @[RegFile.scala 66:20:@42277.4]
  wire  regs_332_io_reset; // @[RegFile.scala 66:20:@42277.4]
  wire [63:0] regs_332_io_out; // @[RegFile.scala 66:20:@42277.4]
  wire  regs_332_io_enable; // @[RegFile.scala 66:20:@42277.4]
  wire  regs_333_clock; // @[RegFile.scala 66:20:@42291.4]
  wire  regs_333_reset; // @[RegFile.scala 66:20:@42291.4]
  wire [63:0] regs_333_io_in; // @[RegFile.scala 66:20:@42291.4]
  wire  regs_333_io_reset; // @[RegFile.scala 66:20:@42291.4]
  wire [63:0] regs_333_io_out; // @[RegFile.scala 66:20:@42291.4]
  wire  regs_333_io_enable; // @[RegFile.scala 66:20:@42291.4]
  wire  regs_334_clock; // @[RegFile.scala 66:20:@42305.4]
  wire  regs_334_reset; // @[RegFile.scala 66:20:@42305.4]
  wire [63:0] regs_334_io_in; // @[RegFile.scala 66:20:@42305.4]
  wire  regs_334_io_reset; // @[RegFile.scala 66:20:@42305.4]
  wire [63:0] regs_334_io_out; // @[RegFile.scala 66:20:@42305.4]
  wire  regs_334_io_enable; // @[RegFile.scala 66:20:@42305.4]
  wire  regs_335_clock; // @[RegFile.scala 66:20:@42319.4]
  wire  regs_335_reset; // @[RegFile.scala 66:20:@42319.4]
  wire [63:0] regs_335_io_in; // @[RegFile.scala 66:20:@42319.4]
  wire  regs_335_io_reset; // @[RegFile.scala 66:20:@42319.4]
  wire [63:0] regs_335_io_out; // @[RegFile.scala 66:20:@42319.4]
  wire  regs_335_io_enable; // @[RegFile.scala 66:20:@42319.4]
  wire  regs_336_clock; // @[RegFile.scala 66:20:@42333.4]
  wire  regs_336_reset; // @[RegFile.scala 66:20:@42333.4]
  wire [63:0] regs_336_io_in; // @[RegFile.scala 66:20:@42333.4]
  wire  regs_336_io_reset; // @[RegFile.scala 66:20:@42333.4]
  wire [63:0] regs_336_io_out; // @[RegFile.scala 66:20:@42333.4]
  wire  regs_336_io_enable; // @[RegFile.scala 66:20:@42333.4]
  wire  regs_337_clock; // @[RegFile.scala 66:20:@42347.4]
  wire  regs_337_reset; // @[RegFile.scala 66:20:@42347.4]
  wire [63:0] regs_337_io_in; // @[RegFile.scala 66:20:@42347.4]
  wire  regs_337_io_reset; // @[RegFile.scala 66:20:@42347.4]
  wire [63:0] regs_337_io_out; // @[RegFile.scala 66:20:@42347.4]
  wire  regs_337_io_enable; // @[RegFile.scala 66:20:@42347.4]
  wire  regs_338_clock; // @[RegFile.scala 66:20:@42361.4]
  wire  regs_338_reset; // @[RegFile.scala 66:20:@42361.4]
  wire [63:0] regs_338_io_in; // @[RegFile.scala 66:20:@42361.4]
  wire  regs_338_io_reset; // @[RegFile.scala 66:20:@42361.4]
  wire [63:0] regs_338_io_out; // @[RegFile.scala 66:20:@42361.4]
  wire  regs_338_io_enable; // @[RegFile.scala 66:20:@42361.4]
  wire  regs_339_clock; // @[RegFile.scala 66:20:@42375.4]
  wire  regs_339_reset; // @[RegFile.scala 66:20:@42375.4]
  wire [63:0] regs_339_io_in; // @[RegFile.scala 66:20:@42375.4]
  wire  regs_339_io_reset; // @[RegFile.scala 66:20:@42375.4]
  wire [63:0] regs_339_io_out; // @[RegFile.scala 66:20:@42375.4]
  wire  regs_339_io_enable; // @[RegFile.scala 66:20:@42375.4]
  wire  regs_340_clock; // @[RegFile.scala 66:20:@42389.4]
  wire  regs_340_reset; // @[RegFile.scala 66:20:@42389.4]
  wire [63:0] regs_340_io_in; // @[RegFile.scala 66:20:@42389.4]
  wire  regs_340_io_reset; // @[RegFile.scala 66:20:@42389.4]
  wire [63:0] regs_340_io_out; // @[RegFile.scala 66:20:@42389.4]
  wire  regs_340_io_enable; // @[RegFile.scala 66:20:@42389.4]
  wire  regs_341_clock; // @[RegFile.scala 66:20:@42403.4]
  wire  regs_341_reset; // @[RegFile.scala 66:20:@42403.4]
  wire [63:0] regs_341_io_in; // @[RegFile.scala 66:20:@42403.4]
  wire  regs_341_io_reset; // @[RegFile.scala 66:20:@42403.4]
  wire [63:0] regs_341_io_out; // @[RegFile.scala 66:20:@42403.4]
  wire  regs_341_io_enable; // @[RegFile.scala 66:20:@42403.4]
  wire  regs_342_clock; // @[RegFile.scala 66:20:@42417.4]
  wire  regs_342_reset; // @[RegFile.scala 66:20:@42417.4]
  wire [63:0] regs_342_io_in; // @[RegFile.scala 66:20:@42417.4]
  wire  regs_342_io_reset; // @[RegFile.scala 66:20:@42417.4]
  wire [63:0] regs_342_io_out; // @[RegFile.scala 66:20:@42417.4]
  wire  regs_342_io_enable; // @[RegFile.scala 66:20:@42417.4]
  wire  regs_343_clock; // @[RegFile.scala 66:20:@42431.4]
  wire  regs_343_reset; // @[RegFile.scala 66:20:@42431.4]
  wire [63:0] regs_343_io_in; // @[RegFile.scala 66:20:@42431.4]
  wire  regs_343_io_reset; // @[RegFile.scala 66:20:@42431.4]
  wire [63:0] regs_343_io_out; // @[RegFile.scala 66:20:@42431.4]
  wire  regs_343_io_enable; // @[RegFile.scala 66:20:@42431.4]
  wire  regs_344_clock; // @[RegFile.scala 66:20:@42445.4]
  wire  regs_344_reset; // @[RegFile.scala 66:20:@42445.4]
  wire [63:0] regs_344_io_in; // @[RegFile.scala 66:20:@42445.4]
  wire  regs_344_io_reset; // @[RegFile.scala 66:20:@42445.4]
  wire [63:0] regs_344_io_out; // @[RegFile.scala 66:20:@42445.4]
  wire  regs_344_io_enable; // @[RegFile.scala 66:20:@42445.4]
  wire  regs_345_clock; // @[RegFile.scala 66:20:@42459.4]
  wire  regs_345_reset; // @[RegFile.scala 66:20:@42459.4]
  wire [63:0] regs_345_io_in; // @[RegFile.scala 66:20:@42459.4]
  wire  regs_345_io_reset; // @[RegFile.scala 66:20:@42459.4]
  wire [63:0] regs_345_io_out; // @[RegFile.scala 66:20:@42459.4]
  wire  regs_345_io_enable; // @[RegFile.scala 66:20:@42459.4]
  wire  regs_346_clock; // @[RegFile.scala 66:20:@42473.4]
  wire  regs_346_reset; // @[RegFile.scala 66:20:@42473.4]
  wire [63:0] regs_346_io_in; // @[RegFile.scala 66:20:@42473.4]
  wire  regs_346_io_reset; // @[RegFile.scala 66:20:@42473.4]
  wire [63:0] regs_346_io_out; // @[RegFile.scala 66:20:@42473.4]
  wire  regs_346_io_enable; // @[RegFile.scala 66:20:@42473.4]
  wire  regs_347_clock; // @[RegFile.scala 66:20:@42487.4]
  wire  regs_347_reset; // @[RegFile.scala 66:20:@42487.4]
  wire [63:0] regs_347_io_in; // @[RegFile.scala 66:20:@42487.4]
  wire  regs_347_io_reset; // @[RegFile.scala 66:20:@42487.4]
  wire [63:0] regs_347_io_out; // @[RegFile.scala 66:20:@42487.4]
  wire  regs_347_io_enable; // @[RegFile.scala 66:20:@42487.4]
  wire  regs_348_clock; // @[RegFile.scala 66:20:@42501.4]
  wire  regs_348_reset; // @[RegFile.scala 66:20:@42501.4]
  wire [63:0] regs_348_io_in; // @[RegFile.scala 66:20:@42501.4]
  wire  regs_348_io_reset; // @[RegFile.scala 66:20:@42501.4]
  wire [63:0] regs_348_io_out; // @[RegFile.scala 66:20:@42501.4]
  wire  regs_348_io_enable; // @[RegFile.scala 66:20:@42501.4]
  wire  regs_349_clock; // @[RegFile.scala 66:20:@42515.4]
  wire  regs_349_reset; // @[RegFile.scala 66:20:@42515.4]
  wire [63:0] regs_349_io_in; // @[RegFile.scala 66:20:@42515.4]
  wire  regs_349_io_reset; // @[RegFile.scala 66:20:@42515.4]
  wire [63:0] regs_349_io_out; // @[RegFile.scala 66:20:@42515.4]
  wire  regs_349_io_enable; // @[RegFile.scala 66:20:@42515.4]
  wire  regs_350_clock; // @[RegFile.scala 66:20:@42529.4]
  wire  regs_350_reset; // @[RegFile.scala 66:20:@42529.4]
  wire [63:0] regs_350_io_in; // @[RegFile.scala 66:20:@42529.4]
  wire  regs_350_io_reset; // @[RegFile.scala 66:20:@42529.4]
  wire [63:0] regs_350_io_out; // @[RegFile.scala 66:20:@42529.4]
  wire  regs_350_io_enable; // @[RegFile.scala 66:20:@42529.4]
  wire  regs_351_clock; // @[RegFile.scala 66:20:@42543.4]
  wire  regs_351_reset; // @[RegFile.scala 66:20:@42543.4]
  wire [63:0] regs_351_io_in; // @[RegFile.scala 66:20:@42543.4]
  wire  regs_351_io_reset; // @[RegFile.scala 66:20:@42543.4]
  wire [63:0] regs_351_io_out; // @[RegFile.scala 66:20:@42543.4]
  wire  regs_351_io_enable; // @[RegFile.scala 66:20:@42543.4]
  wire  regs_352_clock; // @[RegFile.scala 66:20:@42557.4]
  wire  regs_352_reset; // @[RegFile.scala 66:20:@42557.4]
  wire [63:0] regs_352_io_in; // @[RegFile.scala 66:20:@42557.4]
  wire  regs_352_io_reset; // @[RegFile.scala 66:20:@42557.4]
  wire [63:0] regs_352_io_out; // @[RegFile.scala 66:20:@42557.4]
  wire  regs_352_io_enable; // @[RegFile.scala 66:20:@42557.4]
  wire  regs_353_clock; // @[RegFile.scala 66:20:@42571.4]
  wire  regs_353_reset; // @[RegFile.scala 66:20:@42571.4]
  wire [63:0] regs_353_io_in; // @[RegFile.scala 66:20:@42571.4]
  wire  regs_353_io_reset; // @[RegFile.scala 66:20:@42571.4]
  wire [63:0] regs_353_io_out; // @[RegFile.scala 66:20:@42571.4]
  wire  regs_353_io_enable; // @[RegFile.scala 66:20:@42571.4]
  wire  regs_354_clock; // @[RegFile.scala 66:20:@42585.4]
  wire  regs_354_reset; // @[RegFile.scala 66:20:@42585.4]
  wire [63:0] regs_354_io_in; // @[RegFile.scala 66:20:@42585.4]
  wire  regs_354_io_reset; // @[RegFile.scala 66:20:@42585.4]
  wire [63:0] regs_354_io_out; // @[RegFile.scala 66:20:@42585.4]
  wire  regs_354_io_enable; // @[RegFile.scala 66:20:@42585.4]
  wire  regs_355_clock; // @[RegFile.scala 66:20:@42599.4]
  wire  regs_355_reset; // @[RegFile.scala 66:20:@42599.4]
  wire [63:0] regs_355_io_in; // @[RegFile.scala 66:20:@42599.4]
  wire  regs_355_io_reset; // @[RegFile.scala 66:20:@42599.4]
  wire [63:0] regs_355_io_out; // @[RegFile.scala 66:20:@42599.4]
  wire  regs_355_io_enable; // @[RegFile.scala 66:20:@42599.4]
  wire  regs_356_clock; // @[RegFile.scala 66:20:@42613.4]
  wire  regs_356_reset; // @[RegFile.scala 66:20:@42613.4]
  wire [63:0] regs_356_io_in; // @[RegFile.scala 66:20:@42613.4]
  wire  regs_356_io_reset; // @[RegFile.scala 66:20:@42613.4]
  wire [63:0] regs_356_io_out; // @[RegFile.scala 66:20:@42613.4]
  wire  regs_356_io_enable; // @[RegFile.scala 66:20:@42613.4]
  wire  regs_357_clock; // @[RegFile.scala 66:20:@42627.4]
  wire  regs_357_reset; // @[RegFile.scala 66:20:@42627.4]
  wire [63:0] regs_357_io_in; // @[RegFile.scala 66:20:@42627.4]
  wire  regs_357_io_reset; // @[RegFile.scala 66:20:@42627.4]
  wire [63:0] regs_357_io_out; // @[RegFile.scala 66:20:@42627.4]
  wire  regs_357_io_enable; // @[RegFile.scala 66:20:@42627.4]
  wire  regs_358_clock; // @[RegFile.scala 66:20:@42641.4]
  wire  regs_358_reset; // @[RegFile.scala 66:20:@42641.4]
  wire [63:0] regs_358_io_in; // @[RegFile.scala 66:20:@42641.4]
  wire  regs_358_io_reset; // @[RegFile.scala 66:20:@42641.4]
  wire [63:0] regs_358_io_out; // @[RegFile.scala 66:20:@42641.4]
  wire  regs_358_io_enable; // @[RegFile.scala 66:20:@42641.4]
  wire  regs_359_clock; // @[RegFile.scala 66:20:@42655.4]
  wire  regs_359_reset; // @[RegFile.scala 66:20:@42655.4]
  wire [63:0] regs_359_io_in; // @[RegFile.scala 66:20:@42655.4]
  wire  regs_359_io_reset; // @[RegFile.scala 66:20:@42655.4]
  wire [63:0] regs_359_io_out; // @[RegFile.scala 66:20:@42655.4]
  wire  regs_359_io_enable; // @[RegFile.scala 66:20:@42655.4]
  wire  regs_360_clock; // @[RegFile.scala 66:20:@42669.4]
  wire  regs_360_reset; // @[RegFile.scala 66:20:@42669.4]
  wire [63:0] regs_360_io_in; // @[RegFile.scala 66:20:@42669.4]
  wire  regs_360_io_reset; // @[RegFile.scala 66:20:@42669.4]
  wire [63:0] regs_360_io_out; // @[RegFile.scala 66:20:@42669.4]
  wire  regs_360_io_enable; // @[RegFile.scala 66:20:@42669.4]
  wire  regs_361_clock; // @[RegFile.scala 66:20:@42683.4]
  wire  regs_361_reset; // @[RegFile.scala 66:20:@42683.4]
  wire [63:0] regs_361_io_in; // @[RegFile.scala 66:20:@42683.4]
  wire  regs_361_io_reset; // @[RegFile.scala 66:20:@42683.4]
  wire [63:0] regs_361_io_out; // @[RegFile.scala 66:20:@42683.4]
  wire  regs_361_io_enable; // @[RegFile.scala 66:20:@42683.4]
  wire  regs_362_clock; // @[RegFile.scala 66:20:@42697.4]
  wire  regs_362_reset; // @[RegFile.scala 66:20:@42697.4]
  wire [63:0] regs_362_io_in; // @[RegFile.scala 66:20:@42697.4]
  wire  regs_362_io_reset; // @[RegFile.scala 66:20:@42697.4]
  wire [63:0] regs_362_io_out; // @[RegFile.scala 66:20:@42697.4]
  wire  regs_362_io_enable; // @[RegFile.scala 66:20:@42697.4]
  wire  regs_363_clock; // @[RegFile.scala 66:20:@42711.4]
  wire  regs_363_reset; // @[RegFile.scala 66:20:@42711.4]
  wire [63:0] regs_363_io_in; // @[RegFile.scala 66:20:@42711.4]
  wire  regs_363_io_reset; // @[RegFile.scala 66:20:@42711.4]
  wire [63:0] regs_363_io_out; // @[RegFile.scala 66:20:@42711.4]
  wire  regs_363_io_enable; // @[RegFile.scala 66:20:@42711.4]
  wire  regs_364_clock; // @[RegFile.scala 66:20:@42725.4]
  wire  regs_364_reset; // @[RegFile.scala 66:20:@42725.4]
  wire [63:0] regs_364_io_in; // @[RegFile.scala 66:20:@42725.4]
  wire  regs_364_io_reset; // @[RegFile.scala 66:20:@42725.4]
  wire [63:0] regs_364_io_out; // @[RegFile.scala 66:20:@42725.4]
  wire  regs_364_io_enable; // @[RegFile.scala 66:20:@42725.4]
  wire  regs_365_clock; // @[RegFile.scala 66:20:@42739.4]
  wire  regs_365_reset; // @[RegFile.scala 66:20:@42739.4]
  wire [63:0] regs_365_io_in; // @[RegFile.scala 66:20:@42739.4]
  wire  regs_365_io_reset; // @[RegFile.scala 66:20:@42739.4]
  wire [63:0] regs_365_io_out; // @[RegFile.scala 66:20:@42739.4]
  wire  regs_365_io_enable; // @[RegFile.scala 66:20:@42739.4]
  wire  regs_366_clock; // @[RegFile.scala 66:20:@42753.4]
  wire  regs_366_reset; // @[RegFile.scala 66:20:@42753.4]
  wire [63:0] regs_366_io_in; // @[RegFile.scala 66:20:@42753.4]
  wire  regs_366_io_reset; // @[RegFile.scala 66:20:@42753.4]
  wire [63:0] regs_366_io_out; // @[RegFile.scala 66:20:@42753.4]
  wire  regs_366_io_enable; // @[RegFile.scala 66:20:@42753.4]
  wire  regs_367_clock; // @[RegFile.scala 66:20:@42767.4]
  wire  regs_367_reset; // @[RegFile.scala 66:20:@42767.4]
  wire [63:0] regs_367_io_in; // @[RegFile.scala 66:20:@42767.4]
  wire  regs_367_io_reset; // @[RegFile.scala 66:20:@42767.4]
  wire [63:0] regs_367_io_out; // @[RegFile.scala 66:20:@42767.4]
  wire  regs_367_io_enable; // @[RegFile.scala 66:20:@42767.4]
  wire  regs_368_clock; // @[RegFile.scala 66:20:@42781.4]
  wire  regs_368_reset; // @[RegFile.scala 66:20:@42781.4]
  wire [63:0] regs_368_io_in; // @[RegFile.scala 66:20:@42781.4]
  wire  regs_368_io_reset; // @[RegFile.scala 66:20:@42781.4]
  wire [63:0] regs_368_io_out; // @[RegFile.scala 66:20:@42781.4]
  wire  regs_368_io_enable; // @[RegFile.scala 66:20:@42781.4]
  wire  regs_369_clock; // @[RegFile.scala 66:20:@42795.4]
  wire  regs_369_reset; // @[RegFile.scala 66:20:@42795.4]
  wire [63:0] regs_369_io_in; // @[RegFile.scala 66:20:@42795.4]
  wire  regs_369_io_reset; // @[RegFile.scala 66:20:@42795.4]
  wire [63:0] regs_369_io_out; // @[RegFile.scala 66:20:@42795.4]
  wire  regs_369_io_enable; // @[RegFile.scala 66:20:@42795.4]
  wire  regs_370_clock; // @[RegFile.scala 66:20:@42809.4]
  wire  regs_370_reset; // @[RegFile.scala 66:20:@42809.4]
  wire [63:0] regs_370_io_in; // @[RegFile.scala 66:20:@42809.4]
  wire  regs_370_io_reset; // @[RegFile.scala 66:20:@42809.4]
  wire [63:0] regs_370_io_out; // @[RegFile.scala 66:20:@42809.4]
  wire  regs_370_io_enable; // @[RegFile.scala 66:20:@42809.4]
  wire  regs_371_clock; // @[RegFile.scala 66:20:@42823.4]
  wire  regs_371_reset; // @[RegFile.scala 66:20:@42823.4]
  wire [63:0] regs_371_io_in; // @[RegFile.scala 66:20:@42823.4]
  wire  regs_371_io_reset; // @[RegFile.scala 66:20:@42823.4]
  wire [63:0] regs_371_io_out; // @[RegFile.scala 66:20:@42823.4]
  wire  regs_371_io_enable; // @[RegFile.scala 66:20:@42823.4]
  wire  regs_372_clock; // @[RegFile.scala 66:20:@42837.4]
  wire  regs_372_reset; // @[RegFile.scala 66:20:@42837.4]
  wire [63:0] regs_372_io_in; // @[RegFile.scala 66:20:@42837.4]
  wire  regs_372_io_reset; // @[RegFile.scala 66:20:@42837.4]
  wire [63:0] regs_372_io_out; // @[RegFile.scala 66:20:@42837.4]
  wire  regs_372_io_enable; // @[RegFile.scala 66:20:@42837.4]
  wire  regs_373_clock; // @[RegFile.scala 66:20:@42851.4]
  wire  regs_373_reset; // @[RegFile.scala 66:20:@42851.4]
  wire [63:0] regs_373_io_in; // @[RegFile.scala 66:20:@42851.4]
  wire  regs_373_io_reset; // @[RegFile.scala 66:20:@42851.4]
  wire [63:0] regs_373_io_out; // @[RegFile.scala 66:20:@42851.4]
  wire  regs_373_io_enable; // @[RegFile.scala 66:20:@42851.4]
  wire  regs_374_clock; // @[RegFile.scala 66:20:@42865.4]
  wire  regs_374_reset; // @[RegFile.scala 66:20:@42865.4]
  wire [63:0] regs_374_io_in; // @[RegFile.scala 66:20:@42865.4]
  wire  regs_374_io_reset; // @[RegFile.scala 66:20:@42865.4]
  wire [63:0] regs_374_io_out; // @[RegFile.scala 66:20:@42865.4]
  wire  regs_374_io_enable; // @[RegFile.scala 66:20:@42865.4]
  wire  regs_375_clock; // @[RegFile.scala 66:20:@42879.4]
  wire  regs_375_reset; // @[RegFile.scala 66:20:@42879.4]
  wire [63:0] regs_375_io_in; // @[RegFile.scala 66:20:@42879.4]
  wire  regs_375_io_reset; // @[RegFile.scala 66:20:@42879.4]
  wire [63:0] regs_375_io_out; // @[RegFile.scala 66:20:@42879.4]
  wire  regs_375_io_enable; // @[RegFile.scala 66:20:@42879.4]
  wire  regs_376_clock; // @[RegFile.scala 66:20:@42893.4]
  wire  regs_376_reset; // @[RegFile.scala 66:20:@42893.4]
  wire [63:0] regs_376_io_in; // @[RegFile.scala 66:20:@42893.4]
  wire  regs_376_io_reset; // @[RegFile.scala 66:20:@42893.4]
  wire [63:0] regs_376_io_out; // @[RegFile.scala 66:20:@42893.4]
  wire  regs_376_io_enable; // @[RegFile.scala 66:20:@42893.4]
  wire  regs_377_clock; // @[RegFile.scala 66:20:@42907.4]
  wire  regs_377_reset; // @[RegFile.scala 66:20:@42907.4]
  wire [63:0] regs_377_io_in; // @[RegFile.scala 66:20:@42907.4]
  wire  regs_377_io_reset; // @[RegFile.scala 66:20:@42907.4]
  wire [63:0] regs_377_io_out; // @[RegFile.scala 66:20:@42907.4]
  wire  regs_377_io_enable; // @[RegFile.scala 66:20:@42907.4]
  wire  regs_378_clock; // @[RegFile.scala 66:20:@42921.4]
  wire  regs_378_reset; // @[RegFile.scala 66:20:@42921.4]
  wire [63:0] regs_378_io_in; // @[RegFile.scala 66:20:@42921.4]
  wire  regs_378_io_reset; // @[RegFile.scala 66:20:@42921.4]
  wire [63:0] regs_378_io_out; // @[RegFile.scala 66:20:@42921.4]
  wire  regs_378_io_enable; // @[RegFile.scala 66:20:@42921.4]
  wire  regs_379_clock; // @[RegFile.scala 66:20:@42935.4]
  wire  regs_379_reset; // @[RegFile.scala 66:20:@42935.4]
  wire [63:0] regs_379_io_in; // @[RegFile.scala 66:20:@42935.4]
  wire  regs_379_io_reset; // @[RegFile.scala 66:20:@42935.4]
  wire [63:0] regs_379_io_out; // @[RegFile.scala 66:20:@42935.4]
  wire  regs_379_io_enable; // @[RegFile.scala 66:20:@42935.4]
  wire  regs_380_clock; // @[RegFile.scala 66:20:@42949.4]
  wire  regs_380_reset; // @[RegFile.scala 66:20:@42949.4]
  wire [63:0] regs_380_io_in; // @[RegFile.scala 66:20:@42949.4]
  wire  regs_380_io_reset; // @[RegFile.scala 66:20:@42949.4]
  wire [63:0] regs_380_io_out; // @[RegFile.scala 66:20:@42949.4]
  wire  regs_380_io_enable; // @[RegFile.scala 66:20:@42949.4]
  wire  regs_381_clock; // @[RegFile.scala 66:20:@42963.4]
  wire  regs_381_reset; // @[RegFile.scala 66:20:@42963.4]
  wire [63:0] regs_381_io_in; // @[RegFile.scala 66:20:@42963.4]
  wire  regs_381_io_reset; // @[RegFile.scala 66:20:@42963.4]
  wire [63:0] regs_381_io_out; // @[RegFile.scala 66:20:@42963.4]
  wire  regs_381_io_enable; // @[RegFile.scala 66:20:@42963.4]
  wire  regs_382_clock; // @[RegFile.scala 66:20:@42977.4]
  wire  regs_382_reset; // @[RegFile.scala 66:20:@42977.4]
  wire [63:0] regs_382_io_in; // @[RegFile.scala 66:20:@42977.4]
  wire  regs_382_io_reset; // @[RegFile.scala 66:20:@42977.4]
  wire [63:0] regs_382_io_out; // @[RegFile.scala 66:20:@42977.4]
  wire  regs_382_io_enable; // @[RegFile.scala 66:20:@42977.4]
  wire  regs_383_clock; // @[RegFile.scala 66:20:@42991.4]
  wire  regs_383_reset; // @[RegFile.scala 66:20:@42991.4]
  wire [63:0] regs_383_io_in; // @[RegFile.scala 66:20:@42991.4]
  wire  regs_383_io_reset; // @[RegFile.scala 66:20:@42991.4]
  wire [63:0] regs_383_io_out; // @[RegFile.scala 66:20:@42991.4]
  wire  regs_383_io_enable; // @[RegFile.scala 66:20:@42991.4]
  wire  regs_384_clock; // @[RegFile.scala 66:20:@43005.4]
  wire  regs_384_reset; // @[RegFile.scala 66:20:@43005.4]
  wire [63:0] regs_384_io_in; // @[RegFile.scala 66:20:@43005.4]
  wire  regs_384_io_reset; // @[RegFile.scala 66:20:@43005.4]
  wire [63:0] regs_384_io_out; // @[RegFile.scala 66:20:@43005.4]
  wire  regs_384_io_enable; // @[RegFile.scala 66:20:@43005.4]
  wire  regs_385_clock; // @[RegFile.scala 66:20:@43019.4]
  wire  regs_385_reset; // @[RegFile.scala 66:20:@43019.4]
  wire [63:0] regs_385_io_in; // @[RegFile.scala 66:20:@43019.4]
  wire  regs_385_io_reset; // @[RegFile.scala 66:20:@43019.4]
  wire [63:0] regs_385_io_out; // @[RegFile.scala 66:20:@43019.4]
  wire  regs_385_io_enable; // @[RegFile.scala 66:20:@43019.4]
  wire  regs_386_clock; // @[RegFile.scala 66:20:@43033.4]
  wire  regs_386_reset; // @[RegFile.scala 66:20:@43033.4]
  wire [63:0] regs_386_io_in; // @[RegFile.scala 66:20:@43033.4]
  wire  regs_386_io_reset; // @[RegFile.scala 66:20:@43033.4]
  wire [63:0] regs_386_io_out; // @[RegFile.scala 66:20:@43033.4]
  wire  regs_386_io_enable; // @[RegFile.scala 66:20:@43033.4]
  wire  regs_387_clock; // @[RegFile.scala 66:20:@43047.4]
  wire  regs_387_reset; // @[RegFile.scala 66:20:@43047.4]
  wire [63:0] regs_387_io_in; // @[RegFile.scala 66:20:@43047.4]
  wire  regs_387_io_reset; // @[RegFile.scala 66:20:@43047.4]
  wire [63:0] regs_387_io_out; // @[RegFile.scala 66:20:@43047.4]
  wire  regs_387_io_enable; // @[RegFile.scala 66:20:@43047.4]
  wire  regs_388_clock; // @[RegFile.scala 66:20:@43061.4]
  wire  regs_388_reset; // @[RegFile.scala 66:20:@43061.4]
  wire [63:0] regs_388_io_in; // @[RegFile.scala 66:20:@43061.4]
  wire  regs_388_io_reset; // @[RegFile.scala 66:20:@43061.4]
  wire [63:0] regs_388_io_out; // @[RegFile.scala 66:20:@43061.4]
  wire  regs_388_io_enable; // @[RegFile.scala 66:20:@43061.4]
  wire  regs_389_clock; // @[RegFile.scala 66:20:@43075.4]
  wire  regs_389_reset; // @[RegFile.scala 66:20:@43075.4]
  wire [63:0] regs_389_io_in; // @[RegFile.scala 66:20:@43075.4]
  wire  regs_389_io_reset; // @[RegFile.scala 66:20:@43075.4]
  wire [63:0] regs_389_io_out; // @[RegFile.scala 66:20:@43075.4]
  wire  regs_389_io_enable; // @[RegFile.scala 66:20:@43075.4]
  wire  regs_390_clock; // @[RegFile.scala 66:20:@43089.4]
  wire  regs_390_reset; // @[RegFile.scala 66:20:@43089.4]
  wire [63:0] regs_390_io_in; // @[RegFile.scala 66:20:@43089.4]
  wire  regs_390_io_reset; // @[RegFile.scala 66:20:@43089.4]
  wire [63:0] regs_390_io_out; // @[RegFile.scala 66:20:@43089.4]
  wire  regs_390_io_enable; // @[RegFile.scala 66:20:@43089.4]
  wire  regs_391_clock; // @[RegFile.scala 66:20:@43103.4]
  wire  regs_391_reset; // @[RegFile.scala 66:20:@43103.4]
  wire [63:0] regs_391_io_in; // @[RegFile.scala 66:20:@43103.4]
  wire  regs_391_io_reset; // @[RegFile.scala 66:20:@43103.4]
  wire [63:0] regs_391_io_out; // @[RegFile.scala 66:20:@43103.4]
  wire  regs_391_io_enable; // @[RegFile.scala 66:20:@43103.4]
  wire  regs_392_clock; // @[RegFile.scala 66:20:@43117.4]
  wire  regs_392_reset; // @[RegFile.scala 66:20:@43117.4]
  wire [63:0] regs_392_io_in; // @[RegFile.scala 66:20:@43117.4]
  wire  regs_392_io_reset; // @[RegFile.scala 66:20:@43117.4]
  wire [63:0] regs_392_io_out; // @[RegFile.scala 66:20:@43117.4]
  wire  regs_392_io_enable; // @[RegFile.scala 66:20:@43117.4]
  wire  regs_393_clock; // @[RegFile.scala 66:20:@43131.4]
  wire  regs_393_reset; // @[RegFile.scala 66:20:@43131.4]
  wire [63:0] regs_393_io_in; // @[RegFile.scala 66:20:@43131.4]
  wire  regs_393_io_reset; // @[RegFile.scala 66:20:@43131.4]
  wire [63:0] regs_393_io_out; // @[RegFile.scala 66:20:@43131.4]
  wire  regs_393_io_enable; // @[RegFile.scala 66:20:@43131.4]
  wire  regs_394_clock; // @[RegFile.scala 66:20:@43145.4]
  wire  regs_394_reset; // @[RegFile.scala 66:20:@43145.4]
  wire [63:0] regs_394_io_in; // @[RegFile.scala 66:20:@43145.4]
  wire  regs_394_io_reset; // @[RegFile.scala 66:20:@43145.4]
  wire [63:0] regs_394_io_out; // @[RegFile.scala 66:20:@43145.4]
  wire  regs_394_io_enable; // @[RegFile.scala 66:20:@43145.4]
  wire  regs_395_clock; // @[RegFile.scala 66:20:@43159.4]
  wire  regs_395_reset; // @[RegFile.scala 66:20:@43159.4]
  wire [63:0] regs_395_io_in; // @[RegFile.scala 66:20:@43159.4]
  wire  regs_395_io_reset; // @[RegFile.scala 66:20:@43159.4]
  wire [63:0] regs_395_io_out; // @[RegFile.scala 66:20:@43159.4]
  wire  regs_395_io_enable; // @[RegFile.scala 66:20:@43159.4]
  wire  regs_396_clock; // @[RegFile.scala 66:20:@43173.4]
  wire  regs_396_reset; // @[RegFile.scala 66:20:@43173.4]
  wire [63:0] regs_396_io_in; // @[RegFile.scala 66:20:@43173.4]
  wire  regs_396_io_reset; // @[RegFile.scala 66:20:@43173.4]
  wire [63:0] regs_396_io_out; // @[RegFile.scala 66:20:@43173.4]
  wire  regs_396_io_enable; // @[RegFile.scala 66:20:@43173.4]
  wire  regs_397_clock; // @[RegFile.scala 66:20:@43187.4]
  wire  regs_397_reset; // @[RegFile.scala 66:20:@43187.4]
  wire [63:0] regs_397_io_in; // @[RegFile.scala 66:20:@43187.4]
  wire  regs_397_io_reset; // @[RegFile.scala 66:20:@43187.4]
  wire [63:0] regs_397_io_out; // @[RegFile.scala 66:20:@43187.4]
  wire  regs_397_io_enable; // @[RegFile.scala 66:20:@43187.4]
  wire  regs_398_clock; // @[RegFile.scala 66:20:@43201.4]
  wire  regs_398_reset; // @[RegFile.scala 66:20:@43201.4]
  wire [63:0] regs_398_io_in; // @[RegFile.scala 66:20:@43201.4]
  wire  regs_398_io_reset; // @[RegFile.scala 66:20:@43201.4]
  wire [63:0] regs_398_io_out; // @[RegFile.scala 66:20:@43201.4]
  wire  regs_398_io_enable; // @[RegFile.scala 66:20:@43201.4]
  wire  regs_399_clock; // @[RegFile.scala 66:20:@43215.4]
  wire  regs_399_reset; // @[RegFile.scala 66:20:@43215.4]
  wire [63:0] regs_399_io_in; // @[RegFile.scala 66:20:@43215.4]
  wire  regs_399_io_reset; // @[RegFile.scala 66:20:@43215.4]
  wire [63:0] regs_399_io_out; // @[RegFile.scala 66:20:@43215.4]
  wire  regs_399_io_enable; // @[RegFile.scala 66:20:@43215.4]
  wire  regs_400_clock; // @[RegFile.scala 66:20:@43229.4]
  wire  regs_400_reset; // @[RegFile.scala 66:20:@43229.4]
  wire [63:0] regs_400_io_in; // @[RegFile.scala 66:20:@43229.4]
  wire  regs_400_io_reset; // @[RegFile.scala 66:20:@43229.4]
  wire [63:0] regs_400_io_out; // @[RegFile.scala 66:20:@43229.4]
  wire  regs_400_io_enable; // @[RegFile.scala 66:20:@43229.4]
  wire  regs_401_clock; // @[RegFile.scala 66:20:@43243.4]
  wire  regs_401_reset; // @[RegFile.scala 66:20:@43243.4]
  wire [63:0] regs_401_io_in; // @[RegFile.scala 66:20:@43243.4]
  wire  regs_401_io_reset; // @[RegFile.scala 66:20:@43243.4]
  wire [63:0] regs_401_io_out; // @[RegFile.scala 66:20:@43243.4]
  wire  regs_401_io_enable; // @[RegFile.scala 66:20:@43243.4]
  wire  regs_402_clock; // @[RegFile.scala 66:20:@43257.4]
  wire  regs_402_reset; // @[RegFile.scala 66:20:@43257.4]
  wire [63:0] regs_402_io_in; // @[RegFile.scala 66:20:@43257.4]
  wire  regs_402_io_reset; // @[RegFile.scala 66:20:@43257.4]
  wire [63:0] regs_402_io_out; // @[RegFile.scala 66:20:@43257.4]
  wire  regs_402_io_enable; // @[RegFile.scala 66:20:@43257.4]
  wire  regs_403_clock; // @[RegFile.scala 66:20:@43271.4]
  wire  regs_403_reset; // @[RegFile.scala 66:20:@43271.4]
  wire [63:0] regs_403_io_in; // @[RegFile.scala 66:20:@43271.4]
  wire  regs_403_io_reset; // @[RegFile.scala 66:20:@43271.4]
  wire [63:0] regs_403_io_out; // @[RegFile.scala 66:20:@43271.4]
  wire  regs_403_io_enable; // @[RegFile.scala 66:20:@43271.4]
  wire  regs_404_clock; // @[RegFile.scala 66:20:@43285.4]
  wire  regs_404_reset; // @[RegFile.scala 66:20:@43285.4]
  wire [63:0] regs_404_io_in; // @[RegFile.scala 66:20:@43285.4]
  wire  regs_404_io_reset; // @[RegFile.scala 66:20:@43285.4]
  wire [63:0] regs_404_io_out; // @[RegFile.scala 66:20:@43285.4]
  wire  regs_404_io_enable; // @[RegFile.scala 66:20:@43285.4]
  wire  regs_405_clock; // @[RegFile.scala 66:20:@43299.4]
  wire  regs_405_reset; // @[RegFile.scala 66:20:@43299.4]
  wire [63:0] regs_405_io_in; // @[RegFile.scala 66:20:@43299.4]
  wire  regs_405_io_reset; // @[RegFile.scala 66:20:@43299.4]
  wire [63:0] regs_405_io_out; // @[RegFile.scala 66:20:@43299.4]
  wire  regs_405_io_enable; // @[RegFile.scala 66:20:@43299.4]
  wire  regs_406_clock; // @[RegFile.scala 66:20:@43313.4]
  wire  regs_406_reset; // @[RegFile.scala 66:20:@43313.4]
  wire [63:0] regs_406_io_in; // @[RegFile.scala 66:20:@43313.4]
  wire  regs_406_io_reset; // @[RegFile.scala 66:20:@43313.4]
  wire [63:0] regs_406_io_out; // @[RegFile.scala 66:20:@43313.4]
  wire  regs_406_io_enable; // @[RegFile.scala 66:20:@43313.4]
  wire  regs_407_clock; // @[RegFile.scala 66:20:@43327.4]
  wire  regs_407_reset; // @[RegFile.scala 66:20:@43327.4]
  wire [63:0] regs_407_io_in; // @[RegFile.scala 66:20:@43327.4]
  wire  regs_407_io_reset; // @[RegFile.scala 66:20:@43327.4]
  wire [63:0] regs_407_io_out; // @[RegFile.scala 66:20:@43327.4]
  wire  regs_407_io_enable; // @[RegFile.scala 66:20:@43327.4]
  wire  regs_408_clock; // @[RegFile.scala 66:20:@43341.4]
  wire  regs_408_reset; // @[RegFile.scala 66:20:@43341.4]
  wire [63:0] regs_408_io_in; // @[RegFile.scala 66:20:@43341.4]
  wire  regs_408_io_reset; // @[RegFile.scala 66:20:@43341.4]
  wire [63:0] regs_408_io_out; // @[RegFile.scala 66:20:@43341.4]
  wire  regs_408_io_enable; // @[RegFile.scala 66:20:@43341.4]
  wire  regs_409_clock; // @[RegFile.scala 66:20:@43355.4]
  wire  regs_409_reset; // @[RegFile.scala 66:20:@43355.4]
  wire [63:0] regs_409_io_in; // @[RegFile.scala 66:20:@43355.4]
  wire  regs_409_io_reset; // @[RegFile.scala 66:20:@43355.4]
  wire [63:0] regs_409_io_out; // @[RegFile.scala 66:20:@43355.4]
  wire  regs_409_io_enable; // @[RegFile.scala 66:20:@43355.4]
  wire  regs_410_clock; // @[RegFile.scala 66:20:@43369.4]
  wire  regs_410_reset; // @[RegFile.scala 66:20:@43369.4]
  wire [63:0] regs_410_io_in; // @[RegFile.scala 66:20:@43369.4]
  wire  regs_410_io_reset; // @[RegFile.scala 66:20:@43369.4]
  wire [63:0] regs_410_io_out; // @[RegFile.scala 66:20:@43369.4]
  wire  regs_410_io_enable; // @[RegFile.scala 66:20:@43369.4]
  wire  regs_411_clock; // @[RegFile.scala 66:20:@43383.4]
  wire  regs_411_reset; // @[RegFile.scala 66:20:@43383.4]
  wire [63:0] regs_411_io_in; // @[RegFile.scala 66:20:@43383.4]
  wire  regs_411_io_reset; // @[RegFile.scala 66:20:@43383.4]
  wire [63:0] regs_411_io_out; // @[RegFile.scala 66:20:@43383.4]
  wire  regs_411_io_enable; // @[RegFile.scala 66:20:@43383.4]
  wire  regs_412_clock; // @[RegFile.scala 66:20:@43397.4]
  wire  regs_412_reset; // @[RegFile.scala 66:20:@43397.4]
  wire [63:0] regs_412_io_in; // @[RegFile.scala 66:20:@43397.4]
  wire  regs_412_io_reset; // @[RegFile.scala 66:20:@43397.4]
  wire [63:0] regs_412_io_out; // @[RegFile.scala 66:20:@43397.4]
  wire  regs_412_io_enable; // @[RegFile.scala 66:20:@43397.4]
  wire  regs_413_clock; // @[RegFile.scala 66:20:@43411.4]
  wire  regs_413_reset; // @[RegFile.scala 66:20:@43411.4]
  wire [63:0] regs_413_io_in; // @[RegFile.scala 66:20:@43411.4]
  wire  regs_413_io_reset; // @[RegFile.scala 66:20:@43411.4]
  wire [63:0] regs_413_io_out; // @[RegFile.scala 66:20:@43411.4]
  wire  regs_413_io_enable; // @[RegFile.scala 66:20:@43411.4]
  wire  regs_414_clock; // @[RegFile.scala 66:20:@43425.4]
  wire  regs_414_reset; // @[RegFile.scala 66:20:@43425.4]
  wire [63:0] regs_414_io_in; // @[RegFile.scala 66:20:@43425.4]
  wire  regs_414_io_reset; // @[RegFile.scala 66:20:@43425.4]
  wire [63:0] regs_414_io_out; // @[RegFile.scala 66:20:@43425.4]
  wire  regs_414_io_enable; // @[RegFile.scala 66:20:@43425.4]
  wire  regs_415_clock; // @[RegFile.scala 66:20:@43439.4]
  wire  regs_415_reset; // @[RegFile.scala 66:20:@43439.4]
  wire [63:0] regs_415_io_in; // @[RegFile.scala 66:20:@43439.4]
  wire  regs_415_io_reset; // @[RegFile.scala 66:20:@43439.4]
  wire [63:0] regs_415_io_out; // @[RegFile.scala 66:20:@43439.4]
  wire  regs_415_io_enable; // @[RegFile.scala 66:20:@43439.4]
  wire  regs_416_clock; // @[RegFile.scala 66:20:@43453.4]
  wire  regs_416_reset; // @[RegFile.scala 66:20:@43453.4]
  wire [63:0] regs_416_io_in; // @[RegFile.scala 66:20:@43453.4]
  wire  regs_416_io_reset; // @[RegFile.scala 66:20:@43453.4]
  wire [63:0] regs_416_io_out; // @[RegFile.scala 66:20:@43453.4]
  wire  regs_416_io_enable; // @[RegFile.scala 66:20:@43453.4]
  wire  regs_417_clock; // @[RegFile.scala 66:20:@43467.4]
  wire  regs_417_reset; // @[RegFile.scala 66:20:@43467.4]
  wire [63:0] regs_417_io_in; // @[RegFile.scala 66:20:@43467.4]
  wire  regs_417_io_reset; // @[RegFile.scala 66:20:@43467.4]
  wire [63:0] regs_417_io_out; // @[RegFile.scala 66:20:@43467.4]
  wire  regs_417_io_enable; // @[RegFile.scala 66:20:@43467.4]
  wire  regs_418_clock; // @[RegFile.scala 66:20:@43481.4]
  wire  regs_418_reset; // @[RegFile.scala 66:20:@43481.4]
  wire [63:0] regs_418_io_in; // @[RegFile.scala 66:20:@43481.4]
  wire  regs_418_io_reset; // @[RegFile.scala 66:20:@43481.4]
  wire [63:0] regs_418_io_out; // @[RegFile.scala 66:20:@43481.4]
  wire  regs_418_io_enable; // @[RegFile.scala 66:20:@43481.4]
  wire  regs_419_clock; // @[RegFile.scala 66:20:@43495.4]
  wire  regs_419_reset; // @[RegFile.scala 66:20:@43495.4]
  wire [63:0] regs_419_io_in; // @[RegFile.scala 66:20:@43495.4]
  wire  regs_419_io_reset; // @[RegFile.scala 66:20:@43495.4]
  wire [63:0] regs_419_io_out; // @[RegFile.scala 66:20:@43495.4]
  wire  regs_419_io_enable; // @[RegFile.scala 66:20:@43495.4]
  wire  regs_420_clock; // @[RegFile.scala 66:20:@43509.4]
  wire  regs_420_reset; // @[RegFile.scala 66:20:@43509.4]
  wire [63:0] regs_420_io_in; // @[RegFile.scala 66:20:@43509.4]
  wire  regs_420_io_reset; // @[RegFile.scala 66:20:@43509.4]
  wire [63:0] regs_420_io_out; // @[RegFile.scala 66:20:@43509.4]
  wire  regs_420_io_enable; // @[RegFile.scala 66:20:@43509.4]
  wire  regs_421_clock; // @[RegFile.scala 66:20:@43523.4]
  wire  regs_421_reset; // @[RegFile.scala 66:20:@43523.4]
  wire [63:0] regs_421_io_in; // @[RegFile.scala 66:20:@43523.4]
  wire  regs_421_io_reset; // @[RegFile.scala 66:20:@43523.4]
  wire [63:0] regs_421_io_out; // @[RegFile.scala 66:20:@43523.4]
  wire  regs_421_io_enable; // @[RegFile.scala 66:20:@43523.4]
  wire  regs_422_clock; // @[RegFile.scala 66:20:@43537.4]
  wire  regs_422_reset; // @[RegFile.scala 66:20:@43537.4]
  wire [63:0] regs_422_io_in; // @[RegFile.scala 66:20:@43537.4]
  wire  regs_422_io_reset; // @[RegFile.scala 66:20:@43537.4]
  wire [63:0] regs_422_io_out; // @[RegFile.scala 66:20:@43537.4]
  wire  regs_422_io_enable; // @[RegFile.scala 66:20:@43537.4]
  wire  regs_423_clock; // @[RegFile.scala 66:20:@43551.4]
  wire  regs_423_reset; // @[RegFile.scala 66:20:@43551.4]
  wire [63:0] regs_423_io_in; // @[RegFile.scala 66:20:@43551.4]
  wire  regs_423_io_reset; // @[RegFile.scala 66:20:@43551.4]
  wire [63:0] regs_423_io_out; // @[RegFile.scala 66:20:@43551.4]
  wire  regs_423_io_enable; // @[RegFile.scala 66:20:@43551.4]
  wire  regs_424_clock; // @[RegFile.scala 66:20:@43565.4]
  wire  regs_424_reset; // @[RegFile.scala 66:20:@43565.4]
  wire [63:0] regs_424_io_in; // @[RegFile.scala 66:20:@43565.4]
  wire  regs_424_io_reset; // @[RegFile.scala 66:20:@43565.4]
  wire [63:0] regs_424_io_out; // @[RegFile.scala 66:20:@43565.4]
  wire  regs_424_io_enable; // @[RegFile.scala 66:20:@43565.4]
  wire  regs_425_clock; // @[RegFile.scala 66:20:@43579.4]
  wire  regs_425_reset; // @[RegFile.scala 66:20:@43579.4]
  wire [63:0] regs_425_io_in; // @[RegFile.scala 66:20:@43579.4]
  wire  regs_425_io_reset; // @[RegFile.scala 66:20:@43579.4]
  wire [63:0] regs_425_io_out; // @[RegFile.scala 66:20:@43579.4]
  wire  regs_425_io_enable; // @[RegFile.scala 66:20:@43579.4]
  wire  regs_426_clock; // @[RegFile.scala 66:20:@43593.4]
  wire  regs_426_reset; // @[RegFile.scala 66:20:@43593.4]
  wire [63:0] regs_426_io_in; // @[RegFile.scala 66:20:@43593.4]
  wire  regs_426_io_reset; // @[RegFile.scala 66:20:@43593.4]
  wire [63:0] regs_426_io_out; // @[RegFile.scala 66:20:@43593.4]
  wire  regs_426_io_enable; // @[RegFile.scala 66:20:@43593.4]
  wire  regs_427_clock; // @[RegFile.scala 66:20:@43607.4]
  wire  regs_427_reset; // @[RegFile.scala 66:20:@43607.4]
  wire [63:0] regs_427_io_in; // @[RegFile.scala 66:20:@43607.4]
  wire  regs_427_io_reset; // @[RegFile.scala 66:20:@43607.4]
  wire [63:0] regs_427_io_out; // @[RegFile.scala 66:20:@43607.4]
  wire  regs_427_io_enable; // @[RegFile.scala 66:20:@43607.4]
  wire  regs_428_clock; // @[RegFile.scala 66:20:@43621.4]
  wire  regs_428_reset; // @[RegFile.scala 66:20:@43621.4]
  wire [63:0] regs_428_io_in; // @[RegFile.scala 66:20:@43621.4]
  wire  regs_428_io_reset; // @[RegFile.scala 66:20:@43621.4]
  wire [63:0] regs_428_io_out; // @[RegFile.scala 66:20:@43621.4]
  wire  regs_428_io_enable; // @[RegFile.scala 66:20:@43621.4]
  wire  regs_429_clock; // @[RegFile.scala 66:20:@43635.4]
  wire  regs_429_reset; // @[RegFile.scala 66:20:@43635.4]
  wire [63:0] regs_429_io_in; // @[RegFile.scala 66:20:@43635.4]
  wire  regs_429_io_reset; // @[RegFile.scala 66:20:@43635.4]
  wire [63:0] regs_429_io_out; // @[RegFile.scala 66:20:@43635.4]
  wire  regs_429_io_enable; // @[RegFile.scala 66:20:@43635.4]
  wire  regs_430_clock; // @[RegFile.scala 66:20:@43649.4]
  wire  regs_430_reset; // @[RegFile.scala 66:20:@43649.4]
  wire [63:0] regs_430_io_in; // @[RegFile.scala 66:20:@43649.4]
  wire  regs_430_io_reset; // @[RegFile.scala 66:20:@43649.4]
  wire [63:0] regs_430_io_out; // @[RegFile.scala 66:20:@43649.4]
  wire  regs_430_io_enable; // @[RegFile.scala 66:20:@43649.4]
  wire  regs_431_clock; // @[RegFile.scala 66:20:@43663.4]
  wire  regs_431_reset; // @[RegFile.scala 66:20:@43663.4]
  wire [63:0] regs_431_io_in; // @[RegFile.scala 66:20:@43663.4]
  wire  regs_431_io_reset; // @[RegFile.scala 66:20:@43663.4]
  wire [63:0] regs_431_io_out; // @[RegFile.scala 66:20:@43663.4]
  wire  regs_431_io_enable; // @[RegFile.scala 66:20:@43663.4]
  wire  regs_432_clock; // @[RegFile.scala 66:20:@43677.4]
  wire  regs_432_reset; // @[RegFile.scala 66:20:@43677.4]
  wire [63:0] regs_432_io_in; // @[RegFile.scala 66:20:@43677.4]
  wire  regs_432_io_reset; // @[RegFile.scala 66:20:@43677.4]
  wire [63:0] regs_432_io_out; // @[RegFile.scala 66:20:@43677.4]
  wire  regs_432_io_enable; // @[RegFile.scala 66:20:@43677.4]
  wire  regs_433_clock; // @[RegFile.scala 66:20:@43691.4]
  wire  regs_433_reset; // @[RegFile.scala 66:20:@43691.4]
  wire [63:0] regs_433_io_in; // @[RegFile.scala 66:20:@43691.4]
  wire  regs_433_io_reset; // @[RegFile.scala 66:20:@43691.4]
  wire [63:0] regs_433_io_out; // @[RegFile.scala 66:20:@43691.4]
  wire  regs_433_io_enable; // @[RegFile.scala 66:20:@43691.4]
  wire  regs_434_clock; // @[RegFile.scala 66:20:@43705.4]
  wire  regs_434_reset; // @[RegFile.scala 66:20:@43705.4]
  wire [63:0] regs_434_io_in; // @[RegFile.scala 66:20:@43705.4]
  wire  regs_434_io_reset; // @[RegFile.scala 66:20:@43705.4]
  wire [63:0] regs_434_io_out; // @[RegFile.scala 66:20:@43705.4]
  wire  regs_434_io_enable; // @[RegFile.scala 66:20:@43705.4]
  wire  regs_435_clock; // @[RegFile.scala 66:20:@43719.4]
  wire  regs_435_reset; // @[RegFile.scala 66:20:@43719.4]
  wire [63:0] regs_435_io_in; // @[RegFile.scala 66:20:@43719.4]
  wire  regs_435_io_reset; // @[RegFile.scala 66:20:@43719.4]
  wire [63:0] regs_435_io_out; // @[RegFile.scala 66:20:@43719.4]
  wire  regs_435_io_enable; // @[RegFile.scala 66:20:@43719.4]
  wire  regs_436_clock; // @[RegFile.scala 66:20:@43733.4]
  wire  regs_436_reset; // @[RegFile.scala 66:20:@43733.4]
  wire [63:0] regs_436_io_in; // @[RegFile.scala 66:20:@43733.4]
  wire  regs_436_io_reset; // @[RegFile.scala 66:20:@43733.4]
  wire [63:0] regs_436_io_out; // @[RegFile.scala 66:20:@43733.4]
  wire  regs_436_io_enable; // @[RegFile.scala 66:20:@43733.4]
  wire  regs_437_clock; // @[RegFile.scala 66:20:@43747.4]
  wire  regs_437_reset; // @[RegFile.scala 66:20:@43747.4]
  wire [63:0] regs_437_io_in; // @[RegFile.scala 66:20:@43747.4]
  wire  regs_437_io_reset; // @[RegFile.scala 66:20:@43747.4]
  wire [63:0] regs_437_io_out; // @[RegFile.scala 66:20:@43747.4]
  wire  regs_437_io_enable; // @[RegFile.scala 66:20:@43747.4]
  wire  regs_438_clock; // @[RegFile.scala 66:20:@43761.4]
  wire  regs_438_reset; // @[RegFile.scala 66:20:@43761.4]
  wire [63:0] regs_438_io_in; // @[RegFile.scala 66:20:@43761.4]
  wire  regs_438_io_reset; // @[RegFile.scala 66:20:@43761.4]
  wire [63:0] regs_438_io_out; // @[RegFile.scala 66:20:@43761.4]
  wire  regs_438_io_enable; // @[RegFile.scala 66:20:@43761.4]
  wire  regs_439_clock; // @[RegFile.scala 66:20:@43775.4]
  wire  regs_439_reset; // @[RegFile.scala 66:20:@43775.4]
  wire [63:0] regs_439_io_in; // @[RegFile.scala 66:20:@43775.4]
  wire  regs_439_io_reset; // @[RegFile.scala 66:20:@43775.4]
  wire [63:0] regs_439_io_out; // @[RegFile.scala 66:20:@43775.4]
  wire  regs_439_io_enable; // @[RegFile.scala 66:20:@43775.4]
  wire  regs_440_clock; // @[RegFile.scala 66:20:@43789.4]
  wire  regs_440_reset; // @[RegFile.scala 66:20:@43789.4]
  wire [63:0] regs_440_io_in; // @[RegFile.scala 66:20:@43789.4]
  wire  regs_440_io_reset; // @[RegFile.scala 66:20:@43789.4]
  wire [63:0] regs_440_io_out; // @[RegFile.scala 66:20:@43789.4]
  wire  regs_440_io_enable; // @[RegFile.scala 66:20:@43789.4]
  wire  regs_441_clock; // @[RegFile.scala 66:20:@43803.4]
  wire  regs_441_reset; // @[RegFile.scala 66:20:@43803.4]
  wire [63:0] regs_441_io_in; // @[RegFile.scala 66:20:@43803.4]
  wire  regs_441_io_reset; // @[RegFile.scala 66:20:@43803.4]
  wire [63:0] regs_441_io_out; // @[RegFile.scala 66:20:@43803.4]
  wire  regs_441_io_enable; // @[RegFile.scala 66:20:@43803.4]
  wire  regs_442_clock; // @[RegFile.scala 66:20:@43817.4]
  wire  regs_442_reset; // @[RegFile.scala 66:20:@43817.4]
  wire [63:0] regs_442_io_in; // @[RegFile.scala 66:20:@43817.4]
  wire  regs_442_io_reset; // @[RegFile.scala 66:20:@43817.4]
  wire [63:0] regs_442_io_out; // @[RegFile.scala 66:20:@43817.4]
  wire  regs_442_io_enable; // @[RegFile.scala 66:20:@43817.4]
  wire  regs_443_clock; // @[RegFile.scala 66:20:@43831.4]
  wire  regs_443_reset; // @[RegFile.scala 66:20:@43831.4]
  wire [63:0] regs_443_io_in; // @[RegFile.scala 66:20:@43831.4]
  wire  regs_443_io_reset; // @[RegFile.scala 66:20:@43831.4]
  wire [63:0] regs_443_io_out; // @[RegFile.scala 66:20:@43831.4]
  wire  regs_443_io_enable; // @[RegFile.scala 66:20:@43831.4]
  wire  regs_444_clock; // @[RegFile.scala 66:20:@43845.4]
  wire  regs_444_reset; // @[RegFile.scala 66:20:@43845.4]
  wire [63:0] regs_444_io_in; // @[RegFile.scala 66:20:@43845.4]
  wire  regs_444_io_reset; // @[RegFile.scala 66:20:@43845.4]
  wire [63:0] regs_444_io_out; // @[RegFile.scala 66:20:@43845.4]
  wire  regs_444_io_enable; // @[RegFile.scala 66:20:@43845.4]
  wire  regs_445_clock; // @[RegFile.scala 66:20:@43859.4]
  wire  regs_445_reset; // @[RegFile.scala 66:20:@43859.4]
  wire [63:0] regs_445_io_in; // @[RegFile.scala 66:20:@43859.4]
  wire  regs_445_io_reset; // @[RegFile.scala 66:20:@43859.4]
  wire [63:0] regs_445_io_out; // @[RegFile.scala 66:20:@43859.4]
  wire  regs_445_io_enable; // @[RegFile.scala 66:20:@43859.4]
  wire  regs_446_clock; // @[RegFile.scala 66:20:@43873.4]
  wire  regs_446_reset; // @[RegFile.scala 66:20:@43873.4]
  wire [63:0] regs_446_io_in; // @[RegFile.scala 66:20:@43873.4]
  wire  regs_446_io_reset; // @[RegFile.scala 66:20:@43873.4]
  wire [63:0] regs_446_io_out; // @[RegFile.scala 66:20:@43873.4]
  wire  regs_446_io_enable; // @[RegFile.scala 66:20:@43873.4]
  wire  regs_447_clock; // @[RegFile.scala 66:20:@43887.4]
  wire  regs_447_reset; // @[RegFile.scala 66:20:@43887.4]
  wire [63:0] regs_447_io_in; // @[RegFile.scala 66:20:@43887.4]
  wire  regs_447_io_reset; // @[RegFile.scala 66:20:@43887.4]
  wire [63:0] regs_447_io_out; // @[RegFile.scala 66:20:@43887.4]
  wire  regs_447_io_enable; // @[RegFile.scala 66:20:@43887.4]
  wire  regs_448_clock; // @[RegFile.scala 66:20:@43901.4]
  wire  regs_448_reset; // @[RegFile.scala 66:20:@43901.4]
  wire [63:0] regs_448_io_in; // @[RegFile.scala 66:20:@43901.4]
  wire  regs_448_io_reset; // @[RegFile.scala 66:20:@43901.4]
  wire [63:0] regs_448_io_out; // @[RegFile.scala 66:20:@43901.4]
  wire  regs_448_io_enable; // @[RegFile.scala 66:20:@43901.4]
  wire  regs_449_clock; // @[RegFile.scala 66:20:@43915.4]
  wire  regs_449_reset; // @[RegFile.scala 66:20:@43915.4]
  wire [63:0] regs_449_io_in; // @[RegFile.scala 66:20:@43915.4]
  wire  regs_449_io_reset; // @[RegFile.scala 66:20:@43915.4]
  wire [63:0] regs_449_io_out; // @[RegFile.scala 66:20:@43915.4]
  wire  regs_449_io_enable; // @[RegFile.scala 66:20:@43915.4]
  wire  regs_450_clock; // @[RegFile.scala 66:20:@43929.4]
  wire  regs_450_reset; // @[RegFile.scala 66:20:@43929.4]
  wire [63:0] regs_450_io_in; // @[RegFile.scala 66:20:@43929.4]
  wire  regs_450_io_reset; // @[RegFile.scala 66:20:@43929.4]
  wire [63:0] regs_450_io_out; // @[RegFile.scala 66:20:@43929.4]
  wire  regs_450_io_enable; // @[RegFile.scala 66:20:@43929.4]
  wire  regs_451_clock; // @[RegFile.scala 66:20:@43943.4]
  wire  regs_451_reset; // @[RegFile.scala 66:20:@43943.4]
  wire [63:0] regs_451_io_in; // @[RegFile.scala 66:20:@43943.4]
  wire  regs_451_io_reset; // @[RegFile.scala 66:20:@43943.4]
  wire [63:0] regs_451_io_out; // @[RegFile.scala 66:20:@43943.4]
  wire  regs_451_io_enable; // @[RegFile.scala 66:20:@43943.4]
  wire  regs_452_clock; // @[RegFile.scala 66:20:@43957.4]
  wire  regs_452_reset; // @[RegFile.scala 66:20:@43957.4]
  wire [63:0] regs_452_io_in; // @[RegFile.scala 66:20:@43957.4]
  wire  regs_452_io_reset; // @[RegFile.scala 66:20:@43957.4]
  wire [63:0] regs_452_io_out; // @[RegFile.scala 66:20:@43957.4]
  wire  regs_452_io_enable; // @[RegFile.scala 66:20:@43957.4]
  wire  regs_453_clock; // @[RegFile.scala 66:20:@43971.4]
  wire  regs_453_reset; // @[RegFile.scala 66:20:@43971.4]
  wire [63:0] regs_453_io_in; // @[RegFile.scala 66:20:@43971.4]
  wire  regs_453_io_reset; // @[RegFile.scala 66:20:@43971.4]
  wire [63:0] regs_453_io_out; // @[RegFile.scala 66:20:@43971.4]
  wire  regs_453_io_enable; // @[RegFile.scala 66:20:@43971.4]
  wire  regs_454_clock; // @[RegFile.scala 66:20:@43985.4]
  wire  regs_454_reset; // @[RegFile.scala 66:20:@43985.4]
  wire [63:0] regs_454_io_in; // @[RegFile.scala 66:20:@43985.4]
  wire  regs_454_io_reset; // @[RegFile.scala 66:20:@43985.4]
  wire [63:0] regs_454_io_out; // @[RegFile.scala 66:20:@43985.4]
  wire  regs_454_io_enable; // @[RegFile.scala 66:20:@43985.4]
  wire  regs_455_clock; // @[RegFile.scala 66:20:@43999.4]
  wire  regs_455_reset; // @[RegFile.scala 66:20:@43999.4]
  wire [63:0] regs_455_io_in; // @[RegFile.scala 66:20:@43999.4]
  wire  regs_455_io_reset; // @[RegFile.scala 66:20:@43999.4]
  wire [63:0] regs_455_io_out; // @[RegFile.scala 66:20:@43999.4]
  wire  regs_455_io_enable; // @[RegFile.scala 66:20:@43999.4]
  wire  regs_456_clock; // @[RegFile.scala 66:20:@44013.4]
  wire  regs_456_reset; // @[RegFile.scala 66:20:@44013.4]
  wire [63:0] regs_456_io_in; // @[RegFile.scala 66:20:@44013.4]
  wire  regs_456_io_reset; // @[RegFile.scala 66:20:@44013.4]
  wire [63:0] regs_456_io_out; // @[RegFile.scala 66:20:@44013.4]
  wire  regs_456_io_enable; // @[RegFile.scala 66:20:@44013.4]
  wire  regs_457_clock; // @[RegFile.scala 66:20:@44027.4]
  wire  regs_457_reset; // @[RegFile.scala 66:20:@44027.4]
  wire [63:0] regs_457_io_in; // @[RegFile.scala 66:20:@44027.4]
  wire  regs_457_io_reset; // @[RegFile.scala 66:20:@44027.4]
  wire [63:0] regs_457_io_out; // @[RegFile.scala 66:20:@44027.4]
  wire  regs_457_io_enable; // @[RegFile.scala 66:20:@44027.4]
  wire  regs_458_clock; // @[RegFile.scala 66:20:@44041.4]
  wire  regs_458_reset; // @[RegFile.scala 66:20:@44041.4]
  wire [63:0] regs_458_io_in; // @[RegFile.scala 66:20:@44041.4]
  wire  regs_458_io_reset; // @[RegFile.scala 66:20:@44041.4]
  wire [63:0] regs_458_io_out; // @[RegFile.scala 66:20:@44041.4]
  wire  regs_458_io_enable; // @[RegFile.scala 66:20:@44041.4]
  wire  regs_459_clock; // @[RegFile.scala 66:20:@44055.4]
  wire  regs_459_reset; // @[RegFile.scala 66:20:@44055.4]
  wire [63:0] regs_459_io_in; // @[RegFile.scala 66:20:@44055.4]
  wire  regs_459_io_reset; // @[RegFile.scala 66:20:@44055.4]
  wire [63:0] regs_459_io_out; // @[RegFile.scala 66:20:@44055.4]
  wire  regs_459_io_enable; // @[RegFile.scala 66:20:@44055.4]
  wire  regs_460_clock; // @[RegFile.scala 66:20:@44069.4]
  wire  regs_460_reset; // @[RegFile.scala 66:20:@44069.4]
  wire [63:0] regs_460_io_in; // @[RegFile.scala 66:20:@44069.4]
  wire  regs_460_io_reset; // @[RegFile.scala 66:20:@44069.4]
  wire [63:0] regs_460_io_out; // @[RegFile.scala 66:20:@44069.4]
  wire  regs_460_io_enable; // @[RegFile.scala 66:20:@44069.4]
  wire  regs_461_clock; // @[RegFile.scala 66:20:@44083.4]
  wire  regs_461_reset; // @[RegFile.scala 66:20:@44083.4]
  wire [63:0] regs_461_io_in; // @[RegFile.scala 66:20:@44083.4]
  wire  regs_461_io_reset; // @[RegFile.scala 66:20:@44083.4]
  wire [63:0] regs_461_io_out; // @[RegFile.scala 66:20:@44083.4]
  wire  regs_461_io_enable; // @[RegFile.scala 66:20:@44083.4]
  wire  regs_462_clock; // @[RegFile.scala 66:20:@44097.4]
  wire  regs_462_reset; // @[RegFile.scala 66:20:@44097.4]
  wire [63:0] regs_462_io_in; // @[RegFile.scala 66:20:@44097.4]
  wire  regs_462_io_reset; // @[RegFile.scala 66:20:@44097.4]
  wire [63:0] regs_462_io_out; // @[RegFile.scala 66:20:@44097.4]
  wire  regs_462_io_enable; // @[RegFile.scala 66:20:@44097.4]
  wire  regs_463_clock; // @[RegFile.scala 66:20:@44111.4]
  wire  regs_463_reset; // @[RegFile.scala 66:20:@44111.4]
  wire [63:0] regs_463_io_in; // @[RegFile.scala 66:20:@44111.4]
  wire  regs_463_io_reset; // @[RegFile.scala 66:20:@44111.4]
  wire [63:0] regs_463_io_out; // @[RegFile.scala 66:20:@44111.4]
  wire  regs_463_io_enable; // @[RegFile.scala 66:20:@44111.4]
  wire  regs_464_clock; // @[RegFile.scala 66:20:@44125.4]
  wire  regs_464_reset; // @[RegFile.scala 66:20:@44125.4]
  wire [63:0] regs_464_io_in; // @[RegFile.scala 66:20:@44125.4]
  wire  regs_464_io_reset; // @[RegFile.scala 66:20:@44125.4]
  wire [63:0] regs_464_io_out; // @[RegFile.scala 66:20:@44125.4]
  wire  regs_464_io_enable; // @[RegFile.scala 66:20:@44125.4]
  wire  regs_465_clock; // @[RegFile.scala 66:20:@44139.4]
  wire  regs_465_reset; // @[RegFile.scala 66:20:@44139.4]
  wire [63:0] regs_465_io_in; // @[RegFile.scala 66:20:@44139.4]
  wire  regs_465_io_reset; // @[RegFile.scala 66:20:@44139.4]
  wire [63:0] regs_465_io_out; // @[RegFile.scala 66:20:@44139.4]
  wire  regs_465_io_enable; // @[RegFile.scala 66:20:@44139.4]
  wire  regs_466_clock; // @[RegFile.scala 66:20:@44153.4]
  wire  regs_466_reset; // @[RegFile.scala 66:20:@44153.4]
  wire [63:0] regs_466_io_in; // @[RegFile.scala 66:20:@44153.4]
  wire  regs_466_io_reset; // @[RegFile.scala 66:20:@44153.4]
  wire [63:0] regs_466_io_out; // @[RegFile.scala 66:20:@44153.4]
  wire  regs_466_io_enable; // @[RegFile.scala 66:20:@44153.4]
  wire  regs_467_clock; // @[RegFile.scala 66:20:@44167.4]
  wire  regs_467_reset; // @[RegFile.scala 66:20:@44167.4]
  wire [63:0] regs_467_io_in; // @[RegFile.scala 66:20:@44167.4]
  wire  regs_467_io_reset; // @[RegFile.scala 66:20:@44167.4]
  wire [63:0] regs_467_io_out; // @[RegFile.scala 66:20:@44167.4]
  wire  regs_467_io_enable; // @[RegFile.scala 66:20:@44167.4]
  wire  regs_468_clock; // @[RegFile.scala 66:20:@44181.4]
  wire  regs_468_reset; // @[RegFile.scala 66:20:@44181.4]
  wire [63:0] regs_468_io_in; // @[RegFile.scala 66:20:@44181.4]
  wire  regs_468_io_reset; // @[RegFile.scala 66:20:@44181.4]
  wire [63:0] regs_468_io_out; // @[RegFile.scala 66:20:@44181.4]
  wire  regs_468_io_enable; // @[RegFile.scala 66:20:@44181.4]
  wire  regs_469_clock; // @[RegFile.scala 66:20:@44195.4]
  wire  regs_469_reset; // @[RegFile.scala 66:20:@44195.4]
  wire [63:0] regs_469_io_in; // @[RegFile.scala 66:20:@44195.4]
  wire  regs_469_io_reset; // @[RegFile.scala 66:20:@44195.4]
  wire [63:0] regs_469_io_out; // @[RegFile.scala 66:20:@44195.4]
  wire  regs_469_io_enable; // @[RegFile.scala 66:20:@44195.4]
  wire  regs_470_clock; // @[RegFile.scala 66:20:@44209.4]
  wire  regs_470_reset; // @[RegFile.scala 66:20:@44209.4]
  wire [63:0] regs_470_io_in; // @[RegFile.scala 66:20:@44209.4]
  wire  regs_470_io_reset; // @[RegFile.scala 66:20:@44209.4]
  wire [63:0] regs_470_io_out; // @[RegFile.scala 66:20:@44209.4]
  wire  regs_470_io_enable; // @[RegFile.scala 66:20:@44209.4]
  wire  regs_471_clock; // @[RegFile.scala 66:20:@44223.4]
  wire  regs_471_reset; // @[RegFile.scala 66:20:@44223.4]
  wire [63:0] regs_471_io_in; // @[RegFile.scala 66:20:@44223.4]
  wire  regs_471_io_reset; // @[RegFile.scala 66:20:@44223.4]
  wire [63:0] regs_471_io_out; // @[RegFile.scala 66:20:@44223.4]
  wire  regs_471_io_enable; // @[RegFile.scala 66:20:@44223.4]
  wire  regs_472_clock; // @[RegFile.scala 66:20:@44237.4]
  wire  regs_472_reset; // @[RegFile.scala 66:20:@44237.4]
  wire [63:0] regs_472_io_in; // @[RegFile.scala 66:20:@44237.4]
  wire  regs_472_io_reset; // @[RegFile.scala 66:20:@44237.4]
  wire [63:0] regs_472_io_out; // @[RegFile.scala 66:20:@44237.4]
  wire  regs_472_io_enable; // @[RegFile.scala 66:20:@44237.4]
  wire  regs_473_clock; // @[RegFile.scala 66:20:@44251.4]
  wire  regs_473_reset; // @[RegFile.scala 66:20:@44251.4]
  wire [63:0] regs_473_io_in; // @[RegFile.scala 66:20:@44251.4]
  wire  regs_473_io_reset; // @[RegFile.scala 66:20:@44251.4]
  wire [63:0] regs_473_io_out; // @[RegFile.scala 66:20:@44251.4]
  wire  regs_473_io_enable; // @[RegFile.scala 66:20:@44251.4]
  wire  regs_474_clock; // @[RegFile.scala 66:20:@44265.4]
  wire  regs_474_reset; // @[RegFile.scala 66:20:@44265.4]
  wire [63:0] regs_474_io_in; // @[RegFile.scala 66:20:@44265.4]
  wire  regs_474_io_reset; // @[RegFile.scala 66:20:@44265.4]
  wire [63:0] regs_474_io_out; // @[RegFile.scala 66:20:@44265.4]
  wire  regs_474_io_enable; // @[RegFile.scala 66:20:@44265.4]
  wire  regs_475_clock; // @[RegFile.scala 66:20:@44279.4]
  wire  regs_475_reset; // @[RegFile.scala 66:20:@44279.4]
  wire [63:0] regs_475_io_in; // @[RegFile.scala 66:20:@44279.4]
  wire  regs_475_io_reset; // @[RegFile.scala 66:20:@44279.4]
  wire [63:0] regs_475_io_out; // @[RegFile.scala 66:20:@44279.4]
  wire  regs_475_io_enable; // @[RegFile.scala 66:20:@44279.4]
  wire  regs_476_clock; // @[RegFile.scala 66:20:@44293.4]
  wire  regs_476_reset; // @[RegFile.scala 66:20:@44293.4]
  wire [63:0] regs_476_io_in; // @[RegFile.scala 66:20:@44293.4]
  wire  regs_476_io_reset; // @[RegFile.scala 66:20:@44293.4]
  wire [63:0] regs_476_io_out; // @[RegFile.scala 66:20:@44293.4]
  wire  regs_476_io_enable; // @[RegFile.scala 66:20:@44293.4]
  wire  regs_477_clock; // @[RegFile.scala 66:20:@44307.4]
  wire  regs_477_reset; // @[RegFile.scala 66:20:@44307.4]
  wire [63:0] regs_477_io_in; // @[RegFile.scala 66:20:@44307.4]
  wire  regs_477_io_reset; // @[RegFile.scala 66:20:@44307.4]
  wire [63:0] regs_477_io_out; // @[RegFile.scala 66:20:@44307.4]
  wire  regs_477_io_enable; // @[RegFile.scala 66:20:@44307.4]
  wire  regs_478_clock; // @[RegFile.scala 66:20:@44321.4]
  wire  regs_478_reset; // @[RegFile.scala 66:20:@44321.4]
  wire [63:0] regs_478_io_in; // @[RegFile.scala 66:20:@44321.4]
  wire  regs_478_io_reset; // @[RegFile.scala 66:20:@44321.4]
  wire [63:0] regs_478_io_out; // @[RegFile.scala 66:20:@44321.4]
  wire  regs_478_io_enable; // @[RegFile.scala 66:20:@44321.4]
  wire  regs_479_clock; // @[RegFile.scala 66:20:@44335.4]
  wire  regs_479_reset; // @[RegFile.scala 66:20:@44335.4]
  wire [63:0] regs_479_io_in; // @[RegFile.scala 66:20:@44335.4]
  wire  regs_479_io_reset; // @[RegFile.scala 66:20:@44335.4]
  wire [63:0] regs_479_io_out; // @[RegFile.scala 66:20:@44335.4]
  wire  regs_479_io_enable; // @[RegFile.scala 66:20:@44335.4]
  wire  regs_480_clock; // @[RegFile.scala 66:20:@44349.4]
  wire  regs_480_reset; // @[RegFile.scala 66:20:@44349.4]
  wire [63:0] regs_480_io_in; // @[RegFile.scala 66:20:@44349.4]
  wire  regs_480_io_reset; // @[RegFile.scala 66:20:@44349.4]
  wire [63:0] regs_480_io_out; // @[RegFile.scala 66:20:@44349.4]
  wire  regs_480_io_enable; // @[RegFile.scala 66:20:@44349.4]
  wire  regs_481_clock; // @[RegFile.scala 66:20:@44363.4]
  wire  regs_481_reset; // @[RegFile.scala 66:20:@44363.4]
  wire [63:0] regs_481_io_in; // @[RegFile.scala 66:20:@44363.4]
  wire  regs_481_io_reset; // @[RegFile.scala 66:20:@44363.4]
  wire [63:0] regs_481_io_out; // @[RegFile.scala 66:20:@44363.4]
  wire  regs_481_io_enable; // @[RegFile.scala 66:20:@44363.4]
  wire  regs_482_clock; // @[RegFile.scala 66:20:@44377.4]
  wire  regs_482_reset; // @[RegFile.scala 66:20:@44377.4]
  wire [63:0] regs_482_io_in; // @[RegFile.scala 66:20:@44377.4]
  wire  regs_482_io_reset; // @[RegFile.scala 66:20:@44377.4]
  wire [63:0] regs_482_io_out; // @[RegFile.scala 66:20:@44377.4]
  wire  regs_482_io_enable; // @[RegFile.scala 66:20:@44377.4]
  wire  regs_483_clock; // @[RegFile.scala 66:20:@44391.4]
  wire  regs_483_reset; // @[RegFile.scala 66:20:@44391.4]
  wire [63:0] regs_483_io_in; // @[RegFile.scala 66:20:@44391.4]
  wire  regs_483_io_reset; // @[RegFile.scala 66:20:@44391.4]
  wire [63:0] regs_483_io_out; // @[RegFile.scala 66:20:@44391.4]
  wire  regs_483_io_enable; // @[RegFile.scala 66:20:@44391.4]
  wire  regs_484_clock; // @[RegFile.scala 66:20:@44405.4]
  wire  regs_484_reset; // @[RegFile.scala 66:20:@44405.4]
  wire [63:0] regs_484_io_in; // @[RegFile.scala 66:20:@44405.4]
  wire  regs_484_io_reset; // @[RegFile.scala 66:20:@44405.4]
  wire [63:0] regs_484_io_out; // @[RegFile.scala 66:20:@44405.4]
  wire  regs_484_io_enable; // @[RegFile.scala 66:20:@44405.4]
  wire  regs_485_clock; // @[RegFile.scala 66:20:@44419.4]
  wire  regs_485_reset; // @[RegFile.scala 66:20:@44419.4]
  wire [63:0] regs_485_io_in; // @[RegFile.scala 66:20:@44419.4]
  wire  regs_485_io_reset; // @[RegFile.scala 66:20:@44419.4]
  wire [63:0] regs_485_io_out; // @[RegFile.scala 66:20:@44419.4]
  wire  regs_485_io_enable; // @[RegFile.scala 66:20:@44419.4]
  wire  regs_486_clock; // @[RegFile.scala 66:20:@44433.4]
  wire  regs_486_reset; // @[RegFile.scala 66:20:@44433.4]
  wire [63:0] regs_486_io_in; // @[RegFile.scala 66:20:@44433.4]
  wire  regs_486_io_reset; // @[RegFile.scala 66:20:@44433.4]
  wire [63:0] regs_486_io_out; // @[RegFile.scala 66:20:@44433.4]
  wire  regs_486_io_enable; // @[RegFile.scala 66:20:@44433.4]
  wire  regs_487_clock; // @[RegFile.scala 66:20:@44447.4]
  wire  regs_487_reset; // @[RegFile.scala 66:20:@44447.4]
  wire [63:0] regs_487_io_in; // @[RegFile.scala 66:20:@44447.4]
  wire  regs_487_io_reset; // @[RegFile.scala 66:20:@44447.4]
  wire [63:0] regs_487_io_out; // @[RegFile.scala 66:20:@44447.4]
  wire  regs_487_io_enable; // @[RegFile.scala 66:20:@44447.4]
  wire  regs_488_clock; // @[RegFile.scala 66:20:@44461.4]
  wire  regs_488_reset; // @[RegFile.scala 66:20:@44461.4]
  wire [63:0] regs_488_io_in; // @[RegFile.scala 66:20:@44461.4]
  wire  regs_488_io_reset; // @[RegFile.scala 66:20:@44461.4]
  wire [63:0] regs_488_io_out; // @[RegFile.scala 66:20:@44461.4]
  wire  regs_488_io_enable; // @[RegFile.scala 66:20:@44461.4]
  wire  regs_489_clock; // @[RegFile.scala 66:20:@44475.4]
  wire  regs_489_reset; // @[RegFile.scala 66:20:@44475.4]
  wire [63:0] regs_489_io_in; // @[RegFile.scala 66:20:@44475.4]
  wire  regs_489_io_reset; // @[RegFile.scala 66:20:@44475.4]
  wire [63:0] regs_489_io_out; // @[RegFile.scala 66:20:@44475.4]
  wire  regs_489_io_enable; // @[RegFile.scala 66:20:@44475.4]
  wire  regs_490_clock; // @[RegFile.scala 66:20:@44489.4]
  wire  regs_490_reset; // @[RegFile.scala 66:20:@44489.4]
  wire [63:0] regs_490_io_in; // @[RegFile.scala 66:20:@44489.4]
  wire  regs_490_io_reset; // @[RegFile.scala 66:20:@44489.4]
  wire [63:0] regs_490_io_out; // @[RegFile.scala 66:20:@44489.4]
  wire  regs_490_io_enable; // @[RegFile.scala 66:20:@44489.4]
  wire  regs_491_clock; // @[RegFile.scala 66:20:@44503.4]
  wire  regs_491_reset; // @[RegFile.scala 66:20:@44503.4]
  wire [63:0] regs_491_io_in; // @[RegFile.scala 66:20:@44503.4]
  wire  regs_491_io_reset; // @[RegFile.scala 66:20:@44503.4]
  wire [63:0] regs_491_io_out; // @[RegFile.scala 66:20:@44503.4]
  wire  regs_491_io_enable; // @[RegFile.scala 66:20:@44503.4]
  wire  regs_492_clock; // @[RegFile.scala 66:20:@44517.4]
  wire  regs_492_reset; // @[RegFile.scala 66:20:@44517.4]
  wire [63:0] regs_492_io_in; // @[RegFile.scala 66:20:@44517.4]
  wire  regs_492_io_reset; // @[RegFile.scala 66:20:@44517.4]
  wire [63:0] regs_492_io_out; // @[RegFile.scala 66:20:@44517.4]
  wire  regs_492_io_enable; // @[RegFile.scala 66:20:@44517.4]
  wire  regs_493_clock; // @[RegFile.scala 66:20:@44531.4]
  wire  regs_493_reset; // @[RegFile.scala 66:20:@44531.4]
  wire [63:0] regs_493_io_in; // @[RegFile.scala 66:20:@44531.4]
  wire  regs_493_io_reset; // @[RegFile.scala 66:20:@44531.4]
  wire [63:0] regs_493_io_out; // @[RegFile.scala 66:20:@44531.4]
  wire  regs_493_io_enable; // @[RegFile.scala 66:20:@44531.4]
  wire  regs_494_clock; // @[RegFile.scala 66:20:@44545.4]
  wire  regs_494_reset; // @[RegFile.scala 66:20:@44545.4]
  wire [63:0] regs_494_io_in; // @[RegFile.scala 66:20:@44545.4]
  wire  regs_494_io_reset; // @[RegFile.scala 66:20:@44545.4]
  wire [63:0] regs_494_io_out; // @[RegFile.scala 66:20:@44545.4]
  wire  regs_494_io_enable; // @[RegFile.scala 66:20:@44545.4]
  wire  regs_495_clock; // @[RegFile.scala 66:20:@44559.4]
  wire  regs_495_reset; // @[RegFile.scala 66:20:@44559.4]
  wire [63:0] regs_495_io_in; // @[RegFile.scala 66:20:@44559.4]
  wire  regs_495_io_reset; // @[RegFile.scala 66:20:@44559.4]
  wire [63:0] regs_495_io_out; // @[RegFile.scala 66:20:@44559.4]
  wire  regs_495_io_enable; // @[RegFile.scala 66:20:@44559.4]
  wire  regs_496_clock; // @[RegFile.scala 66:20:@44573.4]
  wire  regs_496_reset; // @[RegFile.scala 66:20:@44573.4]
  wire [63:0] regs_496_io_in; // @[RegFile.scala 66:20:@44573.4]
  wire  regs_496_io_reset; // @[RegFile.scala 66:20:@44573.4]
  wire [63:0] regs_496_io_out; // @[RegFile.scala 66:20:@44573.4]
  wire  regs_496_io_enable; // @[RegFile.scala 66:20:@44573.4]
  wire  regs_497_clock; // @[RegFile.scala 66:20:@44587.4]
  wire  regs_497_reset; // @[RegFile.scala 66:20:@44587.4]
  wire [63:0] regs_497_io_in; // @[RegFile.scala 66:20:@44587.4]
  wire  regs_497_io_reset; // @[RegFile.scala 66:20:@44587.4]
  wire [63:0] regs_497_io_out; // @[RegFile.scala 66:20:@44587.4]
  wire  regs_497_io_enable; // @[RegFile.scala 66:20:@44587.4]
  wire  regs_498_clock; // @[RegFile.scala 66:20:@44601.4]
  wire  regs_498_reset; // @[RegFile.scala 66:20:@44601.4]
  wire [63:0] regs_498_io_in; // @[RegFile.scala 66:20:@44601.4]
  wire  regs_498_io_reset; // @[RegFile.scala 66:20:@44601.4]
  wire [63:0] regs_498_io_out; // @[RegFile.scala 66:20:@44601.4]
  wire  regs_498_io_enable; // @[RegFile.scala 66:20:@44601.4]
  wire  regs_499_clock; // @[RegFile.scala 66:20:@44615.4]
  wire  regs_499_reset; // @[RegFile.scala 66:20:@44615.4]
  wire [63:0] regs_499_io_in; // @[RegFile.scala 66:20:@44615.4]
  wire  regs_499_io_reset; // @[RegFile.scala 66:20:@44615.4]
  wire [63:0] regs_499_io_out; // @[RegFile.scala 66:20:@44615.4]
  wire  regs_499_io_enable; // @[RegFile.scala 66:20:@44615.4]
  wire  regs_500_clock; // @[RegFile.scala 66:20:@44629.4]
  wire  regs_500_reset; // @[RegFile.scala 66:20:@44629.4]
  wire [63:0] regs_500_io_in; // @[RegFile.scala 66:20:@44629.4]
  wire  regs_500_io_reset; // @[RegFile.scala 66:20:@44629.4]
  wire [63:0] regs_500_io_out; // @[RegFile.scala 66:20:@44629.4]
  wire  regs_500_io_enable; // @[RegFile.scala 66:20:@44629.4]
  wire  regs_501_clock; // @[RegFile.scala 66:20:@44643.4]
  wire  regs_501_reset; // @[RegFile.scala 66:20:@44643.4]
  wire [63:0] regs_501_io_in; // @[RegFile.scala 66:20:@44643.4]
  wire  regs_501_io_reset; // @[RegFile.scala 66:20:@44643.4]
  wire [63:0] regs_501_io_out; // @[RegFile.scala 66:20:@44643.4]
  wire  regs_501_io_enable; // @[RegFile.scala 66:20:@44643.4]
  wire  regs_502_clock; // @[RegFile.scala 66:20:@44657.4]
  wire  regs_502_reset; // @[RegFile.scala 66:20:@44657.4]
  wire [63:0] regs_502_io_in; // @[RegFile.scala 66:20:@44657.4]
  wire  regs_502_io_reset; // @[RegFile.scala 66:20:@44657.4]
  wire [63:0] regs_502_io_out; // @[RegFile.scala 66:20:@44657.4]
  wire  regs_502_io_enable; // @[RegFile.scala 66:20:@44657.4]
  wire  regs_503_clock; // @[RegFile.scala 66:20:@44671.4]
  wire  regs_503_reset; // @[RegFile.scala 66:20:@44671.4]
  wire [63:0] regs_503_io_in; // @[RegFile.scala 66:20:@44671.4]
  wire  regs_503_io_reset; // @[RegFile.scala 66:20:@44671.4]
  wire [63:0] regs_503_io_out; // @[RegFile.scala 66:20:@44671.4]
  wire  regs_503_io_enable; // @[RegFile.scala 66:20:@44671.4]
  wire  regs_504_clock; // @[RegFile.scala 66:20:@44685.4]
  wire  regs_504_reset; // @[RegFile.scala 66:20:@44685.4]
  wire [63:0] regs_504_io_in; // @[RegFile.scala 66:20:@44685.4]
  wire  regs_504_io_reset; // @[RegFile.scala 66:20:@44685.4]
  wire [63:0] regs_504_io_out; // @[RegFile.scala 66:20:@44685.4]
  wire  regs_504_io_enable; // @[RegFile.scala 66:20:@44685.4]
  wire  regs_505_clock; // @[RegFile.scala 66:20:@44699.4]
  wire  regs_505_reset; // @[RegFile.scala 66:20:@44699.4]
  wire [63:0] regs_505_io_in; // @[RegFile.scala 66:20:@44699.4]
  wire  regs_505_io_reset; // @[RegFile.scala 66:20:@44699.4]
  wire [63:0] regs_505_io_out; // @[RegFile.scala 66:20:@44699.4]
  wire  regs_505_io_enable; // @[RegFile.scala 66:20:@44699.4]
  wire  regs_506_clock; // @[RegFile.scala 66:20:@44713.4]
  wire  regs_506_reset; // @[RegFile.scala 66:20:@44713.4]
  wire [63:0] regs_506_io_in; // @[RegFile.scala 66:20:@44713.4]
  wire  regs_506_io_reset; // @[RegFile.scala 66:20:@44713.4]
  wire [63:0] regs_506_io_out; // @[RegFile.scala 66:20:@44713.4]
  wire  regs_506_io_enable; // @[RegFile.scala 66:20:@44713.4]
  wire  regs_507_clock; // @[RegFile.scala 66:20:@44727.4]
  wire  regs_507_reset; // @[RegFile.scala 66:20:@44727.4]
  wire [63:0] regs_507_io_in; // @[RegFile.scala 66:20:@44727.4]
  wire  regs_507_io_reset; // @[RegFile.scala 66:20:@44727.4]
  wire [63:0] regs_507_io_out; // @[RegFile.scala 66:20:@44727.4]
  wire  regs_507_io_enable; // @[RegFile.scala 66:20:@44727.4]
  wire  regs_508_clock; // @[RegFile.scala 66:20:@44741.4]
  wire  regs_508_reset; // @[RegFile.scala 66:20:@44741.4]
  wire [63:0] regs_508_io_in; // @[RegFile.scala 66:20:@44741.4]
  wire  regs_508_io_reset; // @[RegFile.scala 66:20:@44741.4]
  wire [63:0] regs_508_io_out; // @[RegFile.scala 66:20:@44741.4]
  wire  regs_508_io_enable; // @[RegFile.scala 66:20:@44741.4]
  wire  regs_509_clock; // @[RegFile.scala 66:20:@44755.4]
  wire  regs_509_reset; // @[RegFile.scala 66:20:@44755.4]
  wire [63:0] regs_509_io_in; // @[RegFile.scala 66:20:@44755.4]
  wire  regs_509_io_reset; // @[RegFile.scala 66:20:@44755.4]
  wire [63:0] regs_509_io_out; // @[RegFile.scala 66:20:@44755.4]
  wire  regs_509_io_enable; // @[RegFile.scala 66:20:@44755.4]
  wire  regs_510_clock; // @[RegFile.scala 66:20:@44769.4]
  wire  regs_510_reset; // @[RegFile.scala 66:20:@44769.4]
  wire [63:0] regs_510_io_in; // @[RegFile.scala 66:20:@44769.4]
  wire  regs_510_io_reset; // @[RegFile.scala 66:20:@44769.4]
  wire [63:0] regs_510_io_out; // @[RegFile.scala 66:20:@44769.4]
  wire  regs_510_io_enable; // @[RegFile.scala 66:20:@44769.4]
  wire  regs_511_clock; // @[RegFile.scala 66:20:@44783.4]
  wire  regs_511_reset; // @[RegFile.scala 66:20:@44783.4]
  wire [63:0] regs_511_io_in; // @[RegFile.scala 66:20:@44783.4]
  wire  regs_511_io_reset; // @[RegFile.scala 66:20:@44783.4]
  wire [63:0] regs_511_io_out; // @[RegFile.scala 66:20:@44783.4]
  wire  regs_511_io_enable; // @[RegFile.scala 66:20:@44783.4]
  wire [63:0] rport_io_ins_0; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_1; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_2; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_3; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_4; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_5; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_6; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_7; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_8; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_9; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_10; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_11; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_12; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_13; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_14; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_15; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_16; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_17; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_18; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_19; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_20; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_21; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_22; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_23; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_24; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_25; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_26; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_27; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_28; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_29; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_30; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_31; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_32; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_33; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_34; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_35; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_36; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_37; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_38; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_39; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_40; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_41; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_42; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_43; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_44; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_45; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_46; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_47; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_48; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_49; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_50; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_51; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_52; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_53; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_54; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_55; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_56; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_57; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_58; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_59; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_60; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_61; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_62; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_63; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_64; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_65; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_66; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_67; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_68; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_69; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_70; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_71; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_72; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_73; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_74; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_75; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_76; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_77; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_78; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_79; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_80; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_81; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_82; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_83; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_84; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_85; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_86; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_87; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_88; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_89; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_90; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_91; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_92; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_93; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_94; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_95; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_96; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_97; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_98; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_99; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_100; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_101; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_102; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_103; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_104; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_105; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_106; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_107; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_108; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_109; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_110; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_111; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_112; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_113; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_114; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_115; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_116; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_117; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_118; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_119; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_120; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_121; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_122; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_123; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_124; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_125; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_126; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_127; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_128; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_129; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_130; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_131; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_132; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_133; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_134; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_135; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_136; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_137; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_138; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_139; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_140; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_141; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_142; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_143; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_144; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_145; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_146; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_147; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_148; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_149; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_150; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_151; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_152; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_153; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_154; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_155; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_156; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_157; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_158; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_159; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_160; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_161; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_162; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_163; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_164; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_165; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_166; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_167; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_168; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_169; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_170; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_171; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_172; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_173; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_174; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_175; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_176; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_177; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_178; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_179; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_180; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_181; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_182; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_183; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_184; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_185; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_186; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_187; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_188; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_189; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_190; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_191; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_192; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_193; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_194; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_195; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_196; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_197; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_198; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_199; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_200; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_201; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_202; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_203; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_204; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_205; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_206; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_207; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_208; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_209; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_210; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_211; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_212; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_213; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_214; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_215; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_216; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_217; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_218; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_219; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_220; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_221; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_222; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_223; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_224; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_225; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_226; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_227; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_228; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_229; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_230; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_231; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_232; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_233; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_234; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_235; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_236; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_237; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_238; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_239; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_240; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_241; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_242; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_243; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_244; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_245; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_246; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_247; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_248; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_249; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_250; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_251; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_252; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_253; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_254; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_255; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_256; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_257; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_258; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_259; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_260; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_261; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_262; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_263; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_264; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_265; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_266; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_267; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_268; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_269; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_270; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_271; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_272; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_273; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_274; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_275; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_276; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_277; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_278; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_279; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_280; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_281; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_282; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_283; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_284; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_285; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_286; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_287; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_288; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_289; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_290; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_291; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_292; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_293; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_294; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_295; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_296; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_297; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_298; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_299; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_300; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_301; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_302; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_303; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_304; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_305; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_306; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_307; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_308; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_309; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_310; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_311; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_312; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_313; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_314; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_315; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_316; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_317; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_318; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_319; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_320; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_321; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_322; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_323; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_324; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_325; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_326; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_327; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_328; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_329; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_330; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_331; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_332; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_333; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_334; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_335; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_336; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_337; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_338; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_339; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_340; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_341; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_342; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_343; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_344; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_345; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_346; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_347; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_348; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_349; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_350; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_351; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_352; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_353; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_354; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_355; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_356; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_357; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_358; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_359; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_360; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_361; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_362; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_363; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_364; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_365; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_366; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_367; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_368; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_369; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_370; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_371; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_372; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_373; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_374; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_375; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_376; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_377; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_378; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_379; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_380; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_381; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_382; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_383; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_384; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_385; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_386; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_387; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_388; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_389; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_390; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_391; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_392; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_393; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_394; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_395; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_396; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_397; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_398; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_399; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_400; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_401; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_402; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_403; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_404; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_405; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_406; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_407; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_408; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_409; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_410; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_411; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_412; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_413; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_414; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_415; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_416; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_417; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_418; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_419; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_420; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_421; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_422; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_423; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_424; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_425; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_426; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_427; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_428; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_429; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_430; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_431; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_432; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_433; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_434; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_435; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_436; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_437; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_438; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_439; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_440; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_441; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_442; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_443; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_444; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_445; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_446; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_447; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_448; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_449; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_450; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_451; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_452; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_453; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_454; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_455; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_456; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_457; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_458; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_459; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_460; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_461; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_462; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_463; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_464; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_465; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_466; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_467; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_468; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_469; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_470; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_471; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_472; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_473; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_474; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_475; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_476; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_477; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_478; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_479; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_480; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_481; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_482; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_483; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_484; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_485; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_486; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_487; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_488; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_489; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_490; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_491; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_492; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_493; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_494; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_495; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_496; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_497; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_498; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_499; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_500; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_501; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_502; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_503; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_504; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_505; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_506; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_507; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_508; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_509; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_510; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_ins_511; // @[RegFile.scala 95:21:@44797.4]
  wire [8:0] rport_io_sel; // @[RegFile.scala 95:21:@44797.4]
  wire [63:0] rport_io_out; // @[RegFile.scala 95:21:@44797.4]
  wire  _T_3130; // @[RegFile.scala 80:42:@37631.4]
  wire  _T_3136; // @[RegFile.scala 68:46:@37643.4]
  wire  _T_3137; // @[RegFile.scala 68:34:@37644.4]
  wire  _T_3150; // @[RegFile.scala 80:42:@37662.4]
  wire  _T_3156; // @[RegFile.scala 74:80:@37674.4]
  wire  _T_3157; // @[RegFile.scala 74:68:@37675.4]
  wire  _T_3163; // @[RegFile.scala 74:80:@37688.4]
  wire  _T_3164; // @[RegFile.scala 74:68:@37689.4]
  wire  _T_3170; // @[RegFile.scala 74:80:@37702.4]
  wire  _T_3171; // @[RegFile.scala 74:68:@37703.4]
  wire  _T_3177; // @[RegFile.scala 74:80:@37716.4]
  wire  _T_3178; // @[RegFile.scala 74:68:@37717.4]
  wire  _T_3184; // @[RegFile.scala 74:80:@37730.4]
  wire  _T_3185; // @[RegFile.scala 74:68:@37731.4]
  wire  _T_3191; // @[RegFile.scala 74:80:@37744.4]
  wire  _T_3192; // @[RegFile.scala 74:68:@37745.4]
  wire  _T_3198; // @[RegFile.scala 74:80:@37758.4]
  wire  _T_3199; // @[RegFile.scala 74:68:@37759.4]
  wire  _T_3205; // @[RegFile.scala 74:80:@37772.4]
  wire  _T_3206; // @[RegFile.scala 74:68:@37773.4]
  wire  _T_3212; // @[RegFile.scala 74:80:@37786.4]
  wire  _T_3213; // @[RegFile.scala 74:68:@37787.4]
  wire  _T_3219; // @[RegFile.scala 74:80:@37800.4]
  wire  _T_3220; // @[RegFile.scala 74:68:@37801.4]
  FringeFF regs_0 ( // @[RegFile.scala 66:20:@37628.4]
    .clock(regs_0_clock),
    .reset(regs_0_reset),
    .io_in(regs_0_io_in),
    .io_reset(regs_0_io_reset),
    .io_out(regs_0_io_out),
    .io_enable(regs_0_io_enable)
  );
  FringeFF regs_1 ( // @[RegFile.scala 66:20:@37640.4]
    .clock(regs_1_clock),
    .reset(regs_1_reset),
    .io_in(regs_1_io_in),
    .io_reset(regs_1_io_reset),
    .io_out(regs_1_io_out),
    .io_enable(regs_1_io_enable)
  );
  FringeFF regs_2 ( // @[RegFile.scala 66:20:@37659.4]
    .clock(regs_2_clock),
    .reset(regs_2_reset),
    .io_in(regs_2_io_in),
    .io_reset(regs_2_io_reset),
    .io_out(regs_2_io_out),
    .io_enable(regs_2_io_enable)
  );
  FringeFF regs_3 ( // @[RegFile.scala 66:20:@37671.4]
    .clock(regs_3_clock),
    .reset(regs_3_reset),
    .io_in(regs_3_io_in),
    .io_reset(regs_3_io_reset),
    .io_out(regs_3_io_out),
    .io_enable(regs_3_io_enable)
  );
  FringeFF regs_4 ( // @[RegFile.scala 66:20:@37685.4]
    .clock(regs_4_clock),
    .reset(regs_4_reset),
    .io_in(regs_4_io_in),
    .io_reset(regs_4_io_reset),
    .io_out(regs_4_io_out),
    .io_enable(regs_4_io_enable)
  );
  FringeFF regs_5 ( // @[RegFile.scala 66:20:@37699.4]
    .clock(regs_5_clock),
    .reset(regs_5_reset),
    .io_in(regs_5_io_in),
    .io_reset(regs_5_io_reset),
    .io_out(regs_5_io_out),
    .io_enable(regs_5_io_enable)
  );
  FringeFF regs_6 ( // @[RegFile.scala 66:20:@37713.4]
    .clock(regs_6_clock),
    .reset(regs_6_reset),
    .io_in(regs_6_io_in),
    .io_reset(regs_6_io_reset),
    .io_out(regs_6_io_out),
    .io_enable(regs_6_io_enable)
  );
  FringeFF regs_7 ( // @[RegFile.scala 66:20:@37727.4]
    .clock(regs_7_clock),
    .reset(regs_7_reset),
    .io_in(regs_7_io_in),
    .io_reset(regs_7_io_reset),
    .io_out(regs_7_io_out),
    .io_enable(regs_7_io_enable)
  );
  FringeFF regs_8 ( // @[RegFile.scala 66:20:@37741.4]
    .clock(regs_8_clock),
    .reset(regs_8_reset),
    .io_in(regs_8_io_in),
    .io_reset(regs_8_io_reset),
    .io_out(regs_8_io_out),
    .io_enable(regs_8_io_enable)
  );
  FringeFF regs_9 ( // @[RegFile.scala 66:20:@37755.4]
    .clock(regs_9_clock),
    .reset(regs_9_reset),
    .io_in(regs_9_io_in),
    .io_reset(regs_9_io_reset),
    .io_out(regs_9_io_out),
    .io_enable(regs_9_io_enable)
  );
  FringeFF regs_10 ( // @[RegFile.scala 66:20:@37769.4]
    .clock(regs_10_clock),
    .reset(regs_10_reset),
    .io_in(regs_10_io_in),
    .io_reset(regs_10_io_reset),
    .io_out(regs_10_io_out),
    .io_enable(regs_10_io_enable)
  );
  FringeFF regs_11 ( // @[RegFile.scala 66:20:@37783.4]
    .clock(regs_11_clock),
    .reset(regs_11_reset),
    .io_in(regs_11_io_in),
    .io_reset(regs_11_io_reset),
    .io_out(regs_11_io_out),
    .io_enable(regs_11_io_enable)
  );
  FringeFF regs_12 ( // @[RegFile.scala 66:20:@37797.4]
    .clock(regs_12_clock),
    .reset(regs_12_reset),
    .io_in(regs_12_io_in),
    .io_reset(regs_12_io_reset),
    .io_out(regs_12_io_out),
    .io_enable(regs_12_io_enable)
  );
  FringeFF regs_13 ( // @[RegFile.scala 66:20:@37811.4]
    .clock(regs_13_clock),
    .reset(regs_13_reset),
    .io_in(regs_13_io_in),
    .io_reset(regs_13_io_reset),
    .io_out(regs_13_io_out),
    .io_enable(regs_13_io_enable)
  );
  FringeFF regs_14 ( // @[RegFile.scala 66:20:@37825.4]
    .clock(regs_14_clock),
    .reset(regs_14_reset),
    .io_in(regs_14_io_in),
    .io_reset(regs_14_io_reset),
    .io_out(regs_14_io_out),
    .io_enable(regs_14_io_enable)
  );
  FringeFF regs_15 ( // @[RegFile.scala 66:20:@37839.4]
    .clock(regs_15_clock),
    .reset(regs_15_reset),
    .io_in(regs_15_io_in),
    .io_reset(regs_15_io_reset),
    .io_out(regs_15_io_out),
    .io_enable(regs_15_io_enable)
  );
  FringeFF regs_16 ( // @[RegFile.scala 66:20:@37853.4]
    .clock(regs_16_clock),
    .reset(regs_16_reset),
    .io_in(regs_16_io_in),
    .io_reset(regs_16_io_reset),
    .io_out(regs_16_io_out),
    .io_enable(regs_16_io_enable)
  );
  FringeFF regs_17 ( // @[RegFile.scala 66:20:@37867.4]
    .clock(regs_17_clock),
    .reset(regs_17_reset),
    .io_in(regs_17_io_in),
    .io_reset(regs_17_io_reset),
    .io_out(regs_17_io_out),
    .io_enable(regs_17_io_enable)
  );
  FringeFF regs_18 ( // @[RegFile.scala 66:20:@37881.4]
    .clock(regs_18_clock),
    .reset(regs_18_reset),
    .io_in(regs_18_io_in),
    .io_reset(regs_18_io_reset),
    .io_out(regs_18_io_out),
    .io_enable(regs_18_io_enable)
  );
  FringeFF regs_19 ( // @[RegFile.scala 66:20:@37895.4]
    .clock(regs_19_clock),
    .reset(regs_19_reset),
    .io_in(regs_19_io_in),
    .io_reset(regs_19_io_reset),
    .io_out(regs_19_io_out),
    .io_enable(regs_19_io_enable)
  );
  FringeFF regs_20 ( // @[RegFile.scala 66:20:@37909.4]
    .clock(regs_20_clock),
    .reset(regs_20_reset),
    .io_in(regs_20_io_in),
    .io_reset(regs_20_io_reset),
    .io_out(regs_20_io_out),
    .io_enable(regs_20_io_enable)
  );
  FringeFF regs_21 ( // @[RegFile.scala 66:20:@37923.4]
    .clock(regs_21_clock),
    .reset(regs_21_reset),
    .io_in(regs_21_io_in),
    .io_reset(regs_21_io_reset),
    .io_out(regs_21_io_out),
    .io_enable(regs_21_io_enable)
  );
  FringeFF regs_22 ( // @[RegFile.scala 66:20:@37937.4]
    .clock(regs_22_clock),
    .reset(regs_22_reset),
    .io_in(regs_22_io_in),
    .io_reset(regs_22_io_reset),
    .io_out(regs_22_io_out),
    .io_enable(regs_22_io_enable)
  );
  FringeFF regs_23 ( // @[RegFile.scala 66:20:@37951.4]
    .clock(regs_23_clock),
    .reset(regs_23_reset),
    .io_in(regs_23_io_in),
    .io_reset(regs_23_io_reset),
    .io_out(regs_23_io_out),
    .io_enable(regs_23_io_enable)
  );
  FringeFF regs_24 ( // @[RegFile.scala 66:20:@37965.4]
    .clock(regs_24_clock),
    .reset(regs_24_reset),
    .io_in(regs_24_io_in),
    .io_reset(regs_24_io_reset),
    .io_out(regs_24_io_out),
    .io_enable(regs_24_io_enable)
  );
  FringeFF regs_25 ( // @[RegFile.scala 66:20:@37979.4]
    .clock(regs_25_clock),
    .reset(regs_25_reset),
    .io_in(regs_25_io_in),
    .io_reset(regs_25_io_reset),
    .io_out(regs_25_io_out),
    .io_enable(regs_25_io_enable)
  );
  FringeFF regs_26 ( // @[RegFile.scala 66:20:@37993.4]
    .clock(regs_26_clock),
    .reset(regs_26_reset),
    .io_in(regs_26_io_in),
    .io_reset(regs_26_io_reset),
    .io_out(regs_26_io_out),
    .io_enable(regs_26_io_enable)
  );
  FringeFF regs_27 ( // @[RegFile.scala 66:20:@38007.4]
    .clock(regs_27_clock),
    .reset(regs_27_reset),
    .io_in(regs_27_io_in),
    .io_reset(regs_27_io_reset),
    .io_out(regs_27_io_out),
    .io_enable(regs_27_io_enable)
  );
  FringeFF regs_28 ( // @[RegFile.scala 66:20:@38021.4]
    .clock(regs_28_clock),
    .reset(regs_28_reset),
    .io_in(regs_28_io_in),
    .io_reset(regs_28_io_reset),
    .io_out(regs_28_io_out),
    .io_enable(regs_28_io_enable)
  );
  FringeFF regs_29 ( // @[RegFile.scala 66:20:@38035.4]
    .clock(regs_29_clock),
    .reset(regs_29_reset),
    .io_in(regs_29_io_in),
    .io_reset(regs_29_io_reset),
    .io_out(regs_29_io_out),
    .io_enable(regs_29_io_enable)
  );
  FringeFF regs_30 ( // @[RegFile.scala 66:20:@38049.4]
    .clock(regs_30_clock),
    .reset(regs_30_reset),
    .io_in(regs_30_io_in),
    .io_reset(regs_30_io_reset),
    .io_out(regs_30_io_out),
    .io_enable(regs_30_io_enable)
  );
  FringeFF regs_31 ( // @[RegFile.scala 66:20:@38063.4]
    .clock(regs_31_clock),
    .reset(regs_31_reset),
    .io_in(regs_31_io_in),
    .io_reset(regs_31_io_reset),
    .io_out(regs_31_io_out),
    .io_enable(regs_31_io_enable)
  );
  FringeFF regs_32 ( // @[RegFile.scala 66:20:@38077.4]
    .clock(regs_32_clock),
    .reset(regs_32_reset),
    .io_in(regs_32_io_in),
    .io_reset(regs_32_io_reset),
    .io_out(regs_32_io_out),
    .io_enable(regs_32_io_enable)
  );
  FringeFF regs_33 ( // @[RegFile.scala 66:20:@38091.4]
    .clock(regs_33_clock),
    .reset(regs_33_reset),
    .io_in(regs_33_io_in),
    .io_reset(regs_33_io_reset),
    .io_out(regs_33_io_out),
    .io_enable(regs_33_io_enable)
  );
  FringeFF regs_34 ( // @[RegFile.scala 66:20:@38105.4]
    .clock(regs_34_clock),
    .reset(regs_34_reset),
    .io_in(regs_34_io_in),
    .io_reset(regs_34_io_reset),
    .io_out(regs_34_io_out),
    .io_enable(regs_34_io_enable)
  );
  FringeFF regs_35 ( // @[RegFile.scala 66:20:@38119.4]
    .clock(regs_35_clock),
    .reset(regs_35_reset),
    .io_in(regs_35_io_in),
    .io_reset(regs_35_io_reset),
    .io_out(regs_35_io_out),
    .io_enable(regs_35_io_enable)
  );
  FringeFF regs_36 ( // @[RegFile.scala 66:20:@38133.4]
    .clock(regs_36_clock),
    .reset(regs_36_reset),
    .io_in(regs_36_io_in),
    .io_reset(regs_36_io_reset),
    .io_out(regs_36_io_out),
    .io_enable(regs_36_io_enable)
  );
  FringeFF regs_37 ( // @[RegFile.scala 66:20:@38147.4]
    .clock(regs_37_clock),
    .reset(regs_37_reset),
    .io_in(regs_37_io_in),
    .io_reset(regs_37_io_reset),
    .io_out(regs_37_io_out),
    .io_enable(regs_37_io_enable)
  );
  FringeFF regs_38 ( // @[RegFile.scala 66:20:@38161.4]
    .clock(regs_38_clock),
    .reset(regs_38_reset),
    .io_in(regs_38_io_in),
    .io_reset(regs_38_io_reset),
    .io_out(regs_38_io_out),
    .io_enable(regs_38_io_enable)
  );
  FringeFF regs_39 ( // @[RegFile.scala 66:20:@38175.4]
    .clock(regs_39_clock),
    .reset(regs_39_reset),
    .io_in(regs_39_io_in),
    .io_reset(regs_39_io_reset),
    .io_out(regs_39_io_out),
    .io_enable(regs_39_io_enable)
  );
  FringeFF regs_40 ( // @[RegFile.scala 66:20:@38189.4]
    .clock(regs_40_clock),
    .reset(regs_40_reset),
    .io_in(regs_40_io_in),
    .io_reset(regs_40_io_reset),
    .io_out(regs_40_io_out),
    .io_enable(regs_40_io_enable)
  );
  FringeFF regs_41 ( // @[RegFile.scala 66:20:@38203.4]
    .clock(regs_41_clock),
    .reset(regs_41_reset),
    .io_in(regs_41_io_in),
    .io_reset(regs_41_io_reset),
    .io_out(regs_41_io_out),
    .io_enable(regs_41_io_enable)
  );
  FringeFF regs_42 ( // @[RegFile.scala 66:20:@38217.4]
    .clock(regs_42_clock),
    .reset(regs_42_reset),
    .io_in(regs_42_io_in),
    .io_reset(regs_42_io_reset),
    .io_out(regs_42_io_out),
    .io_enable(regs_42_io_enable)
  );
  FringeFF regs_43 ( // @[RegFile.scala 66:20:@38231.4]
    .clock(regs_43_clock),
    .reset(regs_43_reset),
    .io_in(regs_43_io_in),
    .io_reset(regs_43_io_reset),
    .io_out(regs_43_io_out),
    .io_enable(regs_43_io_enable)
  );
  FringeFF regs_44 ( // @[RegFile.scala 66:20:@38245.4]
    .clock(regs_44_clock),
    .reset(regs_44_reset),
    .io_in(regs_44_io_in),
    .io_reset(regs_44_io_reset),
    .io_out(regs_44_io_out),
    .io_enable(regs_44_io_enable)
  );
  FringeFF regs_45 ( // @[RegFile.scala 66:20:@38259.4]
    .clock(regs_45_clock),
    .reset(regs_45_reset),
    .io_in(regs_45_io_in),
    .io_reset(regs_45_io_reset),
    .io_out(regs_45_io_out),
    .io_enable(regs_45_io_enable)
  );
  FringeFF regs_46 ( // @[RegFile.scala 66:20:@38273.4]
    .clock(regs_46_clock),
    .reset(regs_46_reset),
    .io_in(regs_46_io_in),
    .io_reset(regs_46_io_reset),
    .io_out(regs_46_io_out),
    .io_enable(regs_46_io_enable)
  );
  FringeFF regs_47 ( // @[RegFile.scala 66:20:@38287.4]
    .clock(regs_47_clock),
    .reset(regs_47_reset),
    .io_in(regs_47_io_in),
    .io_reset(regs_47_io_reset),
    .io_out(regs_47_io_out),
    .io_enable(regs_47_io_enable)
  );
  FringeFF regs_48 ( // @[RegFile.scala 66:20:@38301.4]
    .clock(regs_48_clock),
    .reset(regs_48_reset),
    .io_in(regs_48_io_in),
    .io_reset(regs_48_io_reset),
    .io_out(regs_48_io_out),
    .io_enable(regs_48_io_enable)
  );
  FringeFF regs_49 ( // @[RegFile.scala 66:20:@38315.4]
    .clock(regs_49_clock),
    .reset(regs_49_reset),
    .io_in(regs_49_io_in),
    .io_reset(regs_49_io_reset),
    .io_out(regs_49_io_out),
    .io_enable(regs_49_io_enable)
  );
  FringeFF regs_50 ( // @[RegFile.scala 66:20:@38329.4]
    .clock(regs_50_clock),
    .reset(regs_50_reset),
    .io_in(regs_50_io_in),
    .io_reset(regs_50_io_reset),
    .io_out(regs_50_io_out),
    .io_enable(regs_50_io_enable)
  );
  FringeFF regs_51 ( // @[RegFile.scala 66:20:@38343.4]
    .clock(regs_51_clock),
    .reset(regs_51_reset),
    .io_in(regs_51_io_in),
    .io_reset(regs_51_io_reset),
    .io_out(regs_51_io_out),
    .io_enable(regs_51_io_enable)
  );
  FringeFF regs_52 ( // @[RegFile.scala 66:20:@38357.4]
    .clock(regs_52_clock),
    .reset(regs_52_reset),
    .io_in(regs_52_io_in),
    .io_reset(regs_52_io_reset),
    .io_out(regs_52_io_out),
    .io_enable(regs_52_io_enable)
  );
  FringeFF regs_53 ( // @[RegFile.scala 66:20:@38371.4]
    .clock(regs_53_clock),
    .reset(regs_53_reset),
    .io_in(regs_53_io_in),
    .io_reset(regs_53_io_reset),
    .io_out(regs_53_io_out),
    .io_enable(regs_53_io_enable)
  );
  FringeFF regs_54 ( // @[RegFile.scala 66:20:@38385.4]
    .clock(regs_54_clock),
    .reset(regs_54_reset),
    .io_in(regs_54_io_in),
    .io_reset(regs_54_io_reset),
    .io_out(regs_54_io_out),
    .io_enable(regs_54_io_enable)
  );
  FringeFF regs_55 ( // @[RegFile.scala 66:20:@38399.4]
    .clock(regs_55_clock),
    .reset(regs_55_reset),
    .io_in(regs_55_io_in),
    .io_reset(regs_55_io_reset),
    .io_out(regs_55_io_out),
    .io_enable(regs_55_io_enable)
  );
  FringeFF regs_56 ( // @[RegFile.scala 66:20:@38413.4]
    .clock(regs_56_clock),
    .reset(regs_56_reset),
    .io_in(regs_56_io_in),
    .io_reset(regs_56_io_reset),
    .io_out(regs_56_io_out),
    .io_enable(regs_56_io_enable)
  );
  FringeFF regs_57 ( // @[RegFile.scala 66:20:@38427.4]
    .clock(regs_57_clock),
    .reset(regs_57_reset),
    .io_in(regs_57_io_in),
    .io_reset(regs_57_io_reset),
    .io_out(regs_57_io_out),
    .io_enable(regs_57_io_enable)
  );
  FringeFF regs_58 ( // @[RegFile.scala 66:20:@38441.4]
    .clock(regs_58_clock),
    .reset(regs_58_reset),
    .io_in(regs_58_io_in),
    .io_reset(regs_58_io_reset),
    .io_out(regs_58_io_out),
    .io_enable(regs_58_io_enable)
  );
  FringeFF regs_59 ( // @[RegFile.scala 66:20:@38455.4]
    .clock(regs_59_clock),
    .reset(regs_59_reset),
    .io_in(regs_59_io_in),
    .io_reset(regs_59_io_reset),
    .io_out(regs_59_io_out),
    .io_enable(regs_59_io_enable)
  );
  FringeFF regs_60 ( // @[RegFile.scala 66:20:@38469.4]
    .clock(regs_60_clock),
    .reset(regs_60_reset),
    .io_in(regs_60_io_in),
    .io_reset(regs_60_io_reset),
    .io_out(regs_60_io_out),
    .io_enable(regs_60_io_enable)
  );
  FringeFF regs_61 ( // @[RegFile.scala 66:20:@38483.4]
    .clock(regs_61_clock),
    .reset(regs_61_reset),
    .io_in(regs_61_io_in),
    .io_reset(regs_61_io_reset),
    .io_out(regs_61_io_out),
    .io_enable(regs_61_io_enable)
  );
  FringeFF regs_62 ( // @[RegFile.scala 66:20:@38497.4]
    .clock(regs_62_clock),
    .reset(regs_62_reset),
    .io_in(regs_62_io_in),
    .io_reset(regs_62_io_reset),
    .io_out(regs_62_io_out),
    .io_enable(regs_62_io_enable)
  );
  FringeFF regs_63 ( // @[RegFile.scala 66:20:@38511.4]
    .clock(regs_63_clock),
    .reset(regs_63_reset),
    .io_in(regs_63_io_in),
    .io_reset(regs_63_io_reset),
    .io_out(regs_63_io_out),
    .io_enable(regs_63_io_enable)
  );
  FringeFF regs_64 ( // @[RegFile.scala 66:20:@38525.4]
    .clock(regs_64_clock),
    .reset(regs_64_reset),
    .io_in(regs_64_io_in),
    .io_reset(regs_64_io_reset),
    .io_out(regs_64_io_out),
    .io_enable(regs_64_io_enable)
  );
  FringeFF regs_65 ( // @[RegFile.scala 66:20:@38539.4]
    .clock(regs_65_clock),
    .reset(regs_65_reset),
    .io_in(regs_65_io_in),
    .io_reset(regs_65_io_reset),
    .io_out(regs_65_io_out),
    .io_enable(regs_65_io_enable)
  );
  FringeFF regs_66 ( // @[RegFile.scala 66:20:@38553.4]
    .clock(regs_66_clock),
    .reset(regs_66_reset),
    .io_in(regs_66_io_in),
    .io_reset(regs_66_io_reset),
    .io_out(regs_66_io_out),
    .io_enable(regs_66_io_enable)
  );
  FringeFF regs_67 ( // @[RegFile.scala 66:20:@38567.4]
    .clock(regs_67_clock),
    .reset(regs_67_reset),
    .io_in(regs_67_io_in),
    .io_reset(regs_67_io_reset),
    .io_out(regs_67_io_out),
    .io_enable(regs_67_io_enable)
  );
  FringeFF regs_68 ( // @[RegFile.scala 66:20:@38581.4]
    .clock(regs_68_clock),
    .reset(regs_68_reset),
    .io_in(regs_68_io_in),
    .io_reset(regs_68_io_reset),
    .io_out(regs_68_io_out),
    .io_enable(regs_68_io_enable)
  );
  FringeFF regs_69 ( // @[RegFile.scala 66:20:@38595.4]
    .clock(regs_69_clock),
    .reset(regs_69_reset),
    .io_in(regs_69_io_in),
    .io_reset(regs_69_io_reset),
    .io_out(regs_69_io_out),
    .io_enable(regs_69_io_enable)
  );
  FringeFF regs_70 ( // @[RegFile.scala 66:20:@38609.4]
    .clock(regs_70_clock),
    .reset(regs_70_reset),
    .io_in(regs_70_io_in),
    .io_reset(regs_70_io_reset),
    .io_out(regs_70_io_out),
    .io_enable(regs_70_io_enable)
  );
  FringeFF regs_71 ( // @[RegFile.scala 66:20:@38623.4]
    .clock(regs_71_clock),
    .reset(regs_71_reset),
    .io_in(regs_71_io_in),
    .io_reset(regs_71_io_reset),
    .io_out(regs_71_io_out),
    .io_enable(regs_71_io_enable)
  );
  FringeFF regs_72 ( // @[RegFile.scala 66:20:@38637.4]
    .clock(regs_72_clock),
    .reset(regs_72_reset),
    .io_in(regs_72_io_in),
    .io_reset(regs_72_io_reset),
    .io_out(regs_72_io_out),
    .io_enable(regs_72_io_enable)
  );
  FringeFF regs_73 ( // @[RegFile.scala 66:20:@38651.4]
    .clock(regs_73_clock),
    .reset(regs_73_reset),
    .io_in(regs_73_io_in),
    .io_reset(regs_73_io_reset),
    .io_out(regs_73_io_out),
    .io_enable(regs_73_io_enable)
  );
  FringeFF regs_74 ( // @[RegFile.scala 66:20:@38665.4]
    .clock(regs_74_clock),
    .reset(regs_74_reset),
    .io_in(regs_74_io_in),
    .io_reset(regs_74_io_reset),
    .io_out(regs_74_io_out),
    .io_enable(regs_74_io_enable)
  );
  FringeFF regs_75 ( // @[RegFile.scala 66:20:@38679.4]
    .clock(regs_75_clock),
    .reset(regs_75_reset),
    .io_in(regs_75_io_in),
    .io_reset(regs_75_io_reset),
    .io_out(regs_75_io_out),
    .io_enable(regs_75_io_enable)
  );
  FringeFF regs_76 ( // @[RegFile.scala 66:20:@38693.4]
    .clock(regs_76_clock),
    .reset(regs_76_reset),
    .io_in(regs_76_io_in),
    .io_reset(regs_76_io_reset),
    .io_out(regs_76_io_out),
    .io_enable(regs_76_io_enable)
  );
  FringeFF regs_77 ( // @[RegFile.scala 66:20:@38707.4]
    .clock(regs_77_clock),
    .reset(regs_77_reset),
    .io_in(regs_77_io_in),
    .io_reset(regs_77_io_reset),
    .io_out(regs_77_io_out),
    .io_enable(regs_77_io_enable)
  );
  FringeFF regs_78 ( // @[RegFile.scala 66:20:@38721.4]
    .clock(regs_78_clock),
    .reset(regs_78_reset),
    .io_in(regs_78_io_in),
    .io_reset(regs_78_io_reset),
    .io_out(regs_78_io_out),
    .io_enable(regs_78_io_enable)
  );
  FringeFF regs_79 ( // @[RegFile.scala 66:20:@38735.4]
    .clock(regs_79_clock),
    .reset(regs_79_reset),
    .io_in(regs_79_io_in),
    .io_reset(regs_79_io_reset),
    .io_out(regs_79_io_out),
    .io_enable(regs_79_io_enable)
  );
  FringeFF regs_80 ( // @[RegFile.scala 66:20:@38749.4]
    .clock(regs_80_clock),
    .reset(regs_80_reset),
    .io_in(regs_80_io_in),
    .io_reset(regs_80_io_reset),
    .io_out(regs_80_io_out),
    .io_enable(regs_80_io_enable)
  );
  FringeFF regs_81 ( // @[RegFile.scala 66:20:@38763.4]
    .clock(regs_81_clock),
    .reset(regs_81_reset),
    .io_in(regs_81_io_in),
    .io_reset(regs_81_io_reset),
    .io_out(regs_81_io_out),
    .io_enable(regs_81_io_enable)
  );
  FringeFF regs_82 ( // @[RegFile.scala 66:20:@38777.4]
    .clock(regs_82_clock),
    .reset(regs_82_reset),
    .io_in(regs_82_io_in),
    .io_reset(regs_82_io_reset),
    .io_out(regs_82_io_out),
    .io_enable(regs_82_io_enable)
  );
  FringeFF regs_83 ( // @[RegFile.scala 66:20:@38791.4]
    .clock(regs_83_clock),
    .reset(regs_83_reset),
    .io_in(regs_83_io_in),
    .io_reset(regs_83_io_reset),
    .io_out(regs_83_io_out),
    .io_enable(regs_83_io_enable)
  );
  FringeFF regs_84 ( // @[RegFile.scala 66:20:@38805.4]
    .clock(regs_84_clock),
    .reset(regs_84_reset),
    .io_in(regs_84_io_in),
    .io_reset(regs_84_io_reset),
    .io_out(regs_84_io_out),
    .io_enable(regs_84_io_enable)
  );
  FringeFF regs_85 ( // @[RegFile.scala 66:20:@38819.4]
    .clock(regs_85_clock),
    .reset(regs_85_reset),
    .io_in(regs_85_io_in),
    .io_reset(regs_85_io_reset),
    .io_out(regs_85_io_out),
    .io_enable(regs_85_io_enable)
  );
  FringeFF regs_86 ( // @[RegFile.scala 66:20:@38833.4]
    .clock(regs_86_clock),
    .reset(regs_86_reset),
    .io_in(regs_86_io_in),
    .io_reset(regs_86_io_reset),
    .io_out(regs_86_io_out),
    .io_enable(regs_86_io_enable)
  );
  FringeFF regs_87 ( // @[RegFile.scala 66:20:@38847.4]
    .clock(regs_87_clock),
    .reset(regs_87_reset),
    .io_in(regs_87_io_in),
    .io_reset(regs_87_io_reset),
    .io_out(regs_87_io_out),
    .io_enable(regs_87_io_enable)
  );
  FringeFF regs_88 ( // @[RegFile.scala 66:20:@38861.4]
    .clock(regs_88_clock),
    .reset(regs_88_reset),
    .io_in(regs_88_io_in),
    .io_reset(regs_88_io_reset),
    .io_out(regs_88_io_out),
    .io_enable(regs_88_io_enable)
  );
  FringeFF regs_89 ( // @[RegFile.scala 66:20:@38875.4]
    .clock(regs_89_clock),
    .reset(regs_89_reset),
    .io_in(regs_89_io_in),
    .io_reset(regs_89_io_reset),
    .io_out(regs_89_io_out),
    .io_enable(regs_89_io_enable)
  );
  FringeFF regs_90 ( // @[RegFile.scala 66:20:@38889.4]
    .clock(regs_90_clock),
    .reset(regs_90_reset),
    .io_in(regs_90_io_in),
    .io_reset(regs_90_io_reset),
    .io_out(regs_90_io_out),
    .io_enable(regs_90_io_enable)
  );
  FringeFF regs_91 ( // @[RegFile.scala 66:20:@38903.4]
    .clock(regs_91_clock),
    .reset(regs_91_reset),
    .io_in(regs_91_io_in),
    .io_reset(regs_91_io_reset),
    .io_out(regs_91_io_out),
    .io_enable(regs_91_io_enable)
  );
  FringeFF regs_92 ( // @[RegFile.scala 66:20:@38917.4]
    .clock(regs_92_clock),
    .reset(regs_92_reset),
    .io_in(regs_92_io_in),
    .io_reset(regs_92_io_reset),
    .io_out(regs_92_io_out),
    .io_enable(regs_92_io_enable)
  );
  FringeFF regs_93 ( // @[RegFile.scala 66:20:@38931.4]
    .clock(regs_93_clock),
    .reset(regs_93_reset),
    .io_in(regs_93_io_in),
    .io_reset(regs_93_io_reset),
    .io_out(regs_93_io_out),
    .io_enable(regs_93_io_enable)
  );
  FringeFF regs_94 ( // @[RegFile.scala 66:20:@38945.4]
    .clock(regs_94_clock),
    .reset(regs_94_reset),
    .io_in(regs_94_io_in),
    .io_reset(regs_94_io_reset),
    .io_out(regs_94_io_out),
    .io_enable(regs_94_io_enable)
  );
  FringeFF regs_95 ( // @[RegFile.scala 66:20:@38959.4]
    .clock(regs_95_clock),
    .reset(regs_95_reset),
    .io_in(regs_95_io_in),
    .io_reset(regs_95_io_reset),
    .io_out(regs_95_io_out),
    .io_enable(regs_95_io_enable)
  );
  FringeFF regs_96 ( // @[RegFile.scala 66:20:@38973.4]
    .clock(regs_96_clock),
    .reset(regs_96_reset),
    .io_in(regs_96_io_in),
    .io_reset(regs_96_io_reset),
    .io_out(regs_96_io_out),
    .io_enable(regs_96_io_enable)
  );
  FringeFF regs_97 ( // @[RegFile.scala 66:20:@38987.4]
    .clock(regs_97_clock),
    .reset(regs_97_reset),
    .io_in(regs_97_io_in),
    .io_reset(regs_97_io_reset),
    .io_out(regs_97_io_out),
    .io_enable(regs_97_io_enable)
  );
  FringeFF regs_98 ( // @[RegFile.scala 66:20:@39001.4]
    .clock(regs_98_clock),
    .reset(regs_98_reset),
    .io_in(regs_98_io_in),
    .io_reset(regs_98_io_reset),
    .io_out(regs_98_io_out),
    .io_enable(regs_98_io_enable)
  );
  FringeFF regs_99 ( // @[RegFile.scala 66:20:@39015.4]
    .clock(regs_99_clock),
    .reset(regs_99_reset),
    .io_in(regs_99_io_in),
    .io_reset(regs_99_io_reset),
    .io_out(regs_99_io_out),
    .io_enable(regs_99_io_enable)
  );
  FringeFF regs_100 ( // @[RegFile.scala 66:20:@39029.4]
    .clock(regs_100_clock),
    .reset(regs_100_reset),
    .io_in(regs_100_io_in),
    .io_reset(regs_100_io_reset),
    .io_out(regs_100_io_out),
    .io_enable(regs_100_io_enable)
  );
  FringeFF regs_101 ( // @[RegFile.scala 66:20:@39043.4]
    .clock(regs_101_clock),
    .reset(regs_101_reset),
    .io_in(regs_101_io_in),
    .io_reset(regs_101_io_reset),
    .io_out(regs_101_io_out),
    .io_enable(regs_101_io_enable)
  );
  FringeFF regs_102 ( // @[RegFile.scala 66:20:@39057.4]
    .clock(regs_102_clock),
    .reset(regs_102_reset),
    .io_in(regs_102_io_in),
    .io_reset(regs_102_io_reset),
    .io_out(regs_102_io_out),
    .io_enable(regs_102_io_enable)
  );
  FringeFF regs_103 ( // @[RegFile.scala 66:20:@39071.4]
    .clock(regs_103_clock),
    .reset(regs_103_reset),
    .io_in(regs_103_io_in),
    .io_reset(regs_103_io_reset),
    .io_out(regs_103_io_out),
    .io_enable(regs_103_io_enable)
  );
  FringeFF regs_104 ( // @[RegFile.scala 66:20:@39085.4]
    .clock(regs_104_clock),
    .reset(regs_104_reset),
    .io_in(regs_104_io_in),
    .io_reset(regs_104_io_reset),
    .io_out(regs_104_io_out),
    .io_enable(regs_104_io_enable)
  );
  FringeFF regs_105 ( // @[RegFile.scala 66:20:@39099.4]
    .clock(regs_105_clock),
    .reset(regs_105_reset),
    .io_in(regs_105_io_in),
    .io_reset(regs_105_io_reset),
    .io_out(regs_105_io_out),
    .io_enable(regs_105_io_enable)
  );
  FringeFF regs_106 ( // @[RegFile.scala 66:20:@39113.4]
    .clock(regs_106_clock),
    .reset(regs_106_reset),
    .io_in(regs_106_io_in),
    .io_reset(regs_106_io_reset),
    .io_out(regs_106_io_out),
    .io_enable(regs_106_io_enable)
  );
  FringeFF regs_107 ( // @[RegFile.scala 66:20:@39127.4]
    .clock(regs_107_clock),
    .reset(regs_107_reset),
    .io_in(regs_107_io_in),
    .io_reset(regs_107_io_reset),
    .io_out(regs_107_io_out),
    .io_enable(regs_107_io_enable)
  );
  FringeFF regs_108 ( // @[RegFile.scala 66:20:@39141.4]
    .clock(regs_108_clock),
    .reset(regs_108_reset),
    .io_in(regs_108_io_in),
    .io_reset(regs_108_io_reset),
    .io_out(regs_108_io_out),
    .io_enable(regs_108_io_enable)
  );
  FringeFF regs_109 ( // @[RegFile.scala 66:20:@39155.4]
    .clock(regs_109_clock),
    .reset(regs_109_reset),
    .io_in(regs_109_io_in),
    .io_reset(regs_109_io_reset),
    .io_out(regs_109_io_out),
    .io_enable(regs_109_io_enable)
  );
  FringeFF regs_110 ( // @[RegFile.scala 66:20:@39169.4]
    .clock(regs_110_clock),
    .reset(regs_110_reset),
    .io_in(regs_110_io_in),
    .io_reset(regs_110_io_reset),
    .io_out(regs_110_io_out),
    .io_enable(regs_110_io_enable)
  );
  FringeFF regs_111 ( // @[RegFile.scala 66:20:@39183.4]
    .clock(regs_111_clock),
    .reset(regs_111_reset),
    .io_in(regs_111_io_in),
    .io_reset(regs_111_io_reset),
    .io_out(regs_111_io_out),
    .io_enable(regs_111_io_enable)
  );
  FringeFF regs_112 ( // @[RegFile.scala 66:20:@39197.4]
    .clock(regs_112_clock),
    .reset(regs_112_reset),
    .io_in(regs_112_io_in),
    .io_reset(regs_112_io_reset),
    .io_out(regs_112_io_out),
    .io_enable(regs_112_io_enable)
  );
  FringeFF regs_113 ( // @[RegFile.scala 66:20:@39211.4]
    .clock(regs_113_clock),
    .reset(regs_113_reset),
    .io_in(regs_113_io_in),
    .io_reset(regs_113_io_reset),
    .io_out(regs_113_io_out),
    .io_enable(regs_113_io_enable)
  );
  FringeFF regs_114 ( // @[RegFile.scala 66:20:@39225.4]
    .clock(regs_114_clock),
    .reset(regs_114_reset),
    .io_in(regs_114_io_in),
    .io_reset(regs_114_io_reset),
    .io_out(regs_114_io_out),
    .io_enable(regs_114_io_enable)
  );
  FringeFF regs_115 ( // @[RegFile.scala 66:20:@39239.4]
    .clock(regs_115_clock),
    .reset(regs_115_reset),
    .io_in(regs_115_io_in),
    .io_reset(regs_115_io_reset),
    .io_out(regs_115_io_out),
    .io_enable(regs_115_io_enable)
  );
  FringeFF regs_116 ( // @[RegFile.scala 66:20:@39253.4]
    .clock(regs_116_clock),
    .reset(regs_116_reset),
    .io_in(regs_116_io_in),
    .io_reset(regs_116_io_reset),
    .io_out(regs_116_io_out),
    .io_enable(regs_116_io_enable)
  );
  FringeFF regs_117 ( // @[RegFile.scala 66:20:@39267.4]
    .clock(regs_117_clock),
    .reset(regs_117_reset),
    .io_in(regs_117_io_in),
    .io_reset(regs_117_io_reset),
    .io_out(regs_117_io_out),
    .io_enable(regs_117_io_enable)
  );
  FringeFF regs_118 ( // @[RegFile.scala 66:20:@39281.4]
    .clock(regs_118_clock),
    .reset(regs_118_reset),
    .io_in(regs_118_io_in),
    .io_reset(regs_118_io_reset),
    .io_out(regs_118_io_out),
    .io_enable(regs_118_io_enable)
  );
  FringeFF regs_119 ( // @[RegFile.scala 66:20:@39295.4]
    .clock(regs_119_clock),
    .reset(regs_119_reset),
    .io_in(regs_119_io_in),
    .io_reset(regs_119_io_reset),
    .io_out(regs_119_io_out),
    .io_enable(regs_119_io_enable)
  );
  FringeFF regs_120 ( // @[RegFile.scala 66:20:@39309.4]
    .clock(regs_120_clock),
    .reset(regs_120_reset),
    .io_in(regs_120_io_in),
    .io_reset(regs_120_io_reset),
    .io_out(regs_120_io_out),
    .io_enable(regs_120_io_enable)
  );
  FringeFF regs_121 ( // @[RegFile.scala 66:20:@39323.4]
    .clock(regs_121_clock),
    .reset(regs_121_reset),
    .io_in(regs_121_io_in),
    .io_reset(regs_121_io_reset),
    .io_out(regs_121_io_out),
    .io_enable(regs_121_io_enable)
  );
  FringeFF regs_122 ( // @[RegFile.scala 66:20:@39337.4]
    .clock(regs_122_clock),
    .reset(regs_122_reset),
    .io_in(regs_122_io_in),
    .io_reset(regs_122_io_reset),
    .io_out(regs_122_io_out),
    .io_enable(regs_122_io_enable)
  );
  FringeFF regs_123 ( // @[RegFile.scala 66:20:@39351.4]
    .clock(regs_123_clock),
    .reset(regs_123_reset),
    .io_in(regs_123_io_in),
    .io_reset(regs_123_io_reset),
    .io_out(regs_123_io_out),
    .io_enable(regs_123_io_enable)
  );
  FringeFF regs_124 ( // @[RegFile.scala 66:20:@39365.4]
    .clock(regs_124_clock),
    .reset(regs_124_reset),
    .io_in(regs_124_io_in),
    .io_reset(regs_124_io_reset),
    .io_out(regs_124_io_out),
    .io_enable(regs_124_io_enable)
  );
  FringeFF regs_125 ( // @[RegFile.scala 66:20:@39379.4]
    .clock(regs_125_clock),
    .reset(regs_125_reset),
    .io_in(regs_125_io_in),
    .io_reset(regs_125_io_reset),
    .io_out(regs_125_io_out),
    .io_enable(regs_125_io_enable)
  );
  FringeFF regs_126 ( // @[RegFile.scala 66:20:@39393.4]
    .clock(regs_126_clock),
    .reset(regs_126_reset),
    .io_in(regs_126_io_in),
    .io_reset(regs_126_io_reset),
    .io_out(regs_126_io_out),
    .io_enable(regs_126_io_enable)
  );
  FringeFF regs_127 ( // @[RegFile.scala 66:20:@39407.4]
    .clock(regs_127_clock),
    .reset(regs_127_reset),
    .io_in(regs_127_io_in),
    .io_reset(regs_127_io_reset),
    .io_out(regs_127_io_out),
    .io_enable(regs_127_io_enable)
  );
  FringeFF regs_128 ( // @[RegFile.scala 66:20:@39421.4]
    .clock(regs_128_clock),
    .reset(regs_128_reset),
    .io_in(regs_128_io_in),
    .io_reset(regs_128_io_reset),
    .io_out(regs_128_io_out),
    .io_enable(regs_128_io_enable)
  );
  FringeFF regs_129 ( // @[RegFile.scala 66:20:@39435.4]
    .clock(regs_129_clock),
    .reset(regs_129_reset),
    .io_in(regs_129_io_in),
    .io_reset(regs_129_io_reset),
    .io_out(regs_129_io_out),
    .io_enable(regs_129_io_enable)
  );
  FringeFF regs_130 ( // @[RegFile.scala 66:20:@39449.4]
    .clock(regs_130_clock),
    .reset(regs_130_reset),
    .io_in(regs_130_io_in),
    .io_reset(regs_130_io_reset),
    .io_out(regs_130_io_out),
    .io_enable(regs_130_io_enable)
  );
  FringeFF regs_131 ( // @[RegFile.scala 66:20:@39463.4]
    .clock(regs_131_clock),
    .reset(regs_131_reset),
    .io_in(regs_131_io_in),
    .io_reset(regs_131_io_reset),
    .io_out(regs_131_io_out),
    .io_enable(regs_131_io_enable)
  );
  FringeFF regs_132 ( // @[RegFile.scala 66:20:@39477.4]
    .clock(regs_132_clock),
    .reset(regs_132_reset),
    .io_in(regs_132_io_in),
    .io_reset(regs_132_io_reset),
    .io_out(regs_132_io_out),
    .io_enable(regs_132_io_enable)
  );
  FringeFF regs_133 ( // @[RegFile.scala 66:20:@39491.4]
    .clock(regs_133_clock),
    .reset(regs_133_reset),
    .io_in(regs_133_io_in),
    .io_reset(regs_133_io_reset),
    .io_out(regs_133_io_out),
    .io_enable(regs_133_io_enable)
  );
  FringeFF regs_134 ( // @[RegFile.scala 66:20:@39505.4]
    .clock(regs_134_clock),
    .reset(regs_134_reset),
    .io_in(regs_134_io_in),
    .io_reset(regs_134_io_reset),
    .io_out(regs_134_io_out),
    .io_enable(regs_134_io_enable)
  );
  FringeFF regs_135 ( // @[RegFile.scala 66:20:@39519.4]
    .clock(regs_135_clock),
    .reset(regs_135_reset),
    .io_in(regs_135_io_in),
    .io_reset(regs_135_io_reset),
    .io_out(regs_135_io_out),
    .io_enable(regs_135_io_enable)
  );
  FringeFF regs_136 ( // @[RegFile.scala 66:20:@39533.4]
    .clock(regs_136_clock),
    .reset(regs_136_reset),
    .io_in(regs_136_io_in),
    .io_reset(regs_136_io_reset),
    .io_out(regs_136_io_out),
    .io_enable(regs_136_io_enable)
  );
  FringeFF regs_137 ( // @[RegFile.scala 66:20:@39547.4]
    .clock(regs_137_clock),
    .reset(regs_137_reset),
    .io_in(regs_137_io_in),
    .io_reset(regs_137_io_reset),
    .io_out(regs_137_io_out),
    .io_enable(regs_137_io_enable)
  );
  FringeFF regs_138 ( // @[RegFile.scala 66:20:@39561.4]
    .clock(regs_138_clock),
    .reset(regs_138_reset),
    .io_in(regs_138_io_in),
    .io_reset(regs_138_io_reset),
    .io_out(regs_138_io_out),
    .io_enable(regs_138_io_enable)
  );
  FringeFF regs_139 ( // @[RegFile.scala 66:20:@39575.4]
    .clock(regs_139_clock),
    .reset(regs_139_reset),
    .io_in(regs_139_io_in),
    .io_reset(regs_139_io_reset),
    .io_out(regs_139_io_out),
    .io_enable(regs_139_io_enable)
  );
  FringeFF regs_140 ( // @[RegFile.scala 66:20:@39589.4]
    .clock(regs_140_clock),
    .reset(regs_140_reset),
    .io_in(regs_140_io_in),
    .io_reset(regs_140_io_reset),
    .io_out(regs_140_io_out),
    .io_enable(regs_140_io_enable)
  );
  FringeFF regs_141 ( // @[RegFile.scala 66:20:@39603.4]
    .clock(regs_141_clock),
    .reset(regs_141_reset),
    .io_in(regs_141_io_in),
    .io_reset(regs_141_io_reset),
    .io_out(regs_141_io_out),
    .io_enable(regs_141_io_enable)
  );
  FringeFF regs_142 ( // @[RegFile.scala 66:20:@39617.4]
    .clock(regs_142_clock),
    .reset(regs_142_reset),
    .io_in(regs_142_io_in),
    .io_reset(regs_142_io_reset),
    .io_out(regs_142_io_out),
    .io_enable(regs_142_io_enable)
  );
  FringeFF regs_143 ( // @[RegFile.scala 66:20:@39631.4]
    .clock(regs_143_clock),
    .reset(regs_143_reset),
    .io_in(regs_143_io_in),
    .io_reset(regs_143_io_reset),
    .io_out(regs_143_io_out),
    .io_enable(regs_143_io_enable)
  );
  FringeFF regs_144 ( // @[RegFile.scala 66:20:@39645.4]
    .clock(regs_144_clock),
    .reset(regs_144_reset),
    .io_in(regs_144_io_in),
    .io_reset(regs_144_io_reset),
    .io_out(regs_144_io_out),
    .io_enable(regs_144_io_enable)
  );
  FringeFF regs_145 ( // @[RegFile.scala 66:20:@39659.4]
    .clock(regs_145_clock),
    .reset(regs_145_reset),
    .io_in(regs_145_io_in),
    .io_reset(regs_145_io_reset),
    .io_out(regs_145_io_out),
    .io_enable(regs_145_io_enable)
  );
  FringeFF regs_146 ( // @[RegFile.scala 66:20:@39673.4]
    .clock(regs_146_clock),
    .reset(regs_146_reset),
    .io_in(regs_146_io_in),
    .io_reset(regs_146_io_reset),
    .io_out(regs_146_io_out),
    .io_enable(regs_146_io_enable)
  );
  FringeFF regs_147 ( // @[RegFile.scala 66:20:@39687.4]
    .clock(regs_147_clock),
    .reset(regs_147_reset),
    .io_in(regs_147_io_in),
    .io_reset(regs_147_io_reset),
    .io_out(regs_147_io_out),
    .io_enable(regs_147_io_enable)
  );
  FringeFF regs_148 ( // @[RegFile.scala 66:20:@39701.4]
    .clock(regs_148_clock),
    .reset(regs_148_reset),
    .io_in(regs_148_io_in),
    .io_reset(regs_148_io_reset),
    .io_out(regs_148_io_out),
    .io_enable(regs_148_io_enable)
  );
  FringeFF regs_149 ( // @[RegFile.scala 66:20:@39715.4]
    .clock(regs_149_clock),
    .reset(regs_149_reset),
    .io_in(regs_149_io_in),
    .io_reset(regs_149_io_reset),
    .io_out(regs_149_io_out),
    .io_enable(regs_149_io_enable)
  );
  FringeFF regs_150 ( // @[RegFile.scala 66:20:@39729.4]
    .clock(regs_150_clock),
    .reset(regs_150_reset),
    .io_in(regs_150_io_in),
    .io_reset(regs_150_io_reset),
    .io_out(regs_150_io_out),
    .io_enable(regs_150_io_enable)
  );
  FringeFF regs_151 ( // @[RegFile.scala 66:20:@39743.4]
    .clock(regs_151_clock),
    .reset(regs_151_reset),
    .io_in(regs_151_io_in),
    .io_reset(regs_151_io_reset),
    .io_out(regs_151_io_out),
    .io_enable(regs_151_io_enable)
  );
  FringeFF regs_152 ( // @[RegFile.scala 66:20:@39757.4]
    .clock(regs_152_clock),
    .reset(regs_152_reset),
    .io_in(regs_152_io_in),
    .io_reset(regs_152_io_reset),
    .io_out(regs_152_io_out),
    .io_enable(regs_152_io_enable)
  );
  FringeFF regs_153 ( // @[RegFile.scala 66:20:@39771.4]
    .clock(regs_153_clock),
    .reset(regs_153_reset),
    .io_in(regs_153_io_in),
    .io_reset(regs_153_io_reset),
    .io_out(regs_153_io_out),
    .io_enable(regs_153_io_enable)
  );
  FringeFF regs_154 ( // @[RegFile.scala 66:20:@39785.4]
    .clock(regs_154_clock),
    .reset(regs_154_reset),
    .io_in(regs_154_io_in),
    .io_reset(regs_154_io_reset),
    .io_out(regs_154_io_out),
    .io_enable(regs_154_io_enable)
  );
  FringeFF regs_155 ( // @[RegFile.scala 66:20:@39799.4]
    .clock(regs_155_clock),
    .reset(regs_155_reset),
    .io_in(regs_155_io_in),
    .io_reset(regs_155_io_reset),
    .io_out(regs_155_io_out),
    .io_enable(regs_155_io_enable)
  );
  FringeFF regs_156 ( // @[RegFile.scala 66:20:@39813.4]
    .clock(regs_156_clock),
    .reset(regs_156_reset),
    .io_in(regs_156_io_in),
    .io_reset(regs_156_io_reset),
    .io_out(regs_156_io_out),
    .io_enable(regs_156_io_enable)
  );
  FringeFF regs_157 ( // @[RegFile.scala 66:20:@39827.4]
    .clock(regs_157_clock),
    .reset(regs_157_reset),
    .io_in(regs_157_io_in),
    .io_reset(regs_157_io_reset),
    .io_out(regs_157_io_out),
    .io_enable(regs_157_io_enable)
  );
  FringeFF regs_158 ( // @[RegFile.scala 66:20:@39841.4]
    .clock(regs_158_clock),
    .reset(regs_158_reset),
    .io_in(regs_158_io_in),
    .io_reset(regs_158_io_reset),
    .io_out(regs_158_io_out),
    .io_enable(regs_158_io_enable)
  );
  FringeFF regs_159 ( // @[RegFile.scala 66:20:@39855.4]
    .clock(regs_159_clock),
    .reset(regs_159_reset),
    .io_in(regs_159_io_in),
    .io_reset(regs_159_io_reset),
    .io_out(regs_159_io_out),
    .io_enable(regs_159_io_enable)
  );
  FringeFF regs_160 ( // @[RegFile.scala 66:20:@39869.4]
    .clock(regs_160_clock),
    .reset(regs_160_reset),
    .io_in(regs_160_io_in),
    .io_reset(regs_160_io_reset),
    .io_out(regs_160_io_out),
    .io_enable(regs_160_io_enable)
  );
  FringeFF regs_161 ( // @[RegFile.scala 66:20:@39883.4]
    .clock(regs_161_clock),
    .reset(regs_161_reset),
    .io_in(regs_161_io_in),
    .io_reset(regs_161_io_reset),
    .io_out(regs_161_io_out),
    .io_enable(regs_161_io_enable)
  );
  FringeFF regs_162 ( // @[RegFile.scala 66:20:@39897.4]
    .clock(regs_162_clock),
    .reset(regs_162_reset),
    .io_in(regs_162_io_in),
    .io_reset(regs_162_io_reset),
    .io_out(regs_162_io_out),
    .io_enable(regs_162_io_enable)
  );
  FringeFF regs_163 ( // @[RegFile.scala 66:20:@39911.4]
    .clock(regs_163_clock),
    .reset(regs_163_reset),
    .io_in(regs_163_io_in),
    .io_reset(regs_163_io_reset),
    .io_out(regs_163_io_out),
    .io_enable(regs_163_io_enable)
  );
  FringeFF regs_164 ( // @[RegFile.scala 66:20:@39925.4]
    .clock(regs_164_clock),
    .reset(regs_164_reset),
    .io_in(regs_164_io_in),
    .io_reset(regs_164_io_reset),
    .io_out(regs_164_io_out),
    .io_enable(regs_164_io_enable)
  );
  FringeFF regs_165 ( // @[RegFile.scala 66:20:@39939.4]
    .clock(regs_165_clock),
    .reset(regs_165_reset),
    .io_in(regs_165_io_in),
    .io_reset(regs_165_io_reset),
    .io_out(regs_165_io_out),
    .io_enable(regs_165_io_enable)
  );
  FringeFF regs_166 ( // @[RegFile.scala 66:20:@39953.4]
    .clock(regs_166_clock),
    .reset(regs_166_reset),
    .io_in(regs_166_io_in),
    .io_reset(regs_166_io_reset),
    .io_out(regs_166_io_out),
    .io_enable(regs_166_io_enable)
  );
  FringeFF regs_167 ( // @[RegFile.scala 66:20:@39967.4]
    .clock(regs_167_clock),
    .reset(regs_167_reset),
    .io_in(regs_167_io_in),
    .io_reset(regs_167_io_reset),
    .io_out(regs_167_io_out),
    .io_enable(regs_167_io_enable)
  );
  FringeFF regs_168 ( // @[RegFile.scala 66:20:@39981.4]
    .clock(regs_168_clock),
    .reset(regs_168_reset),
    .io_in(regs_168_io_in),
    .io_reset(regs_168_io_reset),
    .io_out(regs_168_io_out),
    .io_enable(regs_168_io_enable)
  );
  FringeFF regs_169 ( // @[RegFile.scala 66:20:@39995.4]
    .clock(regs_169_clock),
    .reset(regs_169_reset),
    .io_in(regs_169_io_in),
    .io_reset(regs_169_io_reset),
    .io_out(regs_169_io_out),
    .io_enable(regs_169_io_enable)
  );
  FringeFF regs_170 ( // @[RegFile.scala 66:20:@40009.4]
    .clock(regs_170_clock),
    .reset(regs_170_reset),
    .io_in(regs_170_io_in),
    .io_reset(regs_170_io_reset),
    .io_out(regs_170_io_out),
    .io_enable(regs_170_io_enable)
  );
  FringeFF regs_171 ( // @[RegFile.scala 66:20:@40023.4]
    .clock(regs_171_clock),
    .reset(regs_171_reset),
    .io_in(regs_171_io_in),
    .io_reset(regs_171_io_reset),
    .io_out(regs_171_io_out),
    .io_enable(regs_171_io_enable)
  );
  FringeFF regs_172 ( // @[RegFile.scala 66:20:@40037.4]
    .clock(regs_172_clock),
    .reset(regs_172_reset),
    .io_in(regs_172_io_in),
    .io_reset(regs_172_io_reset),
    .io_out(regs_172_io_out),
    .io_enable(regs_172_io_enable)
  );
  FringeFF regs_173 ( // @[RegFile.scala 66:20:@40051.4]
    .clock(regs_173_clock),
    .reset(regs_173_reset),
    .io_in(regs_173_io_in),
    .io_reset(regs_173_io_reset),
    .io_out(regs_173_io_out),
    .io_enable(regs_173_io_enable)
  );
  FringeFF regs_174 ( // @[RegFile.scala 66:20:@40065.4]
    .clock(regs_174_clock),
    .reset(regs_174_reset),
    .io_in(regs_174_io_in),
    .io_reset(regs_174_io_reset),
    .io_out(regs_174_io_out),
    .io_enable(regs_174_io_enable)
  );
  FringeFF regs_175 ( // @[RegFile.scala 66:20:@40079.4]
    .clock(regs_175_clock),
    .reset(regs_175_reset),
    .io_in(regs_175_io_in),
    .io_reset(regs_175_io_reset),
    .io_out(regs_175_io_out),
    .io_enable(regs_175_io_enable)
  );
  FringeFF regs_176 ( // @[RegFile.scala 66:20:@40093.4]
    .clock(regs_176_clock),
    .reset(regs_176_reset),
    .io_in(regs_176_io_in),
    .io_reset(regs_176_io_reset),
    .io_out(regs_176_io_out),
    .io_enable(regs_176_io_enable)
  );
  FringeFF regs_177 ( // @[RegFile.scala 66:20:@40107.4]
    .clock(regs_177_clock),
    .reset(regs_177_reset),
    .io_in(regs_177_io_in),
    .io_reset(regs_177_io_reset),
    .io_out(regs_177_io_out),
    .io_enable(regs_177_io_enable)
  );
  FringeFF regs_178 ( // @[RegFile.scala 66:20:@40121.4]
    .clock(regs_178_clock),
    .reset(regs_178_reset),
    .io_in(regs_178_io_in),
    .io_reset(regs_178_io_reset),
    .io_out(regs_178_io_out),
    .io_enable(regs_178_io_enable)
  );
  FringeFF regs_179 ( // @[RegFile.scala 66:20:@40135.4]
    .clock(regs_179_clock),
    .reset(regs_179_reset),
    .io_in(regs_179_io_in),
    .io_reset(regs_179_io_reset),
    .io_out(regs_179_io_out),
    .io_enable(regs_179_io_enable)
  );
  FringeFF regs_180 ( // @[RegFile.scala 66:20:@40149.4]
    .clock(regs_180_clock),
    .reset(regs_180_reset),
    .io_in(regs_180_io_in),
    .io_reset(regs_180_io_reset),
    .io_out(regs_180_io_out),
    .io_enable(regs_180_io_enable)
  );
  FringeFF regs_181 ( // @[RegFile.scala 66:20:@40163.4]
    .clock(regs_181_clock),
    .reset(regs_181_reset),
    .io_in(regs_181_io_in),
    .io_reset(regs_181_io_reset),
    .io_out(regs_181_io_out),
    .io_enable(regs_181_io_enable)
  );
  FringeFF regs_182 ( // @[RegFile.scala 66:20:@40177.4]
    .clock(regs_182_clock),
    .reset(regs_182_reset),
    .io_in(regs_182_io_in),
    .io_reset(regs_182_io_reset),
    .io_out(regs_182_io_out),
    .io_enable(regs_182_io_enable)
  );
  FringeFF regs_183 ( // @[RegFile.scala 66:20:@40191.4]
    .clock(regs_183_clock),
    .reset(regs_183_reset),
    .io_in(regs_183_io_in),
    .io_reset(regs_183_io_reset),
    .io_out(regs_183_io_out),
    .io_enable(regs_183_io_enable)
  );
  FringeFF regs_184 ( // @[RegFile.scala 66:20:@40205.4]
    .clock(regs_184_clock),
    .reset(regs_184_reset),
    .io_in(regs_184_io_in),
    .io_reset(regs_184_io_reset),
    .io_out(regs_184_io_out),
    .io_enable(regs_184_io_enable)
  );
  FringeFF regs_185 ( // @[RegFile.scala 66:20:@40219.4]
    .clock(regs_185_clock),
    .reset(regs_185_reset),
    .io_in(regs_185_io_in),
    .io_reset(regs_185_io_reset),
    .io_out(regs_185_io_out),
    .io_enable(regs_185_io_enable)
  );
  FringeFF regs_186 ( // @[RegFile.scala 66:20:@40233.4]
    .clock(regs_186_clock),
    .reset(regs_186_reset),
    .io_in(regs_186_io_in),
    .io_reset(regs_186_io_reset),
    .io_out(regs_186_io_out),
    .io_enable(regs_186_io_enable)
  );
  FringeFF regs_187 ( // @[RegFile.scala 66:20:@40247.4]
    .clock(regs_187_clock),
    .reset(regs_187_reset),
    .io_in(regs_187_io_in),
    .io_reset(regs_187_io_reset),
    .io_out(regs_187_io_out),
    .io_enable(regs_187_io_enable)
  );
  FringeFF regs_188 ( // @[RegFile.scala 66:20:@40261.4]
    .clock(regs_188_clock),
    .reset(regs_188_reset),
    .io_in(regs_188_io_in),
    .io_reset(regs_188_io_reset),
    .io_out(regs_188_io_out),
    .io_enable(regs_188_io_enable)
  );
  FringeFF regs_189 ( // @[RegFile.scala 66:20:@40275.4]
    .clock(regs_189_clock),
    .reset(regs_189_reset),
    .io_in(regs_189_io_in),
    .io_reset(regs_189_io_reset),
    .io_out(regs_189_io_out),
    .io_enable(regs_189_io_enable)
  );
  FringeFF regs_190 ( // @[RegFile.scala 66:20:@40289.4]
    .clock(regs_190_clock),
    .reset(regs_190_reset),
    .io_in(regs_190_io_in),
    .io_reset(regs_190_io_reset),
    .io_out(regs_190_io_out),
    .io_enable(regs_190_io_enable)
  );
  FringeFF regs_191 ( // @[RegFile.scala 66:20:@40303.4]
    .clock(regs_191_clock),
    .reset(regs_191_reset),
    .io_in(regs_191_io_in),
    .io_reset(regs_191_io_reset),
    .io_out(regs_191_io_out),
    .io_enable(regs_191_io_enable)
  );
  FringeFF regs_192 ( // @[RegFile.scala 66:20:@40317.4]
    .clock(regs_192_clock),
    .reset(regs_192_reset),
    .io_in(regs_192_io_in),
    .io_reset(regs_192_io_reset),
    .io_out(regs_192_io_out),
    .io_enable(regs_192_io_enable)
  );
  FringeFF regs_193 ( // @[RegFile.scala 66:20:@40331.4]
    .clock(regs_193_clock),
    .reset(regs_193_reset),
    .io_in(regs_193_io_in),
    .io_reset(regs_193_io_reset),
    .io_out(regs_193_io_out),
    .io_enable(regs_193_io_enable)
  );
  FringeFF regs_194 ( // @[RegFile.scala 66:20:@40345.4]
    .clock(regs_194_clock),
    .reset(regs_194_reset),
    .io_in(regs_194_io_in),
    .io_reset(regs_194_io_reset),
    .io_out(regs_194_io_out),
    .io_enable(regs_194_io_enable)
  );
  FringeFF regs_195 ( // @[RegFile.scala 66:20:@40359.4]
    .clock(regs_195_clock),
    .reset(regs_195_reset),
    .io_in(regs_195_io_in),
    .io_reset(regs_195_io_reset),
    .io_out(regs_195_io_out),
    .io_enable(regs_195_io_enable)
  );
  FringeFF regs_196 ( // @[RegFile.scala 66:20:@40373.4]
    .clock(regs_196_clock),
    .reset(regs_196_reset),
    .io_in(regs_196_io_in),
    .io_reset(regs_196_io_reset),
    .io_out(regs_196_io_out),
    .io_enable(regs_196_io_enable)
  );
  FringeFF regs_197 ( // @[RegFile.scala 66:20:@40387.4]
    .clock(regs_197_clock),
    .reset(regs_197_reset),
    .io_in(regs_197_io_in),
    .io_reset(regs_197_io_reset),
    .io_out(regs_197_io_out),
    .io_enable(regs_197_io_enable)
  );
  FringeFF regs_198 ( // @[RegFile.scala 66:20:@40401.4]
    .clock(regs_198_clock),
    .reset(regs_198_reset),
    .io_in(regs_198_io_in),
    .io_reset(regs_198_io_reset),
    .io_out(regs_198_io_out),
    .io_enable(regs_198_io_enable)
  );
  FringeFF regs_199 ( // @[RegFile.scala 66:20:@40415.4]
    .clock(regs_199_clock),
    .reset(regs_199_reset),
    .io_in(regs_199_io_in),
    .io_reset(regs_199_io_reset),
    .io_out(regs_199_io_out),
    .io_enable(regs_199_io_enable)
  );
  FringeFF regs_200 ( // @[RegFile.scala 66:20:@40429.4]
    .clock(regs_200_clock),
    .reset(regs_200_reset),
    .io_in(regs_200_io_in),
    .io_reset(regs_200_io_reset),
    .io_out(regs_200_io_out),
    .io_enable(regs_200_io_enable)
  );
  FringeFF regs_201 ( // @[RegFile.scala 66:20:@40443.4]
    .clock(regs_201_clock),
    .reset(regs_201_reset),
    .io_in(regs_201_io_in),
    .io_reset(regs_201_io_reset),
    .io_out(regs_201_io_out),
    .io_enable(regs_201_io_enable)
  );
  FringeFF regs_202 ( // @[RegFile.scala 66:20:@40457.4]
    .clock(regs_202_clock),
    .reset(regs_202_reset),
    .io_in(regs_202_io_in),
    .io_reset(regs_202_io_reset),
    .io_out(regs_202_io_out),
    .io_enable(regs_202_io_enable)
  );
  FringeFF regs_203 ( // @[RegFile.scala 66:20:@40471.4]
    .clock(regs_203_clock),
    .reset(regs_203_reset),
    .io_in(regs_203_io_in),
    .io_reset(regs_203_io_reset),
    .io_out(regs_203_io_out),
    .io_enable(regs_203_io_enable)
  );
  FringeFF regs_204 ( // @[RegFile.scala 66:20:@40485.4]
    .clock(regs_204_clock),
    .reset(regs_204_reset),
    .io_in(regs_204_io_in),
    .io_reset(regs_204_io_reset),
    .io_out(regs_204_io_out),
    .io_enable(regs_204_io_enable)
  );
  FringeFF regs_205 ( // @[RegFile.scala 66:20:@40499.4]
    .clock(regs_205_clock),
    .reset(regs_205_reset),
    .io_in(regs_205_io_in),
    .io_reset(regs_205_io_reset),
    .io_out(regs_205_io_out),
    .io_enable(regs_205_io_enable)
  );
  FringeFF regs_206 ( // @[RegFile.scala 66:20:@40513.4]
    .clock(regs_206_clock),
    .reset(regs_206_reset),
    .io_in(regs_206_io_in),
    .io_reset(regs_206_io_reset),
    .io_out(regs_206_io_out),
    .io_enable(regs_206_io_enable)
  );
  FringeFF regs_207 ( // @[RegFile.scala 66:20:@40527.4]
    .clock(regs_207_clock),
    .reset(regs_207_reset),
    .io_in(regs_207_io_in),
    .io_reset(regs_207_io_reset),
    .io_out(regs_207_io_out),
    .io_enable(regs_207_io_enable)
  );
  FringeFF regs_208 ( // @[RegFile.scala 66:20:@40541.4]
    .clock(regs_208_clock),
    .reset(regs_208_reset),
    .io_in(regs_208_io_in),
    .io_reset(regs_208_io_reset),
    .io_out(regs_208_io_out),
    .io_enable(regs_208_io_enable)
  );
  FringeFF regs_209 ( // @[RegFile.scala 66:20:@40555.4]
    .clock(regs_209_clock),
    .reset(regs_209_reset),
    .io_in(regs_209_io_in),
    .io_reset(regs_209_io_reset),
    .io_out(regs_209_io_out),
    .io_enable(regs_209_io_enable)
  );
  FringeFF regs_210 ( // @[RegFile.scala 66:20:@40569.4]
    .clock(regs_210_clock),
    .reset(regs_210_reset),
    .io_in(regs_210_io_in),
    .io_reset(regs_210_io_reset),
    .io_out(regs_210_io_out),
    .io_enable(regs_210_io_enable)
  );
  FringeFF regs_211 ( // @[RegFile.scala 66:20:@40583.4]
    .clock(regs_211_clock),
    .reset(regs_211_reset),
    .io_in(regs_211_io_in),
    .io_reset(regs_211_io_reset),
    .io_out(regs_211_io_out),
    .io_enable(regs_211_io_enable)
  );
  FringeFF regs_212 ( // @[RegFile.scala 66:20:@40597.4]
    .clock(regs_212_clock),
    .reset(regs_212_reset),
    .io_in(regs_212_io_in),
    .io_reset(regs_212_io_reset),
    .io_out(regs_212_io_out),
    .io_enable(regs_212_io_enable)
  );
  FringeFF regs_213 ( // @[RegFile.scala 66:20:@40611.4]
    .clock(regs_213_clock),
    .reset(regs_213_reset),
    .io_in(regs_213_io_in),
    .io_reset(regs_213_io_reset),
    .io_out(regs_213_io_out),
    .io_enable(regs_213_io_enable)
  );
  FringeFF regs_214 ( // @[RegFile.scala 66:20:@40625.4]
    .clock(regs_214_clock),
    .reset(regs_214_reset),
    .io_in(regs_214_io_in),
    .io_reset(regs_214_io_reset),
    .io_out(regs_214_io_out),
    .io_enable(regs_214_io_enable)
  );
  FringeFF regs_215 ( // @[RegFile.scala 66:20:@40639.4]
    .clock(regs_215_clock),
    .reset(regs_215_reset),
    .io_in(regs_215_io_in),
    .io_reset(regs_215_io_reset),
    .io_out(regs_215_io_out),
    .io_enable(regs_215_io_enable)
  );
  FringeFF regs_216 ( // @[RegFile.scala 66:20:@40653.4]
    .clock(regs_216_clock),
    .reset(regs_216_reset),
    .io_in(regs_216_io_in),
    .io_reset(regs_216_io_reset),
    .io_out(regs_216_io_out),
    .io_enable(regs_216_io_enable)
  );
  FringeFF regs_217 ( // @[RegFile.scala 66:20:@40667.4]
    .clock(regs_217_clock),
    .reset(regs_217_reset),
    .io_in(regs_217_io_in),
    .io_reset(regs_217_io_reset),
    .io_out(regs_217_io_out),
    .io_enable(regs_217_io_enable)
  );
  FringeFF regs_218 ( // @[RegFile.scala 66:20:@40681.4]
    .clock(regs_218_clock),
    .reset(regs_218_reset),
    .io_in(regs_218_io_in),
    .io_reset(regs_218_io_reset),
    .io_out(regs_218_io_out),
    .io_enable(regs_218_io_enable)
  );
  FringeFF regs_219 ( // @[RegFile.scala 66:20:@40695.4]
    .clock(regs_219_clock),
    .reset(regs_219_reset),
    .io_in(regs_219_io_in),
    .io_reset(regs_219_io_reset),
    .io_out(regs_219_io_out),
    .io_enable(regs_219_io_enable)
  );
  FringeFF regs_220 ( // @[RegFile.scala 66:20:@40709.4]
    .clock(regs_220_clock),
    .reset(regs_220_reset),
    .io_in(regs_220_io_in),
    .io_reset(regs_220_io_reset),
    .io_out(regs_220_io_out),
    .io_enable(regs_220_io_enable)
  );
  FringeFF regs_221 ( // @[RegFile.scala 66:20:@40723.4]
    .clock(regs_221_clock),
    .reset(regs_221_reset),
    .io_in(regs_221_io_in),
    .io_reset(regs_221_io_reset),
    .io_out(regs_221_io_out),
    .io_enable(regs_221_io_enable)
  );
  FringeFF regs_222 ( // @[RegFile.scala 66:20:@40737.4]
    .clock(regs_222_clock),
    .reset(regs_222_reset),
    .io_in(regs_222_io_in),
    .io_reset(regs_222_io_reset),
    .io_out(regs_222_io_out),
    .io_enable(regs_222_io_enable)
  );
  FringeFF regs_223 ( // @[RegFile.scala 66:20:@40751.4]
    .clock(regs_223_clock),
    .reset(regs_223_reset),
    .io_in(regs_223_io_in),
    .io_reset(regs_223_io_reset),
    .io_out(regs_223_io_out),
    .io_enable(regs_223_io_enable)
  );
  FringeFF regs_224 ( // @[RegFile.scala 66:20:@40765.4]
    .clock(regs_224_clock),
    .reset(regs_224_reset),
    .io_in(regs_224_io_in),
    .io_reset(regs_224_io_reset),
    .io_out(regs_224_io_out),
    .io_enable(regs_224_io_enable)
  );
  FringeFF regs_225 ( // @[RegFile.scala 66:20:@40779.4]
    .clock(regs_225_clock),
    .reset(regs_225_reset),
    .io_in(regs_225_io_in),
    .io_reset(regs_225_io_reset),
    .io_out(regs_225_io_out),
    .io_enable(regs_225_io_enable)
  );
  FringeFF regs_226 ( // @[RegFile.scala 66:20:@40793.4]
    .clock(regs_226_clock),
    .reset(regs_226_reset),
    .io_in(regs_226_io_in),
    .io_reset(regs_226_io_reset),
    .io_out(regs_226_io_out),
    .io_enable(regs_226_io_enable)
  );
  FringeFF regs_227 ( // @[RegFile.scala 66:20:@40807.4]
    .clock(regs_227_clock),
    .reset(regs_227_reset),
    .io_in(regs_227_io_in),
    .io_reset(regs_227_io_reset),
    .io_out(regs_227_io_out),
    .io_enable(regs_227_io_enable)
  );
  FringeFF regs_228 ( // @[RegFile.scala 66:20:@40821.4]
    .clock(regs_228_clock),
    .reset(regs_228_reset),
    .io_in(regs_228_io_in),
    .io_reset(regs_228_io_reset),
    .io_out(regs_228_io_out),
    .io_enable(regs_228_io_enable)
  );
  FringeFF regs_229 ( // @[RegFile.scala 66:20:@40835.4]
    .clock(regs_229_clock),
    .reset(regs_229_reset),
    .io_in(regs_229_io_in),
    .io_reset(regs_229_io_reset),
    .io_out(regs_229_io_out),
    .io_enable(regs_229_io_enable)
  );
  FringeFF regs_230 ( // @[RegFile.scala 66:20:@40849.4]
    .clock(regs_230_clock),
    .reset(regs_230_reset),
    .io_in(regs_230_io_in),
    .io_reset(regs_230_io_reset),
    .io_out(regs_230_io_out),
    .io_enable(regs_230_io_enable)
  );
  FringeFF regs_231 ( // @[RegFile.scala 66:20:@40863.4]
    .clock(regs_231_clock),
    .reset(regs_231_reset),
    .io_in(regs_231_io_in),
    .io_reset(regs_231_io_reset),
    .io_out(regs_231_io_out),
    .io_enable(regs_231_io_enable)
  );
  FringeFF regs_232 ( // @[RegFile.scala 66:20:@40877.4]
    .clock(regs_232_clock),
    .reset(regs_232_reset),
    .io_in(regs_232_io_in),
    .io_reset(regs_232_io_reset),
    .io_out(regs_232_io_out),
    .io_enable(regs_232_io_enable)
  );
  FringeFF regs_233 ( // @[RegFile.scala 66:20:@40891.4]
    .clock(regs_233_clock),
    .reset(regs_233_reset),
    .io_in(regs_233_io_in),
    .io_reset(regs_233_io_reset),
    .io_out(regs_233_io_out),
    .io_enable(regs_233_io_enable)
  );
  FringeFF regs_234 ( // @[RegFile.scala 66:20:@40905.4]
    .clock(regs_234_clock),
    .reset(regs_234_reset),
    .io_in(regs_234_io_in),
    .io_reset(regs_234_io_reset),
    .io_out(regs_234_io_out),
    .io_enable(regs_234_io_enable)
  );
  FringeFF regs_235 ( // @[RegFile.scala 66:20:@40919.4]
    .clock(regs_235_clock),
    .reset(regs_235_reset),
    .io_in(regs_235_io_in),
    .io_reset(regs_235_io_reset),
    .io_out(regs_235_io_out),
    .io_enable(regs_235_io_enable)
  );
  FringeFF regs_236 ( // @[RegFile.scala 66:20:@40933.4]
    .clock(regs_236_clock),
    .reset(regs_236_reset),
    .io_in(regs_236_io_in),
    .io_reset(regs_236_io_reset),
    .io_out(regs_236_io_out),
    .io_enable(regs_236_io_enable)
  );
  FringeFF regs_237 ( // @[RegFile.scala 66:20:@40947.4]
    .clock(regs_237_clock),
    .reset(regs_237_reset),
    .io_in(regs_237_io_in),
    .io_reset(regs_237_io_reset),
    .io_out(regs_237_io_out),
    .io_enable(regs_237_io_enable)
  );
  FringeFF regs_238 ( // @[RegFile.scala 66:20:@40961.4]
    .clock(regs_238_clock),
    .reset(regs_238_reset),
    .io_in(regs_238_io_in),
    .io_reset(regs_238_io_reset),
    .io_out(regs_238_io_out),
    .io_enable(regs_238_io_enable)
  );
  FringeFF regs_239 ( // @[RegFile.scala 66:20:@40975.4]
    .clock(regs_239_clock),
    .reset(regs_239_reset),
    .io_in(regs_239_io_in),
    .io_reset(regs_239_io_reset),
    .io_out(regs_239_io_out),
    .io_enable(regs_239_io_enable)
  );
  FringeFF regs_240 ( // @[RegFile.scala 66:20:@40989.4]
    .clock(regs_240_clock),
    .reset(regs_240_reset),
    .io_in(regs_240_io_in),
    .io_reset(regs_240_io_reset),
    .io_out(regs_240_io_out),
    .io_enable(regs_240_io_enable)
  );
  FringeFF regs_241 ( // @[RegFile.scala 66:20:@41003.4]
    .clock(regs_241_clock),
    .reset(regs_241_reset),
    .io_in(regs_241_io_in),
    .io_reset(regs_241_io_reset),
    .io_out(regs_241_io_out),
    .io_enable(regs_241_io_enable)
  );
  FringeFF regs_242 ( // @[RegFile.scala 66:20:@41017.4]
    .clock(regs_242_clock),
    .reset(regs_242_reset),
    .io_in(regs_242_io_in),
    .io_reset(regs_242_io_reset),
    .io_out(regs_242_io_out),
    .io_enable(regs_242_io_enable)
  );
  FringeFF regs_243 ( // @[RegFile.scala 66:20:@41031.4]
    .clock(regs_243_clock),
    .reset(regs_243_reset),
    .io_in(regs_243_io_in),
    .io_reset(regs_243_io_reset),
    .io_out(regs_243_io_out),
    .io_enable(regs_243_io_enable)
  );
  FringeFF regs_244 ( // @[RegFile.scala 66:20:@41045.4]
    .clock(regs_244_clock),
    .reset(regs_244_reset),
    .io_in(regs_244_io_in),
    .io_reset(regs_244_io_reset),
    .io_out(regs_244_io_out),
    .io_enable(regs_244_io_enable)
  );
  FringeFF regs_245 ( // @[RegFile.scala 66:20:@41059.4]
    .clock(regs_245_clock),
    .reset(regs_245_reset),
    .io_in(regs_245_io_in),
    .io_reset(regs_245_io_reset),
    .io_out(regs_245_io_out),
    .io_enable(regs_245_io_enable)
  );
  FringeFF regs_246 ( // @[RegFile.scala 66:20:@41073.4]
    .clock(regs_246_clock),
    .reset(regs_246_reset),
    .io_in(regs_246_io_in),
    .io_reset(regs_246_io_reset),
    .io_out(regs_246_io_out),
    .io_enable(regs_246_io_enable)
  );
  FringeFF regs_247 ( // @[RegFile.scala 66:20:@41087.4]
    .clock(regs_247_clock),
    .reset(regs_247_reset),
    .io_in(regs_247_io_in),
    .io_reset(regs_247_io_reset),
    .io_out(regs_247_io_out),
    .io_enable(regs_247_io_enable)
  );
  FringeFF regs_248 ( // @[RegFile.scala 66:20:@41101.4]
    .clock(regs_248_clock),
    .reset(regs_248_reset),
    .io_in(regs_248_io_in),
    .io_reset(regs_248_io_reset),
    .io_out(regs_248_io_out),
    .io_enable(regs_248_io_enable)
  );
  FringeFF regs_249 ( // @[RegFile.scala 66:20:@41115.4]
    .clock(regs_249_clock),
    .reset(regs_249_reset),
    .io_in(regs_249_io_in),
    .io_reset(regs_249_io_reset),
    .io_out(regs_249_io_out),
    .io_enable(regs_249_io_enable)
  );
  FringeFF regs_250 ( // @[RegFile.scala 66:20:@41129.4]
    .clock(regs_250_clock),
    .reset(regs_250_reset),
    .io_in(regs_250_io_in),
    .io_reset(regs_250_io_reset),
    .io_out(regs_250_io_out),
    .io_enable(regs_250_io_enable)
  );
  FringeFF regs_251 ( // @[RegFile.scala 66:20:@41143.4]
    .clock(regs_251_clock),
    .reset(regs_251_reset),
    .io_in(regs_251_io_in),
    .io_reset(regs_251_io_reset),
    .io_out(regs_251_io_out),
    .io_enable(regs_251_io_enable)
  );
  FringeFF regs_252 ( // @[RegFile.scala 66:20:@41157.4]
    .clock(regs_252_clock),
    .reset(regs_252_reset),
    .io_in(regs_252_io_in),
    .io_reset(regs_252_io_reset),
    .io_out(regs_252_io_out),
    .io_enable(regs_252_io_enable)
  );
  FringeFF regs_253 ( // @[RegFile.scala 66:20:@41171.4]
    .clock(regs_253_clock),
    .reset(regs_253_reset),
    .io_in(regs_253_io_in),
    .io_reset(regs_253_io_reset),
    .io_out(regs_253_io_out),
    .io_enable(regs_253_io_enable)
  );
  FringeFF regs_254 ( // @[RegFile.scala 66:20:@41185.4]
    .clock(regs_254_clock),
    .reset(regs_254_reset),
    .io_in(regs_254_io_in),
    .io_reset(regs_254_io_reset),
    .io_out(regs_254_io_out),
    .io_enable(regs_254_io_enable)
  );
  FringeFF regs_255 ( // @[RegFile.scala 66:20:@41199.4]
    .clock(regs_255_clock),
    .reset(regs_255_reset),
    .io_in(regs_255_io_in),
    .io_reset(regs_255_io_reset),
    .io_out(regs_255_io_out),
    .io_enable(regs_255_io_enable)
  );
  FringeFF regs_256 ( // @[RegFile.scala 66:20:@41213.4]
    .clock(regs_256_clock),
    .reset(regs_256_reset),
    .io_in(regs_256_io_in),
    .io_reset(regs_256_io_reset),
    .io_out(regs_256_io_out),
    .io_enable(regs_256_io_enable)
  );
  FringeFF regs_257 ( // @[RegFile.scala 66:20:@41227.4]
    .clock(regs_257_clock),
    .reset(regs_257_reset),
    .io_in(regs_257_io_in),
    .io_reset(regs_257_io_reset),
    .io_out(regs_257_io_out),
    .io_enable(regs_257_io_enable)
  );
  FringeFF regs_258 ( // @[RegFile.scala 66:20:@41241.4]
    .clock(regs_258_clock),
    .reset(regs_258_reset),
    .io_in(regs_258_io_in),
    .io_reset(regs_258_io_reset),
    .io_out(regs_258_io_out),
    .io_enable(regs_258_io_enable)
  );
  FringeFF regs_259 ( // @[RegFile.scala 66:20:@41255.4]
    .clock(regs_259_clock),
    .reset(regs_259_reset),
    .io_in(regs_259_io_in),
    .io_reset(regs_259_io_reset),
    .io_out(regs_259_io_out),
    .io_enable(regs_259_io_enable)
  );
  FringeFF regs_260 ( // @[RegFile.scala 66:20:@41269.4]
    .clock(regs_260_clock),
    .reset(regs_260_reset),
    .io_in(regs_260_io_in),
    .io_reset(regs_260_io_reset),
    .io_out(regs_260_io_out),
    .io_enable(regs_260_io_enable)
  );
  FringeFF regs_261 ( // @[RegFile.scala 66:20:@41283.4]
    .clock(regs_261_clock),
    .reset(regs_261_reset),
    .io_in(regs_261_io_in),
    .io_reset(regs_261_io_reset),
    .io_out(regs_261_io_out),
    .io_enable(regs_261_io_enable)
  );
  FringeFF regs_262 ( // @[RegFile.scala 66:20:@41297.4]
    .clock(regs_262_clock),
    .reset(regs_262_reset),
    .io_in(regs_262_io_in),
    .io_reset(regs_262_io_reset),
    .io_out(regs_262_io_out),
    .io_enable(regs_262_io_enable)
  );
  FringeFF regs_263 ( // @[RegFile.scala 66:20:@41311.4]
    .clock(regs_263_clock),
    .reset(regs_263_reset),
    .io_in(regs_263_io_in),
    .io_reset(regs_263_io_reset),
    .io_out(regs_263_io_out),
    .io_enable(regs_263_io_enable)
  );
  FringeFF regs_264 ( // @[RegFile.scala 66:20:@41325.4]
    .clock(regs_264_clock),
    .reset(regs_264_reset),
    .io_in(regs_264_io_in),
    .io_reset(regs_264_io_reset),
    .io_out(regs_264_io_out),
    .io_enable(regs_264_io_enable)
  );
  FringeFF regs_265 ( // @[RegFile.scala 66:20:@41339.4]
    .clock(regs_265_clock),
    .reset(regs_265_reset),
    .io_in(regs_265_io_in),
    .io_reset(regs_265_io_reset),
    .io_out(regs_265_io_out),
    .io_enable(regs_265_io_enable)
  );
  FringeFF regs_266 ( // @[RegFile.scala 66:20:@41353.4]
    .clock(regs_266_clock),
    .reset(regs_266_reset),
    .io_in(regs_266_io_in),
    .io_reset(regs_266_io_reset),
    .io_out(regs_266_io_out),
    .io_enable(regs_266_io_enable)
  );
  FringeFF regs_267 ( // @[RegFile.scala 66:20:@41367.4]
    .clock(regs_267_clock),
    .reset(regs_267_reset),
    .io_in(regs_267_io_in),
    .io_reset(regs_267_io_reset),
    .io_out(regs_267_io_out),
    .io_enable(regs_267_io_enable)
  );
  FringeFF regs_268 ( // @[RegFile.scala 66:20:@41381.4]
    .clock(regs_268_clock),
    .reset(regs_268_reset),
    .io_in(regs_268_io_in),
    .io_reset(regs_268_io_reset),
    .io_out(regs_268_io_out),
    .io_enable(regs_268_io_enable)
  );
  FringeFF regs_269 ( // @[RegFile.scala 66:20:@41395.4]
    .clock(regs_269_clock),
    .reset(regs_269_reset),
    .io_in(regs_269_io_in),
    .io_reset(regs_269_io_reset),
    .io_out(regs_269_io_out),
    .io_enable(regs_269_io_enable)
  );
  FringeFF regs_270 ( // @[RegFile.scala 66:20:@41409.4]
    .clock(regs_270_clock),
    .reset(regs_270_reset),
    .io_in(regs_270_io_in),
    .io_reset(regs_270_io_reset),
    .io_out(regs_270_io_out),
    .io_enable(regs_270_io_enable)
  );
  FringeFF regs_271 ( // @[RegFile.scala 66:20:@41423.4]
    .clock(regs_271_clock),
    .reset(regs_271_reset),
    .io_in(regs_271_io_in),
    .io_reset(regs_271_io_reset),
    .io_out(regs_271_io_out),
    .io_enable(regs_271_io_enable)
  );
  FringeFF regs_272 ( // @[RegFile.scala 66:20:@41437.4]
    .clock(regs_272_clock),
    .reset(regs_272_reset),
    .io_in(regs_272_io_in),
    .io_reset(regs_272_io_reset),
    .io_out(regs_272_io_out),
    .io_enable(regs_272_io_enable)
  );
  FringeFF regs_273 ( // @[RegFile.scala 66:20:@41451.4]
    .clock(regs_273_clock),
    .reset(regs_273_reset),
    .io_in(regs_273_io_in),
    .io_reset(regs_273_io_reset),
    .io_out(regs_273_io_out),
    .io_enable(regs_273_io_enable)
  );
  FringeFF regs_274 ( // @[RegFile.scala 66:20:@41465.4]
    .clock(regs_274_clock),
    .reset(regs_274_reset),
    .io_in(regs_274_io_in),
    .io_reset(regs_274_io_reset),
    .io_out(regs_274_io_out),
    .io_enable(regs_274_io_enable)
  );
  FringeFF regs_275 ( // @[RegFile.scala 66:20:@41479.4]
    .clock(regs_275_clock),
    .reset(regs_275_reset),
    .io_in(regs_275_io_in),
    .io_reset(regs_275_io_reset),
    .io_out(regs_275_io_out),
    .io_enable(regs_275_io_enable)
  );
  FringeFF regs_276 ( // @[RegFile.scala 66:20:@41493.4]
    .clock(regs_276_clock),
    .reset(regs_276_reset),
    .io_in(regs_276_io_in),
    .io_reset(regs_276_io_reset),
    .io_out(regs_276_io_out),
    .io_enable(regs_276_io_enable)
  );
  FringeFF regs_277 ( // @[RegFile.scala 66:20:@41507.4]
    .clock(regs_277_clock),
    .reset(regs_277_reset),
    .io_in(regs_277_io_in),
    .io_reset(regs_277_io_reset),
    .io_out(regs_277_io_out),
    .io_enable(regs_277_io_enable)
  );
  FringeFF regs_278 ( // @[RegFile.scala 66:20:@41521.4]
    .clock(regs_278_clock),
    .reset(regs_278_reset),
    .io_in(regs_278_io_in),
    .io_reset(regs_278_io_reset),
    .io_out(regs_278_io_out),
    .io_enable(regs_278_io_enable)
  );
  FringeFF regs_279 ( // @[RegFile.scala 66:20:@41535.4]
    .clock(regs_279_clock),
    .reset(regs_279_reset),
    .io_in(regs_279_io_in),
    .io_reset(regs_279_io_reset),
    .io_out(regs_279_io_out),
    .io_enable(regs_279_io_enable)
  );
  FringeFF regs_280 ( // @[RegFile.scala 66:20:@41549.4]
    .clock(regs_280_clock),
    .reset(regs_280_reset),
    .io_in(regs_280_io_in),
    .io_reset(regs_280_io_reset),
    .io_out(regs_280_io_out),
    .io_enable(regs_280_io_enable)
  );
  FringeFF regs_281 ( // @[RegFile.scala 66:20:@41563.4]
    .clock(regs_281_clock),
    .reset(regs_281_reset),
    .io_in(regs_281_io_in),
    .io_reset(regs_281_io_reset),
    .io_out(regs_281_io_out),
    .io_enable(regs_281_io_enable)
  );
  FringeFF regs_282 ( // @[RegFile.scala 66:20:@41577.4]
    .clock(regs_282_clock),
    .reset(regs_282_reset),
    .io_in(regs_282_io_in),
    .io_reset(regs_282_io_reset),
    .io_out(regs_282_io_out),
    .io_enable(regs_282_io_enable)
  );
  FringeFF regs_283 ( // @[RegFile.scala 66:20:@41591.4]
    .clock(regs_283_clock),
    .reset(regs_283_reset),
    .io_in(regs_283_io_in),
    .io_reset(regs_283_io_reset),
    .io_out(regs_283_io_out),
    .io_enable(regs_283_io_enable)
  );
  FringeFF regs_284 ( // @[RegFile.scala 66:20:@41605.4]
    .clock(regs_284_clock),
    .reset(regs_284_reset),
    .io_in(regs_284_io_in),
    .io_reset(regs_284_io_reset),
    .io_out(regs_284_io_out),
    .io_enable(regs_284_io_enable)
  );
  FringeFF regs_285 ( // @[RegFile.scala 66:20:@41619.4]
    .clock(regs_285_clock),
    .reset(regs_285_reset),
    .io_in(regs_285_io_in),
    .io_reset(regs_285_io_reset),
    .io_out(regs_285_io_out),
    .io_enable(regs_285_io_enable)
  );
  FringeFF regs_286 ( // @[RegFile.scala 66:20:@41633.4]
    .clock(regs_286_clock),
    .reset(regs_286_reset),
    .io_in(regs_286_io_in),
    .io_reset(regs_286_io_reset),
    .io_out(regs_286_io_out),
    .io_enable(regs_286_io_enable)
  );
  FringeFF regs_287 ( // @[RegFile.scala 66:20:@41647.4]
    .clock(regs_287_clock),
    .reset(regs_287_reset),
    .io_in(regs_287_io_in),
    .io_reset(regs_287_io_reset),
    .io_out(regs_287_io_out),
    .io_enable(regs_287_io_enable)
  );
  FringeFF regs_288 ( // @[RegFile.scala 66:20:@41661.4]
    .clock(regs_288_clock),
    .reset(regs_288_reset),
    .io_in(regs_288_io_in),
    .io_reset(regs_288_io_reset),
    .io_out(regs_288_io_out),
    .io_enable(regs_288_io_enable)
  );
  FringeFF regs_289 ( // @[RegFile.scala 66:20:@41675.4]
    .clock(regs_289_clock),
    .reset(regs_289_reset),
    .io_in(regs_289_io_in),
    .io_reset(regs_289_io_reset),
    .io_out(regs_289_io_out),
    .io_enable(regs_289_io_enable)
  );
  FringeFF regs_290 ( // @[RegFile.scala 66:20:@41689.4]
    .clock(regs_290_clock),
    .reset(regs_290_reset),
    .io_in(regs_290_io_in),
    .io_reset(regs_290_io_reset),
    .io_out(regs_290_io_out),
    .io_enable(regs_290_io_enable)
  );
  FringeFF regs_291 ( // @[RegFile.scala 66:20:@41703.4]
    .clock(regs_291_clock),
    .reset(regs_291_reset),
    .io_in(regs_291_io_in),
    .io_reset(regs_291_io_reset),
    .io_out(regs_291_io_out),
    .io_enable(regs_291_io_enable)
  );
  FringeFF regs_292 ( // @[RegFile.scala 66:20:@41717.4]
    .clock(regs_292_clock),
    .reset(regs_292_reset),
    .io_in(regs_292_io_in),
    .io_reset(regs_292_io_reset),
    .io_out(regs_292_io_out),
    .io_enable(regs_292_io_enable)
  );
  FringeFF regs_293 ( // @[RegFile.scala 66:20:@41731.4]
    .clock(regs_293_clock),
    .reset(regs_293_reset),
    .io_in(regs_293_io_in),
    .io_reset(regs_293_io_reset),
    .io_out(regs_293_io_out),
    .io_enable(regs_293_io_enable)
  );
  FringeFF regs_294 ( // @[RegFile.scala 66:20:@41745.4]
    .clock(regs_294_clock),
    .reset(regs_294_reset),
    .io_in(regs_294_io_in),
    .io_reset(regs_294_io_reset),
    .io_out(regs_294_io_out),
    .io_enable(regs_294_io_enable)
  );
  FringeFF regs_295 ( // @[RegFile.scala 66:20:@41759.4]
    .clock(regs_295_clock),
    .reset(regs_295_reset),
    .io_in(regs_295_io_in),
    .io_reset(regs_295_io_reset),
    .io_out(regs_295_io_out),
    .io_enable(regs_295_io_enable)
  );
  FringeFF regs_296 ( // @[RegFile.scala 66:20:@41773.4]
    .clock(regs_296_clock),
    .reset(regs_296_reset),
    .io_in(regs_296_io_in),
    .io_reset(regs_296_io_reset),
    .io_out(regs_296_io_out),
    .io_enable(regs_296_io_enable)
  );
  FringeFF regs_297 ( // @[RegFile.scala 66:20:@41787.4]
    .clock(regs_297_clock),
    .reset(regs_297_reset),
    .io_in(regs_297_io_in),
    .io_reset(regs_297_io_reset),
    .io_out(regs_297_io_out),
    .io_enable(regs_297_io_enable)
  );
  FringeFF regs_298 ( // @[RegFile.scala 66:20:@41801.4]
    .clock(regs_298_clock),
    .reset(regs_298_reset),
    .io_in(regs_298_io_in),
    .io_reset(regs_298_io_reset),
    .io_out(regs_298_io_out),
    .io_enable(regs_298_io_enable)
  );
  FringeFF regs_299 ( // @[RegFile.scala 66:20:@41815.4]
    .clock(regs_299_clock),
    .reset(regs_299_reset),
    .io_in(regs_299_io_in),
    .io_reset(regs_299_io_reset),
    .io_out(regs_299_io_out),
    .io_enable(regs_299_io_enable)
  );
  FringeFF regs_300 ( // @[RegFile.scala 66:20:@41829.4]
    .clock(regs_300_clock),
    .reset(regs_300_reset),
    .io_in(regs_300_io_in),
    .io_reset(regs_300_io_reset),
    .io_out(regs_300_io_out),
    .io_enable(regs_300_io_enable)
  );
  FringeFF regs_301 ( // @[RegFile.scala 66:20:@41843.4]
    .clock(regs_301_clock),
    .reset(regs_301_reset),
    .io_in(regs_301_io_in),
    .io_reset(regs_301_io_reset),
    .io_out(regs_301_io_out),
    .io_enable(regs_301_io_enable)
  );
  FringeFF regs_302 ( // @[RegFile.scala 66:20:@41857.4]
    .clock(regs_302_clock),
    .reset(regs_302_reset),
    .io_in(regs_302_io_in),
    .io_reset(regs_302_io_reset),
    .io_out(regs_302_io_out),
    .io_enable(regs_302_io_enable)
  );
  FringeFF regs_303 ( // @[RegFile.scala 66:20:@41871.4]
    .clock(regs_303_clock),
    .reset(regs_303_reset),
    .io_in(regs_303_io_in),
    .io_reset(regs_303_io_reset),
    .io_out(regs_303_io_out),
    .io_enable(regs_303_io_enable)
  );
  FringeFF regs_304 ( // @[RegFile.scala 66:20:@41885.4]
    .clock(regs_304_clock),
    .reset(regs_304_reset),
    .io_in(regs_304_io_in),
    .io_reset(regs_304_io_reset),
    .io_out(regs_304_io_out),
    .io_enable(regs_304_io_enable)
  );
  FringeFF regs_305 ( // @[RegFile.scala 66:20:@41899.4]
    .clock(regs_305_clock),
    .reset(regs_305_reset),
    .io_in(regs_305_io_in),
    .io_reset(regs_305_io_reset),
    .io_out(regs_305_io_out),
    .io_enable(regs_305_io_enable)
  );
  FringeFF regs_306 ( // @[RegFile.scala 66:20:@41913.4]
    .clock(regs_306_clock),
    .reset(regs_306_reset),
    .io_in(regs_306_io_in),
    .io_reset(regs_306_io_reset),
    .io_out(regs_306_io_out),
    .io_enable(regs_306_io_enable)
  );
  FringeFF regs_307 ( // @[RegFile.scala 66:20:@41927.4]
    .clock(regs_307_clock),
    .reset(regs_307_reset),
    .io_in(regs_307_io_in),
    .io_reset(regs_307_io_reset),
    .io_out(regs_307_io_out),
    .io_enable(regs_307_io_enable)
  );
  FringeFF regs_308 ( // @[RegFile.scala 66:20:@41941.4]
    .clock(regs_308_clock),
    .reset(regs_308_reset),
    .io_in(regs_308_io_in),
    .io_reset(regs_308_io_reset),
    .io_out(regs_308_io_out),
    .io_enable(regs_308_io_enable)
  );
  FringeFF regs_309 ( // @[RegFile.scala 66:20:@41955.4]
    .clock(regs_309_clock),
    .reset(regs_309_reset),
    .io_in(regs_309_io_in),
    .io_reset(regs_309_io_reset),
    .io_out(regs_309_io_out),
    .io_enable(regs_309_io_enable)
  );
  FringeFF regs_310 ( // @[RegFile.scala 66:20:@41969.4]
    .clock(regs_310_clock),
    .reset(regs_310_reset),
    .io_in(regs_310_io_in),
    .io_reset(regs_310_io_reset),
    .io_out(regs_310_io_out),
    .io_enable(regs_310_io_enable)
  );
  FringeFF regs_311 ( // @[RegFile.scala 66:20:@41983.4]
    .clock(regs_311_clock),
    .reset(regs_311_reset),
    .io_in(regs_311_io_in),
    .io_reset(regs_311_io_reset),
    .io_out(regs_311_io_out),
    .io_enable(regs_311_io_enable)
  );
  FringeFF regs_312 ( // @[RegFile.scala 66:20:@41997.4]
    .clock(regs_312_clock),
    .reset(regs_312_reset),
    .io_in(regs_312_io_in),
    .io_reset(regs_312_io_reset),
    .io_out(regs_312_io_out),
    .io_enable(regs_312_io_enable)
  );
  FringeFF regs_313 ( // @[RegFile.scala 66:20:@42011.4]
    .clock(regs_313_clock),
    .reset(regs_313_reset),
    .io_in(regs_313_io_in),
    .io_reset(regs_313_io_reset),
    .io_out(regs_313_io_out),
    .io_enable(regs_313_io_enable)
  );
  FringeFF regs_314 ( // @[RegFile.scala 66:20:@42025.4]
    .clock(regs_314_clock),
    .reset(regs_314_reset),
    .io_in(regs_314_io_in),
    .io_reset(regs_314_io_reset),
    .io_out(regs_314_io_out),
    .io_enable(regs_314_io_enable)
  );
  FringeFF regs_315 ( // @[RegFile.scala 66:20:@42039.4]
    .clock(regs_315_clock),
    .reset(regs_315_reset),
    .io_in(regs_315_io_in),
    .io_reset(regs_315_io_reset),
    .io_out(regs_315_io_out),
    .io_enable(regs_315_io_enable)
  );
  FringeFF regs_316 ( // @[RegFile.scala 66:20:@42053.4]
    .clock(regs_316_clock),
    .reset(regs_316_reset),
    .io_in(regs_316_io_in),
    .io_reset(regs_316_io_reset),
    .io_out(regs_316_io_out),
    .io_enable(regs_316_io_enable)
  );
  FringeFF regs_317 ( // @[RegFile.scala 66:20:@42067.4]
    .clock(regs_317_clock),
    .reset(regs_317_reset),
    .io_in(regs_317_io_in),
    .io_reset(regs_317_io_reset),
    .io_out(regs_317_io_out),
    .io_enable(regs_317_io_enable)
  );
  FringeFF regs_318 ( // @[RegFile.scala 66:20:@42081.4]
    .clock(regs_318_clock),
    .reset(regs_318_reset),
    .io_in(regs_318_io_in),
    .io_reset(regs_318_io_reset),
    .io_out(regs_318_io_out),
    .io_enable(regs_318_io_enable)
  );
  FringeFF regs_319 ( // @[RegFile.scala 66:20:@42095.4]
    .clock(regs_319_clock),
    .reset(regs_319_reset),
    .io_in(regs_319_io_in),
    .io_reset(regs_319_io_reset),
    .io_out(regs_319_io_out),
    .io_enable(regs_319_io_enable)
  );
  FringeFF regs_320 ( // @[RegFile.scala 66:20:@42109.4]
    .clock(regs_320_clock),
    .reset(regs_320_reset),
    .io_in(regs_320_io_in),
    .io_reset(regs_320_io_reset),
    .io_out(regs_320_io_out),
    .io_enable(regs_320_io_enable)
  );
  FringeFF regs_321 ( // @[RegFile.scala 66:20:@42123.4]
    .clock(regs_321_clock),
    .reset(regs_321_reset),
    .io_in(regs_321_io_in),
    .io_reset(regs_321_io_reset),
    .io_out(regs_321_io_out),
    .io_enable(regs_321_io_enable)
  );
  FringeFF regs_322 ( // @[RegFile.scala 66:20:@42137.4]
    .clock(regs_322_clock),
    .reset(regs_322_reset),
    .io_in(regs_322_io_in),
    .io_reset(regs_322_io_reset),
    .io_out(regs_322_io_out),
    .io_enable(regs_322_io_enable)
  );
  FringeFF regs_323 ( // @[RegFile.scala 66:20:@42151.4]
    .clock(regs_323_clock),
    .reset(regs_323_reset),
    .io_in(regs_323_io_in),
    .io_reset(regs_323_io_reset),
    .io_out(regs_323_io_out),
    .io_enable(regs_323_io_enable)
  );
  FringeFF regs_324 ( // @[RegFile.scala 66:20:@42165.4]
    .clock(regs_324_clock),
    .reset(regs_324_reset),
    .io_in(regs_324_io_in),
    .io_reset(regs_324_io_reset),
    .io_out(regs_324_io_out),
    .io_enable(regs_324_io_enable)
  );
  FringeFF regs_325 ( // @[RegFile.scala 66:20:@42179.4]
    .clock(regs_325_clock),
    .reset(regs_325_reset),
    .io_in(regs_325_io_in),
    .io_reset(regs_325_io_reset),
    .io_out(regs_325_io_out),
    .io_enable(regs_325_io_enable)
  );
  FringeFF regs_326 ( // @[RegFile.scala 66:20:@42193.4]
    .clock(regs_326_clock),
    .reset(regs_326_reset),
    .io_in(regs_326_io_in),
    .io_reset(regs_326_io_reset),
    .io_out(regs_326_io_out),
    .io_enable(regs_326_io_enable)
  );
  FringeFF regs_327 ( // @[RegFile.scala 66:20:@42207.4]
    .clock(regs_327_clock),
    .reset(regs_327_reset),
    .io_in(regs_327_io_in),
    .io_reset(regs_327_io_reset),
    .io_out(regs_327_io_out),
    .io_enable(regs_327_io_enable)
  );
  FringeFF regs_328 ( // @[RegFile.scala 66:20:@42221.4]
    .clock(regs_328_clock),
    .reset(regs_328_reset),
    .io_in(regs_328_io_in),
    .io_reset(regs_328_io_reset),
    .io_out(regs_328_io_out),
    .io_enable(regs_328_io_enable)
  );
  FringeFF regs_329 ( // @[RegFile.scala 66:20:@42235.4]
    .clock(regs_329_clock),
    .reset(regs_329_reset),
    .io_in(regs_329_io_in),
    .io_reset(regs_329_io_reset),
    .io_out(regs_329_io_out),
    .io_enable(regs_329_io_enable)
  );
  FringeFF regs_330 ( // @[RegFile.scala 66:20:@42249.4]
    .clock(regs_330_clock),
    .reset(regs_330_reset),
    .io_in(regs_330_io_in),
    .io_reset(regs_330_io_reset),
    .io_out(regs_330_io_out),
    .io_enable(regs_330_io_enable)
  );
  FringeFF regs_331 ( // @[RegFile.scala 66:20:@42263.4]
    .clock(regs_331_clock),
    .reset(regs_331_reset),
    .io_in(regs_331_io_in),
    .io_reset(regs_331_io_reset),
    .io_out(regs_331_io_out),
    .io_enable(regs_331_io_enable)
  );
  FringeFF regs_332 ( // @[RegFile.scala 66:20:@42277.4]
    .clock(regs_332_clock),
    .reset(regs_332_reset),
    .io_in(regs_332_io_in),
    .io_reset(regs_332_io_reset),
    .io_out(regs_332_io_out),
    .io_enable(regs_332_io_enable)
  );
  FringeFF regs_333 ( // @[RegFile.scala 66:20:@42291.4]
    .clock(regs_333_clock),
    .reset(regs_333_reset),
    .io_in(regs_333_io_in),
    .io_reset(regs_333_io_reset),
    .io_out(regs_333_io_out),
    .io_enable(regs_333_io_enable)
  );
  FringeFF regs_334 ( // @[RegFile.scala 66:20:@42305.4]
    .clock(regs_334_clock),
    .reset(regs_334_reset),
    .io_in(regs_334_io_in),
    .io_reset(regs_334_io_reset),
    .io_out(regs_334_io_out),
    .io_enable(regs_334_io_enable)
  );
  FringeFF regs_335 ( // @[RegFile.scala 66:20:@42319.4]
    .clock(regs_335_clock),
    .reset(regs_335_reset),
    .io_in(regs_335_io_in),
    .io_reset(regs_335_io_reset),
    .io_out(regs_335_io_out),
    .io_enable(regs_335_io_enable)
  );
  FringeFF regs_336 ( // @[RegFile.scala 66:20:@42333.4]
    .clock(regs_336_clock),
    .reset(regs_336_reset),
    .io_in(regs_336_io_in),
    .io_reset(regs_336_io_reset),
    .io_out(regs_336_io_out),
    .io_enable(regs_336_io_enable)
  );
  FringeFF regs_337 ( // @[RegFile.scala 66:20:@42347.4]
    .clock(regs_337_clock),
    .reset(regs_337_reset),
    .io_in(regs_337_io_in),
    .io_reset(regs_337_io_reset),
    .io_out(regs_337_io_out),
    .io_enable(regs_337_io_enable)
  );
  FringeFF regs_338 ( // @[RegFile.scala 66:20:@42361.4]
    .clock(regs_338_clock),
    .reset(regs_338_reset),
    .io_in(regs_338_io_in),
    .io_reset(regs_338_io_reset),
    .io_out(regs_338_io_out),
    .io_enable(regs_338_io_enable)
  );
  FringeFF regs_339 ( // @[RegFile.scala 66:20:@42375.4]
    .clock(regs_339_clock),
    .reset(regs_339_reset),
    .io_in(regs_339_io_in),
    .io_reset(regs_339_io_reset),
    .io_out(regs_339_io_out),
    .io_enable(regs_339_io_enable)
  );
  FringeFF regs_340 ( // @[RegFile.scala 66:20:@42389.4]
    .clock(regs_340_clock),
    .reset(regs_340_reset),
    .io_in(regs_340_io_in),
    .io_reset(regs_340_io_reset),
    .io_out(regs_340_io_out),
    .io_enable(regs_340_io_enable)
  );
  FringeFF regs_341 ( // @[RegFile.scala 66:20:@42403.4]
    .clock(regs_341_clock),
    .reset(regs_341_reset),
    .io_in(regs_341_io_in),
    .io_reset(regs_341_io_reset),
    .io_out(regs_341_io_out),
    .io_enable(regs_341_io_enable)
  );
  FringeFF regs_342 ( // @[RegFile.scala 66:20:@42417.4]
    .clock(regs_342_clock),
    .reset(regs_342_reset),
    .io_in(regs_342_io_in),
    .io_reset(regs_342_io_reset),
    .io_out(regs_342_io_out),
    .io_enable(regs_342_io_enable)
  );
  FringeFF regs_343 ( // @[RegFile.scala 66:20:@42431.4]
    .clock(regs_343_clock),
    .reset(regs_343_reset),
    .io_in(regs_343_io_in),
    .io_reset(regs_343_io_reset),
    .io_out(regs_343_io_out),
    .io_enable(regs_343_io_enable)
  );
  FringeFF regs_344 ( // @[RegFile.scala 66:20:@42445.4]
    .clock(regs_344_clock),
    .reset(regs_344_reset),
    .io_in(regs_344_io_in),
    .io_reset(regs_344_io_reset),
    .io_out(regs_344_io_out),
    .io_enable(regs_344_io_enable)
  );
  FringeFF regs_345 ( // @[RegFile.scala 66:20:@42459.4]
    .clock(regs_345_clock),
    .reset(regs_345_reset),
    .io_in(regs_345_io_in),
    .io_reset(regs_345_io_reset),
    .io_out(regs_345_io_out),
    .io_enable(regs_345_io_enable)
  );
  FringeFF regs_346 ( // @[RegFile.scala 66:20:@42473.4]
    .clock(regs_346_clock),
    .reset(regs_346_reset),
    .io_in(regs_346_io_in),
    .io_reset(regs_346_io_reset),
    .io_out(regs_346_io_out),
    .io_enable(regs_346_io_enable)
  );
  FringeFF regs_347 ( // @[RegFile.scala 66:20:@42487.4]
    .clock(regs_347_clock),
    .reset(regs_347_reset),
    .io_in(regs_347_io_in),
    .io_reset(regs_347_io_reset),
    .io_out(regs_347_io_out),
    .io_enable(regs_347_io_enable)
  );
  FringeFF regs_348 ( // @[RegFile.scala 66:20:@42501.4]
    .clock(regs_348_clock),
    .reset(regs_348_reset),
    .io_in(regs_348_io_in),
    .io_reset(regs_348_io_reset),
    .io_out(regs_348_io_out),
    .io_enable(regs_348_io_enable)
  );
  FringeFF regs_349 ( // @[RegFile.scala 66:20:@42515.4]
    .clock(regs_349_clock),
    .reset(regs_349_reset),
    .io_in(regs_349_io_in),
    .io_reset(regs_349_io_reset),
    .io_out(regs_349_io_out),
    .io_enable(regs_349_io_enable)
  );
  FringeFF regs_350 ( // @[RegFile.scala 66:20:@42529.4]
    .clock(regs_350_clock),
    .reset(regs_350_reset),
    .io_in(regs_350_io_in),
    .io_reset(regs_350_io_reset),
    .io_out(regs_350_io_out),
    .io_enable(regs_350_io_enable)
  );
  FringeFF regs_351 ( // @[RegFile.scala 66:20:@42543.4]
    .clock(regs_351_clock),
    .reset(regs_351_reset),
    .io_in(regs_351_io_in),
    .io_reset(regs_351_io_reset),
    .io_out(regs_351_io_out),
    .io_enable(regs_351_io_enable)
  );
  FringeFF regs_352 ( // @[RegFile.scala 66:20:@42557.4]
    .clock(regs_352_clock),
    .reset(regs_352_reset),
    .io_in(regs_352_io_in),
    .io_reset(regs_352_io_reset),
    .io_out(regs_352_io_out),
    .io_enable(regs_352_io_enable)
  );
  FringeFF regs_353 ( // @[RegFile.scala 66:20:@42571.4]
    .clock(regs_353_clock),
    .reset(regs_353_reset),
    .io_in(regs_353_io_in),
    .io_reset(regs_353_io_reset),
    .io_out(regs_353_io_out),
    .io_enable(regs_353_io_enable)
  );
  FringeFF regs_354 ( // @[RegFile.scala 66:20:@42585.4]
    .clock(regs_354_clock),
    .reset(regs_354_reset),
    .io_in(regs_354_io_in),
    .io_reset(regs_354_io_reset),
    .io_out(regs_354_io_out),
    .io_enable(regs_354_io_enable)
  );
  FringeFF regs_355 ( // @[RegFile.scala 66:20:@42599.4]
    .clock(regs_355_clock),
    .reset(regs_355_reset),
    .io_in(regs_355_io_in),
    .io_reset(regs_355_io_reset),
    .io_out(regs_355_io_out),
    .io_enable(regs_355_io_enable)
  );
  FringeFF regs_356 ( // @[RegFile.scala 66:20:@42613.4]
    .clock(regs_356_clock),
    .reset(regs_356_reset),
    .io_in(regs_356_io_in),
    .io_reset(regs_356_io_reset),
    .io_out(regs_356_io_out),
    .io_enable(regs_356_io_enable)
  );
  FringeFF regs_357 ( // @[RegFile.scala 66:20:@42627.4]
    .clock(regs_357_clock),
    .reset(regs_357_reset),
    .io_in(regs_357_io_in),
    .io_reset(regs_357_io_reset),
    .io_out(regs_357_io_out),
    .io_enable(regs_357_io_enable)
  );
  FringeFF regs_358 ( // @[RegFile.scala 66:20:@42641.4]
    .clock(regs_358_clock),
    .reset(regs_358_reset),
    .io_in(regs_358_io_in),
    .io_reset(regs_358_io_reset),
    .io_out(regs_358_io_out),
    .io_enable(regs_358_io_enable)
  );
  FringeFF regs_359 ( // @[RegFile.scala 66:20:@42655.4]
    .clock(regs_359_clock),
    .reset(regs_359_reset),
    .io_in(regs_359_io_in),
    .io_reset(regs_359_io_reset),
    .io_out(regs_359_io_out),
    .io_enable(regs_359_io_enable)
  );
  FringeFF regs_360 ( // @[RegFile.scala 66:20:@42669.4]
    .clock(regs_360_clock),
    .reset(regs_360_reset),
    .io_in(regs_360_io_in),
    .io_reset(regs_360_io_reset),
    .io_out(regs_360_io_out),
    .io_enable(regs_360_io_enable)
  );
  FringeFF regs_361 ( // @[RegFile.scala 66:20:@42683.4]
    .clock(regs_361_clock),
    .reset(regs_361_reset),
    .io_in(regs_361_io_in),
    .io_reset(regs_361_io_reset),
    .io_out(regs_361_io_out),
    .io_enable(regs_361_io_enable)
  );
  FringeFF regs_362 ( // @[RegFile.scala 66:20:@42697.4]
    .clock(regs_362_clock),
    .reset(regs_362_reset),
    .io_in(regs_362_io_in),
    .io_reset(regs_362_io_reset),
    .io_out(regs_362_io_out),
    .io_enable(regs_362_io_enable)
  );
  FringeFF regs_363 ( // @[RegFile.scala 66:20:@42711.4]
    .clock(regs_363_clock),
    .reset(regs_363_reset),
    .io_in(regs_363_io_in),
    .io_reset(regs_363_io_reset),
    .io_out(regs_363_io_out),
    .io_enable(regs_363_io_enable)
  );
  FringeFF regs_364 ( // @[RegFile.scala 66:20:@42725.4]
    .clock(regs_364_clock),
    .reset(regs_364_reset),
    .io_in(regs_364_io_in),
    .io_reset(regs_364_io_reset),
    .io_out(regs_364_io_out),
    .io_enable(regs_364_io_enable)
  );
  FringeFF regs_365 ( // @[RegFile.scala 66:20:@42739.4]
    .clock(regs_365_clock),
    .reset(regs_365_reset),
    .io_in(regs_365_io_in),
    .io_reset(regs_365_io_reset),
    .io_out(regs_365_io_out),
    .io_enable(regs_365_io_enable)
  );
  FringeFF regs_366 ( // @[RegFile.scala 66:20:@42753.4]
    .clock(regs_366_clock),
    .reset(regs_366_reset),
    .io_in(regs_366_io_in),
    .io_reset(regs_366_io_reset),
    .io_out(regs_366_io_out),
    .io_enable(regs_366_io_enable)
  );
  FringeFF regs_367 ( // @[RegFile.scala 66:20:@42767.4]
    .clock(regs_367_clock),
    .reset(regs_367_reset),
    .io_in(regs_367_io_in),
    .io_reset(regs_367_io_reset),
    .io_out(regs_367_io_out),
    .io_enable(regs_367_io_enable)
  );
  FringeFF regs_368 ( // @[RegFile.scala 66:20:@42781.4]
    .clock(regs_368_clock),
    .reset(regs_368_reset),
    .io_in(regs_368_io_in),
    .io_reset(regs_368_io_reset),
    .io_out(regs_368_io_out),
    .io_enable(regs_368_io_enable)
  );
  FringeFF regs_369 ( // @[RegFile.scala 66:20:@42795.4]
    .clock(regs_369_clock),
    .reset(regs_369_reset),
    .io_in(regs_369_io_in),
    .io_reset(regs_369_io_reset),
    .io_out(regs_369_io_out),
    .io_enable(regs_369_io_enable)
  );
  FringeFF regs_370 ( // @[RegFile.scala 66:20:@42809.4]
    .clock(regs_370_clock),
    .reset(regs_370_reset),
    .io_in(regs_370_io_in),
    .io_reset(regs_370_io_reset),
    .io_out(regs_370_io_out),
    .io_enable(regs_370_io_enable)
  );
  FringeFF regs_371 ( // @[RegFile.scala 66:20:@42823.4]
    .clock(regs_371_clock),
    .reset(regs_371_reset),
    .io_in(regs_371_io_in),
    .io_reset(regs_371_io_reset),
    .io_out(regs_371_io_out),
    .io_enable(regs_371_io_enable)
  );
  FringeFF regs_372 ( // @[RegFile.scala 66:20:@42837.4]
    .clock(regs_372_clock),
    .reset(regs_372_reset),
    .io_in(regs_372_io_in),
    .io_reset(regs_372_io_reset),
    .io_out(regs_372_io_out),
    .io_enable(regs_372_io_enable)
  );
  FringeFF regs_373 ( // @[RegFile.scala 66:20:@42851.4]
    .clock(regs_373_clock),
    .reset(regs_373_reset),
    .io_in(regs_373_io_in),
    .io_reset(regs_373_io_reset),
    .io_out(regs_373_io_out),
    .io_enable(regs_373_io_enable)
  );
  FringeFF regs_374 ( // @[RegFile.scala 66:20:@42865.4]
    .clock(regs_374_clock),
    .reset(regs_374_reset),
    .io_in(regs_374_io_in),
    .io_reset(regs_374_io_reset),
    .io_out(regs_374_io_out),
    .io_enable(regs_374_io_enable)
  );
  FringeFF regs_375 ( // @[RegFile.scala 66:20:@42879.4]
    .clock(regs_375_clock),
    .reset(regs_375_reset),
    .io_in(regs_375_io_in),
    .io_reset(regs_375_io_reset),
    .io_out(regs_375_io_out),
    .io_enable(regs_375_io_enable)
  );
  FringeFF regs_376 ( // @[RegFile.scala 66:20:@42893.4]
    .clock(regs_376_clock),
    .reset(regs_376_reset),
    .io_in(regs_376_io_in),
    .io_reset(regs_376_io_reset),
    .io_out(regs_376_io_out),
    .io_enable(regs_376_io_enable)
  );
  FringeFF regs_377 ( // @[RegFile.scala 66:20:@42907.4]
    .clock(regs_377_clock),
    .reset(regs_377_reset),
    .io_in(regs_377_io_in),
    .io_reset(regs_377_io_reset),
    .io_out(regs_377_io_out),
    .io_enable(regs_377_io_enable)
  );
  FringeFF regs_378 ( // @[RegFile.scala 66:20:@42921.4]
    .clock(regs_378_clock),
    .reset(regs_378_reset),
    .io_in(regs_378_io_in),
    .io_reset(regs_378_io_reset),
    .io_out(regs_378_io_out),
    .io_enable(regs_378_io_enable)
  );
  FringeFF regs_379 ( // @[RegFile.scala 66:20:@42935.4]
    .clock(regs_379_clock),
    .reset(regs_379_reset),
    .io_in(regs_379_io_in),
    .io_reset(regs_379_io_reset),
    .io_out(regs_379_io_out),
    .io_enable(regs_379_io_enable)
  );
  FringeFF regs_380 ( // @[RegFile.scala 66:20:@42949.4]
    .clock(regs_380_clock),
    .reset(regs_380_reset),
    .io_in(regs_380_io_in),
    .io_reset(regs_380_io_reset),
    .io_out(regs_380_io_out),
    .io_enable(regs_380_io_enable)
  );
  FringeFF regs_381 ( // @[RegFile.scala 66:20:@42963.4]
    .clock(regs_381_clock),
    .reset(regs_381_reset),
    .io_in(regs_381_io_in),
    .io_reset(regs_381_io_reset),
    .io_out(regs_381_io_out),
    .io_enable(regs_381_io_enable)
  );
  FringeFF regs_382 ( // @[RegFile.scala 66:20:@42977.4]
    .clock(regs_382_clock),
    .reset(regs_382_reset),
    .io_in(regs_382_io_in),
    .io_reset(regs_382_io_reset),
    .io_out(regs_382_io_out),
    .io_enable(regs_382_io_enable)
  );
  FringeFF regs_383 ( // @[RegFile.scala 66:20:@42991.4]
    .clock(regs_383_clock),
    .reset(regs_383_reset),
    .io_in(regs_383_io_in),
    .io_reset(regs_383_io_reset),
    .io_out(regs_383_io_out),
    .io_enable(regs_383_io_enable)
  );
  FringeFF regs_384 ( // @[RegFile.scala 66:20:@43005.4]
    .clock(regs_384_clock),
    .reset(regs_384_reset),
    .io_in(regs_384_io_in),
    .io_reset(regs_384_io_reset),
    .io_out(regs_384_io_out),
    .io_enable(regs_384_io_enable)
  );
  FringeFF regs_385 ( // @[RegFile.scala 66:20:@43019.4]
    .clock(regs_385_clock),
    .reset(regs_385_reset),
    .io_in(regs_385_io_in),
    .io_reset(regs_385_io_reset),
    .io_out(regs_385_io_out),
    .io_enable(regs_385_io_enable)
  );
  FringeFF regs_386 ( // @[RegFile.scala 66:20:@43033.4]
    .clock(regs_386_clock),
    .reset(regs_386_reset),
    .io_in(regs_386_io_in),
    .io_reset(regs_386_io_reset),
    .io_out(regs_386_io_out),
    .io_enable(regs_386_io_enable)
  );
  FringeFF regs_387 ( // @[RegFile.scala 66:20:@43047.4]
    .clock(regs_387_clock),
    .reset(regs_387_reset),
    .io_in(regs_387_io_in),
    .io_reset(regs_387_io_reset),
    .io_out(regs_387_io_out),
    .io_enable(regs_387_io_enable)
  );
  FringeFF regs_388 ( // @[RegFile.scala 66:20:@43061.4]
    .clock(regs_388_clock),
    .reset(regs_388_reset),
    .io_in(regs_388_io_in),
    .io_reset(regs_388_io_reset),
    .io_out(regs_388_io_out),
    .io_enable(regs_388_io_enable)
  );
  FringeFF regs_389 ( // @[RegFile.scala 66:20:@43075.4]
    .clock(regs_389_clock),
    .reset(regs_389_reset),
    .io_in(regs_389_io_in),
    .io_reset(regs_389_io_reset),
    .io_out(regs_389_io_out),
    .io_enable(regs_389_io_enable)
  );
  FringeFF regs_390 ( // @[RegFile.scala 66:20:@43089.4]
    .clock(regs_390_clock),
    .reset(regs_390_reset),
    .io_in(regs_390_io_in),
    .io_reset(regs_390_io_reset),
    .io_out(regs_390_io_out),
    .io_enable(regs_390_io_enable)
  );
  FringeFF regs_391 ( // @[RegFile.scala 66:20:@43103.4]
    .clock(regs_391_clock),
    .reset(regs_391_reset),
    .io_in(regs_391_io_in),
    .io_reset(regs_391_io_reset),
    .io_out(regs_391_io_out),
    .io_enable(regs_391_io_enable)
  );
  FringeFF regs_392 ( // @[RegFile.scala 66:20:@43117.4]
    .clock(regs_392_clock),
    .reset(regs_392_reset),
    .io_in(regs_392_io_in),
    .io_reset(regs_392_io_reset),
    .io_out(regs_392_io_out),
    .io_enable(regs_392_io_enable)
  );
  FringeFF regs_393 ( // @[RegFile.scala 66:20:@43131.4]
    .clock(regs_393_clock),
    .reset(regs_393_reset),
    .io_in(regs_393_io_in),
    .io_reset(regs_393_io_reset),
    .io_out(regs_393_io_out),
    .io_enable(regs_393_io_enable)
  );
  FringeFF regs_394 ( // @[RegFile.scala 66:20:@43145.4]
    .clock(regs_394_clock),
    .reset(regs_394_reset),
    .io_in(regs_394_io_in),
    .io_reset(regs_394_io_reset),
    .io_out(regs_394_io_out),
    .io_enable(regs_394_io_enable)
  );
  FringeFF regs_395 ( // @[RegFile.scala 66:20:@43159.4]
    .clock(regs_395_clock),
    .reset(regs_395_reset),
    .io_in(regs_395_io_in),
    .io_reset(regs_395_io_reset),
    .io_out(regs_395_io_out),
    .io_enable(regs_395_io_enable)
  );
  FringeFF regs_396 ( // @[RegFile.scala 66:20:@43173.4]
    .clock(regs_396_clock),
    .reset(regs_396_reset),
    .io_in(regs_396_io_in),
    .io_reset(regs_396_io_reset),
    .io_out(regs_396_io_out),
    .io_enable(regs_396_io_enable)
  );
  FringeFF regs_397 ( // @[RegFile.scala 66:20:@43187.4]
    .clock(regs_397_clock),
    .reset(regs_397_reset),
    .io_in(regs_397_io_in),
    .io_reset(regs_397_io_reset),
    .io_out(regs_397_io_out),
    .io_enable(regs_397_io_enable)
  );
  FringeFF regs_398 ( // @[RegFile.scala 66:20:@43201.4]
    .clock(regs_398_clock),
    .reset(regs_398_reset),
    .io_in(regs_398_io_in),
    .io_reset(regs_398_io_reset),
    .io_out(regs_398_io_out),
    .io_enable(regs_398_io_enable)
  );
  FringeFF regs_399 ( // @[RegFile.scala 66:20:@43215.4]
    .clock(regs_399_clock),
    .reset(regs_399_reset),
    .io_in(regs_399_io_in),
    .io_reset(regs_399_io_reset),
    .io_out(regs_399_io_out),
    .io_enable(regs_399_io_enable)
  );
  FringeFF regs_400 ( // @[RegFile.scala 66:20:@43229.4]
    .clock(regs_400_clock),
    .reset(regs_400_reset),
    .io_in(regs_400_io_in),
    .io_reset(regs_400_io_reset),
    .io_out(regs_400_io_out),
    .io_enable(regs_400_io_enable)
  );
  FringeFF regs_401 ( // @[RegFile.scala 66:20:@43243.4]
    .clock(regs_401_clock),
    .reset(regs_401_reset),
    .io_in(regs_401_io_in),
    .io_reset(regs_401_io_reset),
    .io_out(regs_401_io_out),
    .io_enable(regs_401_io_enable)
  );
  FringeFF regs_402 ( // @[RegFile.scala 66:20:@43257.4]
    .clock(regs_402_clock),
    .reset(regs_402_reset),
    .io_in(regs_402_io_in),
    .io_reset(regs_402_io_reset),
    .io_out(regs_402_io_out),
    .io_enable(regs_402_io_enable)
  );
  FringeFF regs_403 ( // @[RegFile.scala 66:20:@43271.4]
    .clock(regs_403_clock),
    .reset(regs_403_reset),
    .io_in(regs_403_io_in),
    .io_reset(regs_403_io_reset),
    .io_out(regs_403_io_out),
    .io_enable(regs_403_io_enable)
  );
  FringeFF regs_404 ( // @[RegFile.scala 66:20:@43285.4]
    .clock(regs_404_clock),
    .reset(regs_404_reset),
    .io_in(regs_404_io_in),
    .io_reset(regs_404_io_reset),
    .io_out(regs_404_io_out),
    .io_enable(regs_404_io_enable)
  );
  FringeFF regs_405 ( // @[RegFile.scala 66:20:@43299.4]
    .clock(regs_405_clock),
    .reset(regs_405_reset),
    .io_in(regs_405_io_in),
    .io_reset(regs_405_io_reset),
    .io_out(regs_405_io_out),
    .io_enable(regs_405_io_enable)
  );
  FringeFF regs_406 ( // @[RegFile.scala 66:20:@43313.4]
    .clock(regs_406_clock),
    .reset(regs_406_reset),
    .io_in(regs_406_io_in),
    .io_reset(regs_406_io_reset),
    .io_out(regs_406_io_out),
    .io_enable(regs_406_io_enable)
  );
  FringeFF regs_407 ( // @[RegFile.scala 66:20:@43327.4]
    .clock(regs_407_clock),
    .reset(regs_407_reset),
    .io_in(regs_407_io_in),
    .io_reset(regs_407_io_reset),
    .io_out(regs_407_io_out),
    .io_enable(regs_407_io_enable)
  );
  FringeFF regs_408 ( // @[RegFile.scala 66:20:@43341.4]
    .clock(regs_408_clock),
    .reset(regs_408_reset),
    .io_in(regs_408_io_in),
    .io_reset(regs_408_io_reset),
    .io_out(regs_408_io_out),
    .io_enable(regs_408_io_enable)
  );
  FringeFF regs_409 ( // @[RegFile.scala 66:20:@43355.4]
    .clock(regs_409_clock),
    .reset(regs_409_reset),
    .io_in(regs_409_io_in),
    .io_reset(regs_409_io_reset),
    .io_out(regs_409_io_out),
    .io_enable(regs_409_io_enable)
  );
  FringeFF regs_410 ( // @[RegFile.scala 66:20:@43369.4]
    .clock(regs_410_clock),
    .reset(regs_410_reset),
    .io_in(regs_410_io_in),
    .io_reset(regs_410_io_reset),
    .io_out(regs_410_io_out),
    .io_enable(regs_410_io_enable)
  );
  FringeFF regs_411 ( // @[RegFile.scala 66:20:@43383.4]
    .clock(regs_411_clock),
    .reset(regs_411_reset),
    .io_in(regs_411_io_in),
    .io_reset(regs_411_io_reset),
    .io_out(regs_411_io_out),
    .io_enable(regs_411_io_enable)
  );
  FringeFF regs_412 ( // @[RegFile.scala 66:20:@43397.4]
    .clock(regs_412_clock),
    .reset(regs_412_reset),
    .io_in(regs_412_io_in),
    .io_reset(regs_412_io_reset),
    .io_out(regs_412_io_out),
    .io_enable(regs_412_io_enable)
  );
  FringeFF regs_413 ( // @[RegFile.scala 66:20:@43411.4]
    .clock(regs_413_clock),
    .reset(regs_413_reset),
    .io_in(regs_413_io_in),
    .io_reset(regs_413_io_reset),
    .io_out(regs_413_io_out),
    .io_enable(regs_413_io_enable)
  );
  FringeFF regs_414 ( // @[RegFile.scala 66:20:@43425.4]
    .clock(regs_414_clock),
    .reset(regs_414_reset),
    .io_in(regs_414_io_in),
    .io_reset(regs_414_io_reset),
    .io_out(regs_414_io_out),
    .io_enable(regs_414_io_enable)
  );
  FringeFF regs_415 ( // @[RegFile.scala 66:20:@43439.4]
    .clock(regs_415_clock),
    .reset(regs_415_reset),
    .io_in(regs_415_io_in),
    .io_reset(regs_415_io_reset),
    .io_out(regs_415_io_out),
    .io_enable(regs_415_io_enable)
  );
  FringeFF regs_416 ( // @[RegFile.scala 66:20:@43453.4]
    .clock(regs_416_clock),
    .reset(regs_416_reset),
    .io_in(regs_416_io_in),
    .io_reset(regs_416_io_reset),
    .io_out(regs_416_io_out),
    .io_enable(regs_416_io_enable)
  );
  FringeFF regs_417 ( // @[RegFile.scala 66:20:@43467.4]
    .clock(regs_417_clock),
    .reset(regs_417_reset),
    .io_in(regs_417_io_in),
    .io_reset(regs_417_io_reset),
    .io_out(regs_417_io_out),
    .io_enable(regs_417_io_enable)
  );
  FringeFF regs_418 ( // @[RegFile.scala 66:20:@43481.4]
    .clock(regs_418_clock),
    .reset(regs_418_reset),
    .io_in(regs_418_io_in),
    .io_reset(regs_418_io_reset),
    .io_out(regs_418_io_out),
    .io_enable(regs_418_io_enable)
  );
  FringeFF regs_419 ( // @[RegFile.scala 66:20:@43495.4]
    .clock(regs_419_clock),
    .reset(regs_419_reset),
    .io_in(regs_419_io_in),
    .io_reset(regs_419_io_reset),
    .io_out(regs_419_io_out),
    .io_enable(regs_419_io_enable)
  );
  FringeFF regs_420 ( // @[RegFile.scala 66:20:@43509.4]
    .clock(regs_420_clock),
    .reset(regs_420_reset),
    .io_in(regs_420_io_in),
    .io_reset(regs_420_io_reset),
    .io_out(regs_420_io_out),
    .io_enable(regs_420_io_enable)
  );
  FringeFF regs_421 ( // @[RegFile.scala 66:20:@43523.4]
    .clock(regs_421_clock),
    .reset(regs_421_reset),
    .io_in(regs_421_io_in),
    .io_reset(regs_421_io_reset),
    .io_out(regs_421_io_out),
    .io_enable(regs_421_io_enable)
  );
  FringeFF regs_422 ( // @[RegFile.scala 66:20:@43537.4]
    .clock(regs_422_clock),
    .reset(regs_422_reset),
    .io_in(regs_422_io_in),
    .io_reset(regs_422_io_reset),
    .io_out(regs_422_io_out),
    .io_enable(regs_422_io_enable)
  );
  FringeFF regs_423 ( // @[RegFile.scala 66:20:@43551.4]
    .clock(regs_423_clock),
    .reset(regs_423_reset),
    .io_in(regs_423_io_in),
    .io_reset(regs_423_io_reset),
    .io_out(regs_423_io_out),
    .io_enable(regs_423_io_enable)
  );
  FringeFF regs_424 ( // @[RegFile.scala 66:20:@43565.4]
    .clock(regs_424_clock),
    .reset(regs_424_reset),
    .io_in(regs_424_io_in),
    .io_reset(regs_424_io_reset),
    .io_out(regs_424_io_out),
    .io_enable(regs_424_io_enable)
  );
  FringeFF regs_425 ( // @[RegFile.scala 66:20:@43579.4]
    .clock(regs_425_clock),
    .reset(regs_425_reset),
    .io_in(regs_425_io_in),
    .io_reset(regs_425_io_reset),
    .io_out(regs_425_io_out),
    .io_enable(regs_425_io_enable)
  );
  FringeFF regs_426 ( // @[RegFile.scala 66:20:@43593.4]
    .clock(regs_426_clock),
    .reset(regs_426_reset),
    .io_in(regs_426_io_in),
    .io_reset(regs_426_io_reset),
    .io_out(regs_426_io_out),
    .io_enable(regs_426_io_enable)
  );
  FringeFF regs_427 ( // @[RegFile.scala 66:20:@43607.4]
    .clock(regs_427_clock),
    .reset(regs_427_reset),
    .io_in(regs_427_io_in),
    .io_reset(regs_427_io_reset),
    .io_out(regs_427_io_out),
    .io_enable(regs_427_io_enable)
  );
  FringeFF regs_428 ( // @[RegFile.scala 66:20:@43621.4]
    .clock(regs_428_clock),
    .reset(regs_428_reset),
    .io_in(regs_428_io_in),
    .io_reset(regs_428_io_reset),
    .io_out(regs_428_io_out),
    .io_enable(regs_428_io_enable)
  );
  FringeFF regs_429 ( // @[RegFile.scala 66:20:@43635.4]
    .clock(regs_429_clock),
    .reset(regs_429_reset),
    .io_in(regs_429_io_in),
    .io_reset(regs_429_io_reset),
    .io_out(regs_429_io_out),
    .io_enable(regs_429_io_enable)
  );
  FringeFF regs_430 ( // @[RegFile.scala 66:20:@43649.4]
    .clock(regs_430_clock),
    .reset(regs_430_reset),
    .io_in(regs_430_io_in),
    .io_reset(regs_430_io_reset),
    .io_out(regs_430_io_out),
    .io_enable(regs_430_io_enable)
  );
  FringeFF regs_431 ( // @[RegFile.scala 66:20:@43663.4]
    .clock(regs_431_clock),
    .reset(regs_431_reset),
    .io_in(regs_431_io_in),
    .io_reset(regs_431_io_reset),
    .io_out(regs_431_io_out),
    .io_enable(regs_431_io_enable)
  );
  FringeFF regs_432 ( // @[RegFile.scala 66:20:@43677.4]
    .clock(regs_432_clock),
    .reset(regs_432_reset),
    .io_in(regs_432_io_in),
    .io_reset(regs_432_io_reset),
    .io_out(regs_432_io_out),
    .io_enable(regs_432_io_enable)
  );
  FringeFF regs_433 ( // @[RegFile.scala 66:20:@43691.4]
    .clock(regs_433_clock),
    .reset(regs_433_reset),
    .io_in(regs_433_io_in),
    .io_reset(regs_433_io_reset),
    .io_out(regs_433_io_out),
    .io_enable(regs_433_io_enable)
  );
  FringeFF regs_434 ( // @[RegFile.scala 66:20:@43705.4]
    .clock(regs_434_clock),
    .reset(regs_434_reset),
    .io_in(regs_434_io_in),
    .io_reset(regs_434_io_reset),
    .io_out(regs_434_io_out),
    .io_enable(regs_434_io_enable)
  );
  FringeFF regs_435 ( // @[RegFile.scala 66:20:@43719.4]
    .clock(regs_435_clock),
    .reset(regs_435_reset),
    .io_in(regs_435_io_in),
    .io_reset(regs_435_io_reset),
    .io_out(regs_435_io_out),
    .io_enable(regs_435_io_enable)
  );
  FringeFF regs_436 ( // @[RegFile.scala 66:20:@43733.4]
    .clock(regs_436_clock),
    .reset(regs_436_reset),
    .io_in(regs_436_io_in),
    .io_reset(regs_436_io_reset),
    .io_out(regs_436_io_out),
    .io_enable(regs_436_io_enable)
  );
  FringeFF regs_437 ( // @[RegFile.scala 66:20:@43747.4]
    .clock(regs_437_clock),
    .reset(regs_437_reset),
    .io_in(regs_437_io_in),
    .io_reset(regs_437_io_reset),
    .io_out(regs_437_io_out),
    .io_enable(regs_437_io_enable)
  );
  FringeFF regs_438 ( // @[RegFile.scala 66:20:@43761.4]
    .clock(regs_438_clock),
    .reset(regs_438_reset),
    .io_in(regs_438_io_in),
    .io_reset(regs_438_io_reset),
    .io_out(regs_438_io_out),
    .io_enable(regs_438_io_enable)
  );
  FringeFF regs_439 ( // @[RegFile.scala 66:20:@43775.4]
    .clock(regs_439_clock),
    .reset(regs_439_reset),
    .io_in(regs_439_io_in),
    .io_reset(regs_439_io_reset),
    .io_out(regs_439_io_out),
    .io_enable(regs_439_io_enable)
  );
  FringeFF regs_440 ( // @[RegFile.scala 66:20:@43789.4]
    .clock(regs_440_clock),
    .reset(regs_440_reset),
    .io_in(regs_440_io_in),
    .io_reset(regs_440_io_reset),
    .io_out(regs_440_io_out),
    .io_enable(regs_440_io_enable)
  );
  FringeFF regs_441 ( // @[RegFile.scala 66:20:@43803.4]
    .clock(regs_441_clock),
    .reset(regs_441_reset),
    .io_in(regs_441_io_in),
    .io_reset(regs_441_io_reset),
    .io_out(regs_441_io_out),
    .io_enable(regs_441_io_enable)
  );
  FringeFF regs_442 ( // @[RegFile.scala 66:20:@43817.4]
    .clock(regs_442_clock),
    .reset(regs_442_reset),
    .io_in(regs_442_io_in),
    .io_reset(regs_442_io_reset),
    .io_out(regs_442_io_out),
    .io_enable(regs_442_io_enable)
  );
  FringeFF regs_443 ( // @[RegFile.scala 66:20:@43831.4]
    .clock(regs_443_clock),
    .reset(regs_443_reset),
    .io_in(regs_443_io_in),
    .io_reset(regs_443_io_reset),
    .io_out(regs_443_io_out),
    .io_enable(regs_443_io_enable)
  );
  FringeFF regs_444 ( // @[RegFile.scala 66:20:@43845.4]
    .clock(regs_444_clock),
    .reset(regs_444_reset),
    .io_in(regs_444_io_in),
    .io_reset(regs_444_io_reset),
    .io_out(regs_444_io_out),
    .io_enable(regs_444_io_enable)
  );
  FringeFF regs_445 ( // @[RegFile.scala 66:20:@43859.4]
    .clock(regs_445_clock),
    .reset(regs_445_reset),
    .io_in(regs_445_io_in),
    .io_reset(regs_445_io_reset),
    .io_out(regs_445_io_out),
    .io_enable(regs_445_io_enable)
  );
  FringeFF regs_446 ( // @[RegFile.scala 66:20:@43873.4]
    .clock(regs_446_clock),
    .reset(regs_446_reset),
    .io_in(regs_446_io_in),
    .io_reset(regs_446_io_reset),
    .io_out(regs_446_io_out),
    .io_enable(regs_446_io_enable)
  );
  FringeFF regs_447 ( // @[RegFile.scala 66:20:@43887.4]
    .clock(regs_447_clock),
    .reset(regs_447_reset),
    .io_in(regs_447_io_in),
    .io_reset(regs_447_io_reset),
    .io_out(regs_447_io_out),
    .io_enable(regs_447_io_enable)
  );
  FringeFF regs_448 ( // @[RegFile.scala 66:20:@43901.4]
    .clock(regs_448_clock),
    .reset(regs_448_reset),
    .io_in(regs_448_io_in),
    .io_reset(regs_448_io_reset),
    .io_out(regs_448_io_out),
    .io_enable(regs_448_io_enable)
  );
  FringeFF regs_449 ( // @[RegFile.scala 66:20:@43915.4]
    .clock(regs_449_clock),
    .reset(regs_449_reset),
    .io_in(regs_449_io_in),
    .io_reset(regs_449_io_reset),
    .io_out(regs_449_io_out),
    .io_enable(regs_449_io_enable)
  );
  FringeFF regs_450 ( // @[RegFile.scala 66:20:@43929.4]
    .clock(regs_450_clock),
    .reset(regs_450_reset),
    .io_in(regs_450_io_in),
    .io_reset(regs_450_io_reset),
    .io_out(regs_450_io_out),
    .io_enable(regs_450_io_enable)
  );
  FringeFF regs_451 ( // @[RegFile.scala 66:20:@43943.4]
    .clock(regs_451_clock),
    .reset(regs_451_reset),
    .io_in(regs_451_io_in),
    .io_reset(regs_451_io_reset),
    .io_out(regs_451_io_out),
    .io_enable(regs_451_io_enable)
  );
  FringeFF regs_452 ( // @[RegFile.scala 66:20:@43957.4]
    .clock(regs_452_clock),
    .reset(regs_452_reset),
    .io_in(regs_452_io_in),
    .io_reset(regs_452_io_reset),
    .io_out(regs_452_io_out),
    .io_enable(regs_452_io_enable)
  );
  FringeFF regs_453 ( // @[RegFile.scala 66:20:@43971.4]
    .clock(regs_453_clock),
    .reset(regs_453_reset),
    .io_in(regs_453_io_in),
    .io_reset(regs_453_io_reset),
    .io_out(regs_453_io_out),
    .io_enable(regs_453_io_enable)
  );
  FringeFF regs_454 ( // @[RegFile.scala 66:20:@43985.4]
    .clock(regs_454_clock),
    .reset(regs_454_reset),
    .io_in(regs_454_io_in),
    .io_reset(regs_454_io_reset),
    .io_out(regs_454_io_out),
    .io_enable(regs_454_io_enable)
  );
  FringeFF regs_455 ( // @[RegFile.scala 66:20:@43999.4]
    .clock(regs_455_clock),
    .reset(regs_455_reset),
    .io_in(regs_455_io_in),
    .io_reset(regs_455_io_reset),
    .io_out(regs_455_io_out),
    .io_enable(regs_455_io_enable)
  );
  FringeFF regs_456 ( // @[RegFile.scala 66:20:@44013.4]
    .clock(regs_456_clock),
    .reset(regs_456_reset),
    .io_in(regs_456_io_in),
    .io_reset(regs_456_io_reset),
    .io_out(regs_456_io_out),
    .io_enable(regs_456_io_enable)
  );
  FringeFF regs_457 ( // @[RegFile.scala 66:20:@44027.4]
    .clock(regs_457_clock),
    .reset(regs_457_reset),
    .io_in(regs_457_io_in),
    .io_reset(regs_457_io_reset),
    .io_out(regs_457_io_out),
    .io_enable(regs_457_io_enable)
  );
  FringeFF regs_458 ( // @[RegFile.scala 66:20:@44041.4]
    .clock(regs_458_clock),
    .reset(regs_458_reset),
    .io_in(regs_458_io_in),
    .io_reset(regs_458_io_reset),
    .io_out(regs_458_io_out),
    .io_enable(regs_458_io_enable)
  );
  FringeFF regs_459 ( // @[RegFile.scala 66:20:@44055.4]
    .clock(regs_459_clock),
    .reset(regs_459_reset),
    .io_in(regs_459_io_in),
    .io_reset(regs_459_io_reset),
    .io_out(regs_459_io_out),
    .io_enable(regs_459_io_enable)
  );
  FringeFF regs_460 ( // @[RegFile.scala 66:20:@44069.4]
    .clock(regs_460_clock),
    .reset(regs_460_reset),
    .io_in(regs_460_io_in),
    .io_reset(regs_460_io_reset),
    .io_out(regs_460_io_out),
    .io_enable(regs_460_io_enable)
  );
  FringeFF regs_461 ( // @[RegFile.scala 66:20:@44083.4]
    .clock(regs_461_clock),
    .reset(regs_461_reset),
    .io_in(regs_461_io_in),
    .io_reset(regs_461_io_reset),
    .io_out(regs_461_io_out),
    .io_enable(regs_461_io_enable)
  );
  FringeFF regs_462 ( // @[RegFile.scala 66:20:@44097.4]
    .clock(regs_462_clock),
    .reset(regs_462_reset),
    .io_in(regs_462_io_in),
    .io_reset(regs_462_io_reset),
    .io_out(regs_462_io_out),
    .io_enable(regs_462_io_enable)
  );
  FringeFF regs_463 ( // @[RegFile.scala 66:20:@44111.4]
    .clock(regs_463_clock),
    .reset(regs_463_reset),
    .io_in(regs_463_io_in),
    .io_reset(regs_463_io_reset),
    .io_out(regs_463_io_out),
    .io_enable(regs_463_io_enable)
  );
  FringeFF regs_464 ( // @[RegFile.scala 66:20:@44125.4]
    .clock(regs_464_clock),
    .reset(regs_464_reset),
    .io_in(regs_464_io_in),
    .io_reset(regs_464_io_reset),
    .io_out(regs_464_io_out),
    .io_enable(regs_464_io_enable)
  );
  FringeFF regs_465 ( // @[RegFile.scala 66:20:@44139.4]
    .clock(regs_465_clock),
    .reset(regs_465_reset),
    .io_in(regs_465_io_in),
    .io_reset(regs_465_io_reset),
    .io_out(regs_465_io_out),
    .io_enable(regs_465_io_enable)
  );
  FringeFF regs_466 ( // @[RegFile.scala 66:20:@44153.4]
    .clock(regs_466_clock),
    .reset(regs_466_reset),
    .io_in(regs_466_io_in),
    .io_reset(regs_466_io_reset),
    .io_out(regs_466_io_out),
    .io_enable(regs_466_io_enable)
  );
  FringeFF regs_467 ( // @[RegFile.scala 66:20:@44167.4]
    .clock(regs_467_clock),
    .reset(regs_467_reset),
    .io_in(regs_467_io_in),
    .io_reset(regs_467_io_reset),
    .io_out(regs_467_io_out),
    .io_enable(regs_467_io_enable)
  );
  FringeFF regs_468 ( // @[RegFile.scala 66:20:@44181.4]
    .clock(regs_468_clock),
    .reset(regs_468_reset),
    .io_in(regs_468_io_in),
    .io_reset(regs_468_io_reset),
    .io_out(regs_468_io_out),
    .io_enable(regs_468_io_enable)
  );
  FringeFF regs_469 ( // @[RegFile.scala 66:20:@44195.4]
    .clock(regs_469_clock),
    .reset(regs_469_reset),
    .io_in(regs_469_io_in),
    .io_reset(regs_469_io_reset),
    .io_out(regs_469_io_out),
    .io_enable(regs_469_io_enable)
  );
  FringeFF regs_470 ( // @[RegFile.scala 66:20:@44209.4]
    .clock(regs_470_clock),
    .reset(regs_470_reset),
    .io_in(regs_470_io_in),
    .io_reset(regs_470_io_reset),
    .io_out(regs_470_io_out),
    .io_enable(regs_470_io_enable)
  );
  FringeFF regs_471 ( // @[RegFile.scala 66:20:@44223.4]
    .clock(regs_471_clock),
    .reset(regs_471_reset),
    .io_in(regs_471_io_in),
    .io_reset(regs_471_io_reset),
    .io_out(regs_471_io_out),
    .io_enable(regs_471_io_enable)
  );
  FringeFF regs_472 ( // @[RegFile.scala 66:20:@44237.4]
    .clock(regs_472_clock),
    .reset(regs_472_reset),
    .io_in(regs_472_io_in),
    .io_reset(regs_472_io_reset),
    .io_out(regs_472_io_out),
    .io_enable(regs_472_io_enable)
  );
  FringeFF regs_473 ( // @[RegFile.scala 66:20:@44251.4]
    .clock(regs_473_clock),
    .reset(regs_473_reset),
    .io_in(regs_473_io_in),
    .io_reset(regs_473_io_reset),
    .io_out(regs_473_io_out),
    .io_enable(regs_473_io_enable)
  );
  FringeFF regs_474 ( // @[RegFile.scala 66:20:@44265.4]
    .clock(regs_474_clock),
    .reset(regs_474_reset),
    .io_in(regs_474_io_in),
    .io_reset(regs_474_io_reset),
    .io_out(regs_474_io_out),
    .io_enable(regs_474_io_enable)
  );
  FringeFF regs_475 ( // @[RegFile.scala 66:20:@44279.4]
    .clock(regs_475_clock),
    .reset(regs_475_reset),
    .io_in(regs_475_io_in),
    .io_reset(regs_475_io_reset),
    .io_out(regs_475_io_out),
    .io_enable(regs_475_io_enable)
  );
  FringeFF regs_476 ( // @[RegFile.scala 66:20:@44293.4]
    .clock(regs_476_clock),
    .reset(regs_476_reset),
    .io_in(regs_476_io_in),
    .io_reset(regs_476_io_reset),
    .io_out(regs_476_io_out),
    .io_enable(regs_476_io_enable)
  );
  FringeFF regs_477 ( // @[RegFile.scala 66:20:@44307.4]
    .clock(regs_477_clock),
    .reset(regs_477_reset),
    .io_in(regs_477_io_in),
    .io_reset(regs_477_io_reset),
    .io_out(regs_477_io_out),
    .io_enable(regs_477_io_enable)
  );
  FringeFF regs_478 ( // @[RegFile.scala 66:20:@44321.4]
    .clock(regs_478_clock),
    .reset(regs_478_reset),
    .io_in(regs_478_io_in),
    .io_reset(regs_478_io_reset),
    .io_out(regs_478_io_out),
    .io_enable(regs_478_io_enable)
  );
  FringeFF regs_479 ( // @[RegFile.scala 66:20:@44335.4]
    .clock(regs_479_clock),
    .reset(regs_479_reset),
    .io_in(regs_479_io_in),
    .io_reset(regs_479_io_reset),
    .io_out(regs_479_io_out),
    .io_enable(regs_479_io_enable)
  );
  FringeFF regs_480 ( // @[RegFile.scala 66:20:@44349.4]
    .clock(regs_480_clock),
    .reset(regs_480_reset),
    .io_in(regs_480_io_in),
    .io_reset(regs_480_io_reset),
    .io_out(regs_480_io_out),
    .io_enable(regs_480_io_enable)
  );
  FringeFF regs_481 ( // @[RegFile.scala 66:20:@44363.4]
    .clock(regs_481_clock),
    .reset(regs_481_reset),
    .io_in(regs_481_io_in),
    .io_reset(regs_481_io_reset),
    .io_out(regs_481_io_out),
    .io_enable(regs_481_io_enable)
  );
  FringeFF regs_482 ( // @[RegFile.scala 66:20:@44377.4]
    .clock(regs_482_clock),
    .reset(regs_482_reset),
    .io_in(regs_482_io_in),
    .io_reset(regs_482_io_reset),
    .io_out(regs_482_io_out),
    .io_enable(regs_482_io_enable)
  );
  FringeFF regs_483 ( // @[RegFile.scala 66:20:@44391.4]
    .clock(regs_483_clock),
    .reset(regs_483_reset),
    .io_in(regs_483_io_in),
    .io_reset(regs_483_io_reset),
    .io_out(regs_483_io_out),
    .io_enable(regs_483_io_enable)
  );
  FringeFF regs_484 ( // @[RegFile.scala 66:20:@44405.4]
    .clock(regs_484_clock),
    .reset(regs_484_reset),
    .io_in(regs_484_io_in),
    .io_reset(regs_484_io_reset),
    .io_out(regs_484_io_out),
    .io_enable(regs_484_io_enable)
  );
  FringeFF regs_485 ( // @[RegFile.scala 66:20:@44419.4]
    .clock(regs_485_clock),
    .reset(regs_485_reset),
    .io_in(regs_485_io_in),
    .io_reset(regs_485_io_reset),
    .io_out(regs_485_io_out),
    .io_enable(regs_485_io_enable)
  );
  FringeFF regs_486 ( // @[RegFile.scala 66:20:@44433.4]
    .clock(regs_486_clock),
    .reset(regs_486_reset),
    .io_in(regs_486_io_in),
    .io_reset(regs_486_io_reset),
    .io_out(regs_486_io_out),
    .io_enable(regs_486_io_enable)
  );
  FringeFF regs_487 ( // @[RegFile.scala 66:20:@44447.4]
    .clock(regs_487_clock),
    .reset(regs_487_reset),
    .io_in(regs_487_io_in),
    .io_reset(regs_487_io_reset),
    .io_out(regs_487_io_out),
    .io_enable(regs_487_io_enable)
  );
  FringeFF regs_488 ( // @[RegFile.scala 66:20:@44461.4]
    .clock(regs_488_clock),
    .reset(regs_488_reset),
    .io_in(regs_488_io_in),
    .io_reset(regs_488_io_reset),
    .io_out(regs_488_io_out),
    .io_enable(regs_488_io_enable)
  );
  FringeFF regs_489 ( // @[RegFile.scala 66:20:@44475.4]
    .clock(regs_489_clock),
    .reset(regs_489_reset),
    .io_in(regs_489_io_in),
    .io_reset(regs_489_io_reset),
    .io_out(regs_489_io_out),
    .io_enable(regs_489_io_enable)
  );
  FringeFF regs_490 ( // @[RegFile.scala 66:20:@44489.4]
    .clock(regs_490_clock),
    .reset(regs_490_reset),
    .io_in(regs_490_io_in),
    .io_reset(regs_490_io_reset),
    .io_out(regs_490_io_out),
    .io_enable(regs_490_io_enable)
  );
  FringeFF regs_491 ( // @[RegFile.scala 66:20:@44503.4]
    .clock(regs_491_clock),
    .reset(regs_491_reset),
    .io_in(regs_491_io_in),
    .io_reset(regs_491_io_reset),
    .io_out(regs_491_io_out),
    .io_enable(regs_491_io_enable)
  );
  FringeFF regs_492 ( // @[RegFile.scala 66:20:@44517.4]
    .clock(regs_492_clock),
    .reset(regs_492_reset),
    .io_in(regs_492_io_in),
    .io_reset(regs_492_io_reset),
    .io_out(regs_492_io_out),
    .io_enable(regs_492_io_enable)
  );
  FringeFF regs_493 ( // @[RegFile.scala 66:20:@44531.4]
    .clock(regs_493_clock),
    .reset(regs_493_reset),
    .io_in(regs_493_io_in),
    .io_reset(regs_493_io_reset),
    .io_out(regs_493_io_out),
    .io_enable(regs_493_io_enable)
  );
  FringeFF regs_494 ( // @[RegFile.scala 66:20:@44545.4]
    .clock(regs_494_clock),
    .reset(regs_494_reset),
    .io_in(regs_494_io_in),
    .io_reset(regs_494_io_reset),
    .io_out(regs_494_io_out),
    .io_enable(regs_494_io_enable)
  );
  FringeFF regs_495 ( // @[RegFile.scala 66:20:@44559.4]
    .clock(regs_495_clock),
    .reset(regs_495_reset),
    .io_in(regs_495_io_in),
    .io_reset(regs_495_io_reset),
    .io_out(regs_495_io_out),
    .io_enable(regs_495_io_enable)
  );
  FringeFF regs_496 ( // @[RegFile.scala 66:20:@44573.4]
    .clock(regs_496_clock),
    .reset(regs_496_reset),
    .io_in(regs_496_io_in),
    .io_reset(regs_496_io_reset),
    .io_out(regs_496_io_out),
    .io_enable(regs_496_io_enable)
  );
  FringeFF regs_497 ( // @[RegFile.scala 66:20:@44587.4]
    .clock(regs_497_clock),
    .reset(regs_497_reset),
    .io_in(regs_497_io_in),
    .io_reset(regs_497_io_reset),
    .io_out(regs_497_io_out),
    .io_enable(regs_497_io_enable)
  );
  FringeFF regs_498 ( // @[RegFile.scala 66:20:@44601.4]
    .clock(regs_498_clock),
    .reset(regs_498_reset),
    .io_in(regs_498_io_in),
    .io_reset(regs_498_io_reset),
    .io_out(regs_498_io_out),
    .io_enable(regs_498_io_enable)
  );
  FringeFF regs_499 ( // @[RegFile.scala 66:20:@44615.4]
    .clock(regs_499_clock),
    .reset(regs_499_reset),
    .io_in(regs_499_io_in),
    .io_reset(regs_499_io_reset),
    .io_out(regs_499_io_out),
    .io_enable(regs_499_io_enable)
  );
  FringeFF regs_500 ( // @[RegFile.scala 66:20:@44629.4]
    .clock(regs_500_clock),
    .reset(regs_500_reset),
    .io_in(regs_500_io_in),
    .io_reset(regs_500_io_reset),
    .io_out(regs_500_io_out),
    .io_enable(regs_500_io_enable)
  );
  FringeFF regs_501 ( // @[RegFile.scala 66:20:@44643.4]
    .clock(regs_501_clock),
    .reset(regs_501_reset),
    .io_in(regs_501_io_in),
    .io_reset(regs_501_io_reset),
    .io_out(regs_501_io_out),
    .io_enable(regs_501_io_enable)
  );
  FringeFF regs_502 ( // @[RegFile.scala 66:20:@44657.4]
    .clock(regs_502_clock),
    .reset(regs_502_reset),
    .io_in(regs_502_io_in),
    .io_reset(regs_502_io_reset),
    .io_out(regs_502_io_out),
    .io_enable(regs_502_io_enable)
  );
  FringeFF regs_503 ( // @[RegFile.scala 66:20:@44671.4]
    .clock(regs_503_clock),
    .reset(regs_503_reset),
    .io_in(regs_503_io_in),
    .io_reset(regs_503_io_reset),
    .io_out(regs_503_io_out),
    .io_enable(regs_503_io_enable)
  );
  FringeFF regs_504 ( // @[RegFile.scala 66:20:@44685.4]
    .clock(regs_504_clock),
    .reset(regs_504_reset),
    .io_in(regs_504_io_in),
    .io_reset(regs_504_io_reset),
    .io_out(regs_504_io_out),
    .io_enable(regs_504_io_enable)
  );
  FringeFF regs_505 ( // @[RegFile.scala 66:20:@44699.4]
    .clock(regs_505_clock),
    .reset(regs_505_reset),
    .io_in(regs_505_io_in),
    .io_reset(regs_505_io_reset),
    .io_out(regs_505_io_out),
    .io_enable(regs_505_io_enable)
  );
  FringeFF regs_506 ( // @[RegFile.scala 66:20:@44713.4]
    .clock(regs_506_clock),
    .reset(regs_506_reset),
    .io_in(regs_506_io_in),
    .io_reset(regs_506_io_reset),
    .io_out(regs_506_io_out),
    .io_enable(regs_506_io_enable)
  );
  FringeFF regs_507 ( // @[RegFile.scala 66:20:@44727.4]
    .clock(regs_507_clock),
    .reset(regs_507_reset),
    .io_in(regs_507_io_in),
    .io_reset(regs_507_io_reset),
    .io_out(regs_507_io_out),
    .io_enable(regs_507_io_enable)
  );
  FringeFF regs_508 ( // @[RegFile.scala 66:20:@44741.4]
    .clock(regs_508_clock),
    .reset(regs_508_reset),
    .io_in(regs_508_io_in),
    .io_reset(regs_508_io_reset),
    .io_out(regs_508_io_out),
    .io_enable(regs_508_io_enable)
  );
  FringeFF regs_509 ( // @[RegFile.scala 66:20:@44755.4]
    .clock(regs_509_clock),
    .reset(regs_509_reset),
    .io_in(regs_509_io_in),
    .io_reset(regs_509_io_reset),
    .io_out(regs_509_io_out),
    .io_enable(regs_509_io_enable)
  );
  FringeFF regs_510 ( // @[RegFile.scala 66:20:@44769.4]
    .clock(regs_510_clock),
    .reset(regs_510_reset),
    .io_in(regs_510_io_in),
    .io_reset(regs_510_io_reset),
    .io_out(regs_510_io_out),
    .io_enable(regs_510_io_enable)
  );
  FringeFF regs_511 ( // @[RegFile.scala 66:20:@44783.4]
    .clock(regs_511_clock),
    .reset(regs_511_reset),
    .io_in(regs_511_io_in),
    .io_reset(regs_511_io_reset),
    .io_out(regs_511_io_out),
    .io_enable(regs_511_io_enable)
  );
  MuxN rport ( // @[RegFile.scala 95:21:@44797.4]
    .io_ins_0(rport_io_ins_0),
    .io_ins_1(rport_io_ins_1),
    .io_ins_2(rport_io_ins_2),
    .io_ins_3(rport_io_ins_3),
    .io_ins_4(rport_io_ins_4),
    .io_ins_5(rport_io_ins_5),
    .io_ins_6(rport_io_ins_6),
    .io_ins_7(rport_io_ins_7),
    .io_ins_8(rport_io_ins_8),
    .io_ins_9(rport_io_ins_9),
    .io_ins_10(rport_io_ins_10),
    .io_ins_11(rport_io_ins_11),
    .io_ins_12(rport_io_ins_12),
    .io_ins_13(rport_io_ins_13),
    .io_ins_14(rport_io_ins_14),
    .io_ins_15(rport_io_ins_15),
    .io_ins_16(rport_io_ins_16),
    .io_ins_17(rport_io_ins_17),
    .io_ins_18(rport_io_ins_18),
    .io_ins_19(rport_io_ins_19),
    .io_ins_20(rport_io_ins_20),
    .io_ins_21(rport_io_ins_21),
    .io_ins_22(rport_io_ins_22),
    .io_ins_23(rport_io_ins_23),
    .io_ins_24(rport_io_ins_24),
    .io_ins_25(rport_io_ins_25),
    .io_ins_26(rport_io_ins_26),
    .io_ins_27(rport_io_ins_27),
    .io_ins_28(rport_io_ins_28),
    .io_ins_29(rport_io_ins_29),
    .io_ins_30(rport_io_ins_30),
    .io_ins_31(rport_io_ins_31),
    .io_ins_32(rport_io_ins_32),
    .io_ins_33(rport_io_ins_33),
    .io_ins_34(rport_io_ins_34),
    .io_ins_35(rport_io_ins_35),
    .io_ins_36(rport_io_ins_36),
    .io_ins_37(rport_io_ins_37),
    .io_ins_38(rport_io_ins_38),
    .io_ins_39(rport_io_ins_39),
    .io_ins_40(rport_io_ins_40),
    .io_ins_41(rport_io_ins_41),
    .io_ins_42(rport_io_ins_42),
    .io_ins_43(rport_io_ins_43),
    .io_ins_44(rport_io_ins_44),
    .io_ins_45(rport_io_ins_45),
    .io_ins_46(rport_io_ins_46),
    .io_ins_47(rport_io_ins_47),
    .io_ins_48(rport_io_ins_48),
    .io_ins_49(rport_io_ins_49),
    .io_ins_50(rport_io_ins_50),
    .io_ins_51(rport_io_ins_51),
    .io_ins_52(rport_io_ins_52),
    .io_ins_53(rport_io_ins_53),
    .io_ins_54(rport_io_ins_54),
    .io_ins_55(rport_io_ins_55),
    .io_ins_56(rport_io_ins_56),
    .io_ins_57(rport_io_ins_57),
    .io_ins_58(rport_io_ins_58),
    .io_ins_59(rport_io_ins_59),
    .io_ins_60(rport_io_ins_60),
    .io_ins_61(rport_io_ins_61),
    .io_ins_62(rport_io_ins_62),
    .io_ins_63(rport_io_ins_63),
    .io_ins_64(rport_io_ins_64),
    .io_ins_65(rport_io_ins_65),
    .io_ins_66(rport_io_ins_66),
    .io_ins_67(rport_io_ins_67),
    .io_ins_68(rport_io_ins_68),
    .io_ins_69(rport_io_ins_69),
    .io_ins_70(rport_io_ins_70),
    .io_ins_71(rport_io_ins_71),
    .io_ins_72(rport_io_ins_72),
    .io_ins_73(rport_io_ins_73),
    .io_ins_74(rport_io_ins_74),
    .io_ins_75(rport_io_ins_75),
    .io_ins_76(rport_io_ins_76),
    .io_ins_77(rport_io_ins_77),
    .io_ins_78(rport_io_ins_78),
    .io_ins_79(rport_io_ins_79),
    .io_ins_80(rport_io_ins_80),
    .io_ins_81(rport_io_ins_81),
    .io_ins_82(rport_io_ins_82),
    .io_ins_83(rport_io_ins_83),
    .io_ins_84(rport_io_ins_84),
    .io_ins_85(rport_io_ins_85),
    .io_ins_86(rport_io_ins_86),
    .io_ins_87(rport_io_ins_87),
    .io_ins_88(rport_io_ins_88),
    .io_ins_89(rport_io_ins_89),
    .io_ins_90(rport_io_ins_90),
    .io_ins_91(rport_io_ins_91),
    .io_ins_92(rport_io_ins_92),
    .io_ins_93(rport_io_ins_93),
    .io_ins_94(rport_io_ins_94),
    .io_ins_95(rport_io_ins_95),
    .io_ins_96(rport_io_ins_96),
    .io_ins_97(rport_io_ins_97),
    .io_ins_98(rport_io_ins_98),
    .io_ins_99(rport_io_ins_99),
    .io_ins_100(rport_io_ins_100),
    .io_ins_101(rport_io_ins_101),
    .io_ins_102(rport_io_ins_102),
    .io_ins_103(rport_io_ins_103),
    .io_ins_104(rport_io_ins_104),
    .io_ins_105(rport_io_ins_105),
    .io_ins_106(rport_io_ins_106),
    .io_ins_107(rport_io_ins_107),
    .io_ins_108(rport_io_ins_108),
    .io_ins_109(rport_io_ins_109),
    .io_ins_110(rport_io_ins_110),
    .io_ins_111(rport_io_ins_111),
    .io_ins_112(rport_io_ins_112),
    .io_ins_113(rport_io_ins_113),
    .io_ins_114(rport_io_ins_114),
    .io_ins_115(rport_io_ins_115),
    .io_ins_116(rport_io_ins_116),
    .io_ins_117(rport_io_ins_117),
    .io_ins_118(rport_io_ins_118),
    .io_ins_119(rport_io_ins_119),
    .io_ins_120(rport_io_ins_120),
    .io_ins_121(rport_io_ins_121),
    .io_ins_122(rport_io_ins_122),
    .io_ins_123(rport_io_ins_123),
    .io_ins_124(rport_io_ins_124),
    .io_ins_125(rport_io_ins_125),
    .io_ins_126(rport_io_ins_126),
    .io_ins_127(rport_io_ins_127),
    .io_ins_128(rport_io_ins_128),
    .io_ins_129(rport_io_ins_129),
    .io_ins_130(rport_io_ins_130),
    .io_ins_131(rport_io_ins_131),
    .io_ins_132(rport_io_ins_132),
    .io_ins_133(rport_io_ins_133),
    .io_ins_134(rport_io_ins_134),
    .io_ins_135(rport_io_ins_135),
    .io_ins_136(rport_io_ins_136),
    .io_ins_137(rport_io_ins_137),
    .io_ins_138(rport_io_ins_138),
    .io_ins_139(rport_io_ins_139),
    .io_ins_140(rport_io_ins_140),
    .io_ins_141(rport_io_ins_141),
    .io_ins_142(rport_io_ins_142),
    .io_ins_143(rport_io_ins_143),
    .io_ins_144(rport_io_ins_144),
    .io_ins_145(rport_io_ins_145),
    .io_ins_146(rport_io_ins_146),
    .io_ins_147(rport_io_ins_147),
    .io_ins_148(rport_io_ins_148),
    .io_ins_149(rport_io_ins_149),
    .io_ins_150(rport_io_ins_150),
    .io_ins_151(rport_io_ins_151),
    .io_ins_152(rport_io_ins_152),
    .io_ins_153(rport_io_ins_153),
    .io_ins_154(rport_io_ins_154),
    .io_ins_155(rport_io_ins_155),
    .io_ins_156(rport_io_ins_156),
    .io_ins_157(rport_io_ins_157),
    .io_ins_158(rport_io_ins_158),
    .io_ins_159(rport_io_ins_159),
    .io_ins_160(rport_io_ins_160),
    .io_ins_161(rport_io_ins_161),
    .io_ins_162(rport_io_ins_162),
    .io_ins_163(rport_io_ins_163),
    .io_ins_164(rport_io_ins_164),
    .io_ins_165(rport_io_ins_165),
    .io_ins_166(rport_io_ins_166),
    .io_ins_167(rport_io_ins_167),
    .io_ins_168(rport_io_ins_168),
    .io_ins_169(rport_io_ins_169),
    .io_ins_170(rport_io_ins_170),
    .io_ins_171(rport_io_ins_171),
    .io_ins_172(rport_io_ins_172),
    .io_ins_173(rport_io_ins_173),
    .io_ins_174(rport_io_ins_174),
    .io_ins_175(rport_io_ins_175),
    .io_ins_176(rport_io_ins_176),
    .io_ins_177(rport_io_ins_177),
    .io_ins_178(rport_io_ins_178),
    .io_ins_179(rport_io_ins_179),
    .io_ins_180(rport_io_ins_180),
    .io_ins_181(rport_io_ins_181),
    .io_ins_182(rport_io_ins_182),
    .io_ins_183(rport_io_ins_183),
    .io_ins_184(rport_io_ins_184),
    .io_ins_185(rport_io_ins_185),
    .io_ins_186(rport_io_ins_186),
    .io_ins_187(rport_io_ins_187),
    .io_ins_188(rport_io_ins_188),
    .io_ins_189(rport_io_ins_189),
    .io_ins_190(rport_io_ins_190),
    .io_ins_191(rport_io_ins_191),
    .io_ins_192(rport_io_ins_192),
    .io_ins_193(rport_io_ins_193),
    .io_ins_194(rport_io_ins_194),
    .io_ins_195(rport_io_ins_195),
    .io_ins_196(rport_io_ins_196),
    .io_ins_197(rport_io_ins_197),
    .io_ins_198(rport_io_ins_198),
    .io_ins_199(rport_io_ins_199),
    .io_ins_200(rport_io_ins_200),
    .io_ins_201(rport_io_ins_201),
    .io_ins_202(rport_io_ins_202),
    .io_ins_203(rport_io_ins_203),
    .io_ins_204(rport_io_ins_204),
    .io_ins_205(rport_io_ins_205),
    .io_ins_206(rport_io_ins_206),
    .io_ins_207(rport_io_ins_207),
    .io_ins_208(rport_io_ins_208),
    .io_ins_209(rport_io_ins_209),
    .io_ins_210(rport_io_ins_210),
    .io_ins_211(rport_io_ins_211),
    .io_ins_212(rport_io_ins_212),
    .io_ins_213(rport_io_ins_213),
    .io_ins_214(rport_io_ins_214),
    .io_ins_215(rport_io_ins_215),
    .io_ins_216(rport_io_ins_216),
    .io_ins_217(rport_io_ins_217),
    .io_ins_218(rport_io_ins_218),
    .io_ins_219(rport_io_ins_219),
    .io_ins_220(rport_io_ins_220),
    .io_ins_221(rport_io_ins_221),
    .io_ins_222(rport_io_ins_222),
    .io_ins_223(rport_io_ins_223),
    .io_ins_224(rport_io_ins_224),
    .io_ins_225(rport_io_ins_225),
    .io_ins_226(rport_io_ins_226),
    .io_ins_227(rport_io_ins_227),
    .io_ins_228(rport_io_ins_228),
    .io_ins_229(rport_io_ins_229),
    .io_ins_230(rport_io_ins_230),
    .io_ins_231(rport_io_ins_231),
    .io_ins_232(rport_io_ins_232),
    .io_ins_233(rport_io_ins_233),
    .io_ins_234(rport_io_ins_234),
    .io_ins_235(rport_io_ins_235),
    .io_ins_236(rport_io_ins_236),
    .io_ins_237(rport_io_ins_237),
    .io_ins_238(rport_io_ins_238),
    .io_ins_239(rport_io_ins_239),
    .io_ins_240(rport_io_ins_240),
    .io_ins_241(rport_io_ins_241),
    .io_ins_242(rport_io_ins_242),
    .io_ins_243(rport_io_ins_243),
    .io_ins_244(rport_io_ins_244),
    .io_ins_245(rport_io_ins_245),
    .io_ins_246(rport_io_ins_246),
    .io_ins_247(rport_io_ins_247),
    .io_ins_248(rport_io_ins_248),
    .io_ins_249(rport_io_ins_249),
    .io_ins_250(rport_io_ins_250),
    .io_ins_251(rport_io_ins_251),
    .io_ins_252(rport_io_ins_252),
    .io_ins_253(rport_io_ins_253),
    .io_ins_254(rport_io_ins_254),
    .io_ins_255(rport_io_ins_255),
    .io_ins_256(rport_io_ins_256),
    .io_ins_257(rport_io_ins_257),
    .io_ins_258(rport_io_ins_258),
    .io_ins_259(rport_io_ins_259),
    .io_ins_260(rport_io_ins_260),
    .io_ins_261(rport_io_ins_261),
    .io_ins_262(rport_io_ins_262),
    .io_ins_263(rport_io_ins_263),
    .io_ins_264(rport_io_ins_264),
    .io_ins_265(rport_io_ins_265),
    .io_ins_266(rport_io_ins_266),
    .io_ins_267(rport_io_ins_267),
    .io_ins_268(rport_io_ins_268),
    .io_ins_269(rport_io_ins_269),
    .io_ins_270(rport_io_ins_270),
    .io_ins_271(rport_io_ins_271),
    .io_ins_272(rport_io_ins_272),
    .io_ins_273(rport_io_ins_273),
    .io_ins_274(rport_io_ins_274),
    .io_ins_275(rport_io_ins_275),
    .io_ins_276(rport_io_ins_276),
    .io_ins_277(rport_io_ins_277),
    .io_ins_278(rport_io_ins_278),
    .io_ins_279(rport_io_ins_279),
    .io_ins_280(rport_io_ins_280),
    .io_ins_281(rport_io_ins_281),
    .io_ins_282(rport_io_ins_282),
    .io_ins_283(rport_io_ins_283),
    .io_ins_284(rport_io_ins_284),
    .io_ins_285(rport_io_ins_285),
    .io_ins_286(rport_io_ins_286),
    .io_ins_287(rport_io_ins_287),
    .io_ins_288(rport_io_ins_288),
    .io_ins_289(rport_io_ins_289),
    .io_ins_290(rport_io_ins_290),
    .io_ins_291(rport_io_ins_291),
    .io_ins_292(rport_io_ins_292),
    .io_ins_293(rport_io_ins_293),
    .io_ins_294(rport_io_ins_294),
    .io_ins_295(rport_io_ins_295),
    .io_ins_296(rport_io_ins_296),
    .io_ins_297(rport_io_ins_297),
    .io_ins_298(rport_io_ins_298),
    .io_ins_299(rport_io_ins_299),
    .io_ins_300(rport_io_ins_300),
    .io_ins_301(rport_io_ins_301),
    .io_ins_302(rport_io_ins_302),
    .io_ins_303(rport_io_ins_303),
    .io_ins_304(rport_io_ins_304),
    .io_ins_305(rport_io_ins_305),
    .io_ins_306(rport_io_ins_306),
    .io_ins_307(rport_io_ins_307),
    .io_ins_308(rport_io_ins_308),
    .io_ins_309(rport_io_ins_309),
    .io_ins_310(rport_io_ins_310),
    .io_ins_311(rport_io_ins_311),
    .io_ins_312(rport_io_ins_312),
    .io_ins_313(rport_io_ins_313),
    .io_ins_314(rport_io_ins_314),
    .io_ins_315(rport_io_ins_315),
    .io_ins_316(rport_io_ins_316),
    .io_ins_317(rport_io_ins_317),
    .io_ins_318(rport_io_ins_318),
    .io_ins_319(rport_io_ins_319),
    .io_ins_320(rport_io_ins_320),
    .io_ins_321(rport_io_ins_321),
    .io_ins_322(rport_io_ins_322),
    .io_ins_323(rport_io_ins_323),
    .io_ins_324(rport_io_ins_324),
    .io_ins_325(rport_io_ins_325),
    .io_ins_326(rport_io_ins_326),
    .io_ins_327(rport_io_ins_327),
    .io_ins_328(rport_io_ins_328),
    .io_ins_329(rport_io_ins_329),
    .io_ins_330(rport_io_ins_330),
    .io_ins_331(rport_io_ins_331),
    .io_ins_332(rport_io_ins_332),
    .io_ins_333(rport_io_ins_333),
    .io_ins_334(rport_io_ins_334),
    .io_ins_335(rport_io_ins_335),
    .io_ins_336(rport_io_ins_336),
    .io_ins_337(rport_io_ins_337),
    .io_ins_338(rport_io_ins_338),
    .io_ins_339(rport_io_ins_339),
    .io_ins_340(rport_io_ins_340),
    .io_ins_341(rport_io_ins_341),
    .io_ins_342(rport_io_ins_342),
    .io_ins_343(rport_io_ins_343),
    .io_ins_344(rport_io_ins_344),
    .io_ins_345(rport_io_ins_345),
    .io_ins_346(rport_io_ins_346),
    .io_ins_347(rport_io_ins_347),
    .io_ins_348(rport_io_ins_348),
    .io_ins_349(rport_io_ins_349),
    .io_ins_350(rport_io_ins_350),
    .io_ins_351(rport_io_ins_351),
    .io_ins_352(rport_io_ins_352),
    .io_ins_353(rport_io_ins_353),
    .io_ins_354(rport_io_ins_354),
    .io_ins_355(rport_io_ins_355),
    .io_ins_356(rport_io_ins_356),
    .io_ins_357(rport_io_ins_357),
    .io_ins_358(rport_io_ins_358),
    .io_ins_359(rport_io_ins_359),
    .io_ins_360(rport_io_ins_360),
    .io_ins_361(rport_io_ins_361),
    .io_ins_362(rport_io_ins_362),
    .io_ins_363(rport_io_ins_363),
    .io_ins_364(rport_io_ins_364),
    .io_ins_365(rport_io_ins_365),
    .io_ins_366(rport_io_ins_366),
    .io_ins_367(rport_io_ins_367),
    .io_ins_368(rport_io_ins_368),
    .io_ins_369(rport_io_ins_369),
    .io_ins_370(rport_io_ins_370),
    .io_ins_371(rport_io_ins_371),
    .io_ins_372(rport_io_ins_372),
    .io_ins_373(rport_io_ins_373),
    .io_ins_374(rport_io_ins_374),
    .io_ins_375(rport_io_ins_375),
    .io_ins_376(rport_io_ins_376),
    .io_ins_377(rport_io_ins_377),
    .io_ins_378(rport_io_ins_378),
    .io_ins_379(rport_io_ins_379),
    .io_ins_380(rport_io_ins_380),
    .io_ins_381(rport_io_ins_381),
    .io_ins_382(rport_io_ins_382),
    .io_ins_383(rport_io_ins_383),
    .io_ins_384(rport_io_ins_384),
    .io_ins_385(rport_io_ins_385),
    .io_ins_386(rport_io_ins_386),
    .io_ins_387(rport_io_ins_387),
    .io_ins_388(rport_io_ins_388),
    .io_ins_389(rport_io_ins_389),
    .io_ins_390(rport_io_ins_390),
    .io_ins_391(rport_io_ins_391),
    .io_ins_392(rport_io_ins_392),
    .io_ins_393(rport_io_ins_393),
    .io_ins_394(rport_io_ins_394),
    .io_ins_395(rport_io_ins_395),
    .io_ins_396(rport_io_ins_396),
    .io_ins_397(rport_io_ins_397),
    .io_ins_398(rport_io_ins_398),
    .io_ins_399(rport_io_ins_399),
    .io_ins_400(rport_io_ins_400),
    .io_ins_401(rport_io_ins_401),
    .io_ins_402(rport_io_ins_402),
    .io_ins_403(rport_io_ins_403),
    .io_ins_404(rport_io_ins_404),
    .io_ins_405(rport_io_ins_405),
    .io_ins_406(rport_io_ins_406),
    .io_ins_407(rport_io_ins_407),
    .io_ins_408(rport_io_ins_408),
    .io_ins_409(rport_io_ins_409),
    .io_ins_410(rport_io_ins_410),
    .io_ins_411(rport_io_ins_411),
    .io_ins_412(rport_io_ins_412),
    .io_ins_413(rport_io_ins_413),
    .io_ins_414(rport_io_ins_414),
    .io_ins_415(rport_io_ins_415),
    .io_ins_416(rport_io_ins_416),
    .io_ins_417(rport_io_ins_417),
    .io_ins_418(rport_io_ins_418),
    .io_ins_419(rport_io_ins_419),
    .io_ins_420(rport_io_ins_420),
    .io_ins_421(rport_io_ins_421),
    .io_ins_422(rport_io_ins_422),
    .io_ins_423(rport_io_ins_423),
    .io_ins_424(rport_io_ins_424),
    .io_ins_425(rport_io_ins_425),
    .io_ins_426(rport_io_ins_426),
    .io_ins_427(rport_io_ins_427),
    .io_ins_428(rport_io_ins_428),
    .io_ins_429(rport_io_ins_429),
    .io_ins_430(rport_io_ins_430),
    .io_ins_431(rport_io_ins_431),
    .io_ins_432(rport_io_ins_432),
    .io_ins_433(rport_io_ins_433),
    .io_ins_434(rport_io_ins_434),
    .io_ins_435(rport_io_ins_435),
    .io_ins_436(rport_io_ins_436),
    .io_ins_437(rport_io_ins_437),
    .io_ins_438(rport_io_ins_438),
    .io_ins_439(rport_io_ins_439),
    .io_ins_440(rport_io_ins_440),
    .io_ins_441(rport_io_ins_441),
    .io_ins_442(rport_io_ins_442),
    .io_ins_443(rport_io_ins_443),
    .io_ins_444(rport_io_ins_444),
    .io_ins_445(rport_io_ins_445),
    .io_ins_446(rport_io_ins_446),
    .io_ins_447(rport_io_ins_447),
    .io_ins_448(rport_io_ins_448),
    .io_ins_449(rport_io_ins_449),
    .io_ins_450(rport_io_ins_450),
    .io_ins_451(rport_io_ins_451),
    .io_ins_452(rport_io_ins_452),
    .io_ins_453(rport_io_ins_453),
    .io_ins_454(rport_io_ins_454),
    .io_ins_455(rport_io_ins_455),
    .io_ins_456(rport_io_ins_456),
    .io_ins_457(rport_io_ins_457),
    .io_ins_458(rport_io_ins_458),
    .io_ins_459(rport_io_ins_459),
    .io_ins_460(rport_io_ins_460),
    .io_ins_461(rport_io_ins_461),
    .io_ins_462(rport_io_ins_462),
    .io_ins_463(rport_io_ins_463),
    .io_ins_464(rport_io_ins_464),
    .io_ins_465(rport_io_ins_465),
    .io_ins_466(rport_io_ins_466),
    .io_ins_467(rport_io_ins_467),
    .io_ins_468(rport_io_ins_468),
    .io_ins_469(rport_io_ins_469),
    .io_ins_470(rport_io_ins_470),
    .io_ins_471(rport_io_ins_471),
    .io_ins_472(rport_io_ins_472),
    .io_ins_473(rport_io_ins_473),
    .io_ins_474(rport_io_ins_474),
    .io_ins_475(rport_io_ins_475),
    .io_ins_476(rport_io_ins_476),
    .io_ins_477(rport_io_ins_477),
    .io_ins_478(rport_io_ins_478),
    .io_ins_479(rport_io_ins_479),
    .io_ins_480(rport_io_ins_480),
    .io_ins_481(rport_io_ins_481),
    .io_ins_482(rport_io_ins_482),
    .io_ins_483(rport_io_ins_483),
    .io_ins_484(rport_io_ins_484),
    .io_ins_485(rport_io_ins_485),
    .io_ins_486(rport_io_ins_486),
    .io_ins_487(rport_io_ins_487),
    .io_ins_488(rport_io_ins_488),
    .io_ins_489(rport_io_ins_489),
    .io_ins_490(rport_io_ins_490),
    .io_ins_491(rport_io_ins_491),
    .io_ins_492(rport_io_ins_492),
    .io_ins_493(rport_io_ins_493),
    .io_ins_494(rport_io_ins_494),
    .io_ins_495(rport_io_ins_495),
    .io_ins_496(rport_io_ins_496),
    .io_ins_497(rport_io_ins_497),
    .io_ins_498(rport_io_ins_498),
    .io_ins_499(rport_io_ins_499),
    .io_ins_500(rport_io_ins_500),
    .io_ins_501(rport_io_ins_501),
    .io_ins_502(rport_io_ins_502),
    .io_ins_503(rport_io_ins_503),
    .io_ins_504(rport_io_ins_504),
    .io_ins_505(rport_io_ins_505),
    .io_ins_506(rport_io_ins_506),
    .io_ins_507(rport_io_ins_507),
    .io_ins_508(rport_io_ins_508),
    .io_ins_509(rport_io_ins_509),
    .io_ins_510(rport_io_ins_510),
    .io_ins_511(rport_io_ins_511),
    .io_sel(rport_io_sel),
    .io_out(rport_io_out)
  );
  assign _T_3130 = io_waddr == 32'h0; // @[RegFile.scala 80:42:@37631.4]
  assign _T_3136 = io_waddr == 32'h1; // @[RegFile.scala 68:46:@37643.4]
  assign _T_3137 = io_wen & _T_3136; // @[RegFile.scala 68:34:@37644.4]
  assign _T_3150 = io_waddr == 32'h2; // @[RegFile.scala 80:42:@37662.4]
  assign _T_3156 = io_waddr == 32'h3; // @[RegFile.scala 74:80:@37674.4]
  assign _T_3157 = io_wen & _T_3156; // @[RegFile.scala 74:68:@37675.4]
  assign _T_3163 = io_waddr == 32'h4; // @[RegFile.scala 74:80:@37688.4]
  assign _T_3164 = io_wen & _T_3163; // @[RegFile.scala 74:68:@37689.4]
  assign _T_3170 = io_waddr == 32'h5; // @[RegFile.scala 74:80:@37702.4]
  assign _T_3171 = io_wen & _T_3170; // @[RegFile.scala 74:68:@37703.4]
  assign _T_3177 = io_waddr == 32'h6; // @[RegFile.scala 74:80:@37716.4]
  assign _T_3178 = io_wen & _T_3177; // @[RegFile.scala 74:68:@37717.4]
  assign _T_3184 = io_waddr == 32'h7; // @[RegFile.scala 74:80:@37730.4]
  assign _T_3185 = io_wen & _T_3184; // @[RegFile.scala 74:68:@37731.4]
  assign _T_3191 = io_waddr == 32'h8; // @[RegFile.scala 74:80:@37744.4]
  assign _T_3192 = io_wen & _T_3191; // @[RegFile.scala 74:68:@37745.4]
  assign _T_3198 = io_waddr == 32'h9; // @[RegFile.scala 74:80:@37758.4]
  assign _T_3199 = io_wen & _T_3198; // @[RegFile.scala 74:68:@37759.4]
  assign _T_3205 = io_waddr == 32'ha; // @[RegFile.scala 74:80:@37772.4]
  assign _T_3206 = io_wen & _T_3205; // @[RegFile.scala 74:68:@37773.4]
  assign _T_3212 = io_waddr == 32'hb; // @[RegFile.scala 74:80:@37786.4]
  assign _T_3213 = io_wen & _T_3212; // @[RegFile.scala 74:68:@37787.4]
  assign _T_3219 = io_waddr == 32'hc; // @[RegFile.scala 74:80:@37800.4]
  assign _T_3220 = io_wen & _T_3219; // @[RegFile.scala 74:68:@37801.4]
  assign io_rdata = rport_io_out; // @[RegFile.scala 107:14:@45826.4]
  assign io_argIns_0 = regs_0_io_out; // @[RegFile.scala 111:13:@45831.4]
  assign io_argIns_1 = regs_1_io_out; // @[RegFile.scala 111:13:@45832.4]
  assign io_argIns_2 = regs_2_io_out; // @[RegFile.scala 111:13:@45833.4]
  assign regs_0_clock = clock; // @[:@37629.4]
  assign regs_0_reset = reset; // @[:@37630.4 RegFile.scala 82:16:@37636.4]
  assign regs_0_io_in = io_wdata; // @[RegFile.scala 81:16:@37634.4]
  assign regs_0_io_reset = reset; // @[RegFile.scala 83:19:@37638.4]
  assign regs_0_io_enable = io_wen & _T_3130; // @[RegFile.scala 80:20:@37633.4]
  assign regs_1_clock = clock; // @[:@37641.4]
  assign regs_1_reset = reset; // @[:@37642.4 RegFile.scala 70:16:@37654.4]
  assign regs_1_io_in = _T_3137 ? io_wdata : io_argOuts_0_bits; // @[RegFile.scala 69:16:@37652.4]
  assign regs_1_io_reset = reset; // @[RegFile.scala 72:19:@37657.4]
  assign regs_1_io_enable = _T_3137 ? _T_3137 : io_argOuts_0_valid; // @[RegFile.scala 68:20:@37648.4]
  assign regs_2_clock = clock; // @[:@37660.4]
  assign regs_2_reset = reset; // @[:@37661.4 RegFile.scala 82:16:@37667.4]
  assign regs_2_io_in = io_wdata; // @[RegFile.scala 81:16:@37665.4]
  assign regs_2_io_reset = reset; // @[RegFile.scala 83:19:@37669.4]
  assign regs_2_io_enable = io_wen & _T_3150; // @[RegFile.scala 80:20:@37664.4]
  assign regs_3_clock = clock; // @[:@37672.4]
  assign regs_3_reset = io_reset; // @[:@37673.4 RegFile.scala 76:16:@37680.4]
  assign regs_3_io_in = io_argOuts_1_valid ? io_argOuts_1_bits : io_wdata; // @[RegFile.scala 75:16:@37679.4]
  assign regs_3_io_reset = reset; // @[RegFile.scala 78:19:@37683.4]
  assign regs_3_io_enable = io_argOuts_1_valid | _T_3157; // @[RegFile.scala 74:20:@37677.4]
  assign regs_4_clock = clock; // @[:@37686.4]
  assign regs_4_reset = io_reset; // @[:@37687.4 RegFile.scala 76:16:@37694.4]
  assign regs_4_io_in = io_argOuts_2_valid ? io_argOuts_2_bits : io_wdata; // @[RegFile.scala 75:16:@37693.4]
  assign regs_4_io_reset = reset; // @[RegFile.scala 78:19:@37697.4]
  assign regs_4_io_enable = io_argOuts_2_valid | _T_3164; // @[RegFile.scala 74:20:@37691.4]
  assign regs_5_clock = clock; // @[:@37700.4]
  assign regs_5_reset = io_reset; // @[:@37701.4 RegFile.scala 76:16:@37708.4]
  assign regs_5_io_in = io_argOuts_3_valid ? io_argOuts_3_bits : io_wdata; // @[RegFile.scala 75:16:@37707.4]
  assign regs_5_io_reset = reset; // @[RegFile.scala 78:19:@37711.4]
  assign regs_5_io_enable = io_argOuts_3_valid | _T_3171; // @[RegFile.scala 74:20:@37705.4]
  assign regs_6_clock = clock; // @[:@37714.4]
  assign regs_6_reset = io_reset; // @[:@37715.4 RegFile.scala 76:16:@37722.4]
  assign regs_6_io_in = io_argOuts_4_valid ? io_argOuts_4_bits : io_wdata; // @[RegFile.scala 75:16:@37721.4]
  assign regs_6_io_reset = reset; // @[RegFile.scala 78:19:@37725.4]
  assign regs_6_io_enable = io_argOuts_4_valid | _T_3178; // @[RegFile.scala 74:20:@37719.4]
  assign regs_7_clock = clock; // @[:@37728.4]
  assign regs_7_reset = io_reset; // @[:@37729.4 RegFile.scala 76:16:@37736.4]
  assign regs_7_io_in = io_argOuts_5_valid ? io_argOuts_5_bits : io_wdata; // @[RegFile.scala 75:16:@37735.4]
  assign regs_7_io_reset = reset; // @[RegFile.scala 78:19:@37739.4]
  assign regs_7_io_enable = io_argOuts_5_valid | _T_3185; // @[RegFile.scala 74:20:@37733.4]
  assign regs_8_clock = clock; // @[:@37742.4]
  assign regs_8_reset = io_reset; // @[:@37743.4 RegFile.scala 76:16:@37750.4]
  assign regs_8_io_in = io_argOuts_6_valid ? io_argOuts_6_bits : io_wdata; // @[RegFile.scala 75:16:@37749.4]
  assign regs_8_io_reset = reset; // @[RegFile.scala 78:19:@37753.4]
  assign regs_8_io_enable = io_argOuts_6_valid | _T_3192; // @[RegFile.scala 74:20:@37747.4]
  assign regs_9_clock = clock; // @[:@37756.4]
  assign regs_9_reset = io_reset; // @[:@37757.4 RegFile.scala 76:16:@37764.4]
  assign regs_9_io_in = io_argOuts_7_valid ? io_argOuts_7_bits : io_wdata; // @[RegFile.scala 75:16:@37763.4]
  assign regs_9_io_reset = reset; // @[RegFile.scala 78:19:@37767.4]
  assign regs_9_io_enable = io_argOuts_7_valid | _T_3199; // @[RegFile.scala 74:20:@37761.4]
  assign regs_10_clock = clock; // @[:@37770.4]
  assign regs_10_reset = io_reset; // @[:@37771.4 RegFile.scala 76:16:@37778.4]
  assign regs_10_io_in = io_argOuts_8_valid ? io_argOuts_8_bits : io_wdata; // @[RegFile.scala 75:16:@37777.4]
  assign regs_10_io_reset = reset; // @[RegFile.scala 78:19:@37781.4]
  assign regs_10_io_enable = io_argOuts_8_valid | _T_3206; // @[RegFile.scala 74:20:@37775.4]
  assign regs_11_clock = clock; // @[:@37784.4]
  assign regs_11_reset = io_reset; // @[:@37785.4 RegFile.scala 76:16:@37792.4]
  assign regs_11_io_in = io_argOuts_9_valid ? io_argOuts_9_bits : io_wdata; // @[RegFile.scala 75:16:@37791.4]
  assign regs_11_io_reset = reset; // @[RegFile.scala 78:19:@37795.4]
  assign regs_11_io_enable = io_argOuts_9_valid | _T_3213; // @[RegFile.scala 74:20:@37789.4]
  assign regs_12_clock = clock; // @[:@37798.4]
  assign regs_12_reset = io_reset; // @[:@37799.4 RegFile.scala 76:16:@37806.4]
  assign regs_12_io_in = io_argOuts_10_valid ? io_argOuts_10_bits : io_wdata; // @[RegFile.scala 75:16:@37805.4]
  assign regs_12_io_reset = reset; // @[RegFile.scala 78:19:@37809.4]
  assign regs_12_io_enable = io_argOuts_10_valid | _T_3220; // @[RegFile.scala 74:20:@37803.4]
  assign regs_13_clock = clock; // @[:@37812.4]
  assign regs_13_reset = io_reset; // @[:@37813.4 RegFile.scala 76:16:@37820.4]
  assign regs_13_io_in = 64'h0; // @[RegFile.scala 75:16:@37819.4]
  assign regs_13_io_reset = reset; // @[RegFile.scala 78:19:@37823.4]
  assign regs_13_io_enable = 1'h1; // @[RegFile.scala 74:20:@37817.4]
  assign regs_14_clock = clock; // @[:@37826.4]
  assign regs_14_reset = io_reset; // @[:@37827.4 RegFile.scala 76:16:@37834.4]
  assign regs_14_io_in = 64'h0; // @[RegFile.scala 75:16:@37833.4]
  assign regs_14_io_reset = reset; // @[RegFile.scala 78:19:@37837.4]
  assign regs_14_io_enable = 1'h1; // @[RegFile.scala 74:20:@37831.4]
  assign regs_15_clock = clock; // @[:@37840.4]
  assign regs_15_reset = io_reset; // @[:@37841.4 RegFile.scala 76:16:@37848.4]
  assign regs_15_io_in = 64'h0; // @[RegFile.scala 75:16:@37847.4]
  assign regs_15_io_reset = reset; // @[RegFile.scala 78:19:@37851.4]
  assign regs_15_io_enable = 1'h1; // @[RegFile.scala 74:20:@37845.4]
  assign regs_16_clock = clock; // @[:@37854.4]
  assign regs_16_reset = io_reset; // @[:@37855.4 RegFile.scala 76:16:@37862.4]
  assign regs_16_io_in = 64'h0; // @[RegFile.scala 75:16:@37861.4]
  assign regs_16_io_reset = reset; // @[RegFile.scala 78:19:@37865.4]
  assign regs_16_io_enable = 1'h1; // @[RegFile.scala 74:20:@37859.4]
  assign regs_17_clock = clock; // @[:@37868.4]
  assign regs_17_reset = io_reset; // @[:@37869.4 RegFile.scala 76:16:@37876.4]
  assign regs_17_io_in = 64'h0; // @[RegFile.scala 75:16:@37875.4]
  assign regs_17_io_reset = reset; // @[RegFile.scala 78:19:@37879.4]
  assign regs_17_io_enable = 1'h1; // @[RegFile.scala 74:20:@37873.4]
  assign regs_18_clock = clock; // @[:@37882.4]
  assign regs_18_reset = io_reset; // @[:@37883.4 RegFile.scala 76:16:@37890.4]
  assign regs_18_io_in = 64'h0; // @[RegFile.scala 75:16:@37889.4]
  assign regs_18_io_reset = reset; // @[RegFile.scala 78:19:@37893.4]
  assign regs_18_io_enable = 1'h1; // @[RegFile.scala 74:20:@37887.4]
  assign regs_19_clock = clock; // @[:@37896.4]
  assign regs_19_reset = io_reset; // @[:@37897.4 RegFile.scala 76:16:@37904.4]
  assign regs_19_io_in = 64'h0; // @[RegFile.scala 75:16:@37903.4]
  assign regs_19_io_reset = reset; // @[RegFile.scala 78:19:@37907.4]
  assign regs_19_io_enable = 1'h1; // @[RegFile.scala 74:20:@37901.4]
  assign regs_20_clock = clock; // @[:@37910.4]
  assign regs_20_reset = io_reset; // @[:@37911.4 RegFile.scala 76:16:@37918.4]
  assign regs_20_io_in = 64'h0; // @[RegFile.scala 75:16:@37917.4]
  assign regs_20_io_reset = reset; // @[RegFile.scala 78:19:@37921.4]
  assign regs_20_io_enable = 1'h1; // @[RegFile.scala 74:20:@37915.4]
  assign regs_21_clock = clock; // @[:@37924.4]
  assign regs_21_reset = io_reset; // @[:@37925.4 RegFile.scala 76:16:@37932.4]
  assign regs_21_io_in = 64'h0; // @[RegFile.scala 75:16:@37931.4]
  assign regs_21_io_reset = reset; // @[RegFile.scala 78:19:@37935.4]
  assign regs_21_io_enable = 1'h1; // @[RegFile.scala 74:20:@37929.4]
  assign regs_22_clock = clock; // @[:@37938.4]
  assign regs_22_reset = io_reset; // @[:@37939.4 RegFile.scala 76:16:@37946.4]
  assign regs_22_io_in = 64'h0; // @[RegFile.scala 75:16:@37945.4]
  assign regs_22_io_reset = reset; // @[RegFile.scala 78:19:@37949.4]
  assign regs_22_io_enable = 1'h1; // @[RegFile.scala 74:20:@37943.4]
  assign regs_23_clock = clock; // @[:@37952.4]
  assign regs_23_reset = io_reset; // @[:@37953.4 RegFile.scala 76:16:@37960.4]
  assign regs_23_io_in = 64'h0; // @[RegFile.scala 75:16:@37959.4]
  assign regs_23_io_reset = reset; // @[RegFile.scala 78:19:@37963.4]
  assign regs_23_io_enable = 1'h1; // @[RegFile.scala 74:20:@37957.4]
  assign regs_24_clock = clock; // @[:@37966.4]
  assign regs_24_reset = io_reset; // @[:@37967.4 RegFile.scala 76:16:@37974.4]
  assign regs_24_io_in = 64'h0; // @[RegFile.scala 75:16:@37973.4]
  assign regs_24_io_reset = reset; // @[RegFile.scala 78:19:@37977.4]
  assign regs_24_io_enable = 1'h1; // @[RegFile.scala 74:20:@37971.4]
  assign regs_25_clock = clock; // @[:@37980.4]
  assign regs_25_reset = io_reset; // @[:@37981.4 RegFile.scala 76:16:@37988.4]
  assign regs_25_io_in = 64'h0; // @[RegFile.scala 75:16:@37987.4]
  assign regs_25_io_reset = reset; // @[RegFile.scala 78:19:@37991.4]
  assign regs_25_io_enable = 1'h1; // @[RegFile.scala 74:20:@37985.4]
  assign regs_26_clock = clock; // @[:@37994.4]
  assign regs_26_reset = io_reset; // @[:@37995.4 RegFile.scala 76:16:@38002.4]
  assign regs_26_io_in = 64'h0; // @[RegFile.scala 75:16:@38001.4]
  assign regs_26_io_reset = reset; // @[RegFile.scala 78:19:@38005.4]
  assign regs_26_io_enable = 1'h1; // @[RegFile.scala 74:20:@37999.4]
  assign regs_27_clock = clock; // @[:@38008.4]
  assign regs_27_reset = io_reset; // @[:@38009.4 RegFile.scala 76:16:@38016.4]
  assign regs_27_io_in = 64'h0; // @[RegFile.scala 75:16:@38015.4]
  assign regs_27_io_reset = reset; // @[RegFile.scala 78:19:@38019.4]
  assign regs_27_io_enable = 1'h1; // @[RegFile.scala 74:20:@38013.4]
  assign regs_28_clock = clock; // @[:@38022.4]
  assign regs_28_reset = io_reset; // @[:@38023.4 RegFile.scala 76:16:@38030.4]
  assign regs_28_io_in = 64'h0; // @[RegFile.scala 75:16:@38029.4]
  assign regs_28_io_reset = reset; // @[RegFile.scala 78:19:@38033.4]
  assign regs_28_io_enable = 1'h1; // @[RegFile.scala 74:20:@38027.4]
  assign regs_29_clock = clock; // @[:@38036.4]
  assign regs_29_reset = io_reset; // @[:@38037.4 RegFile.scala 76:16:@38044.4]
  assign regs_29_io_in = 64'h0; // @[RegFile.scala 75:16:@38043.4]
  assign regs_29_io_reset = reset; // @[RegFile.scala 78:19:@38047.4]
  assign regs_29_io_enable = 1'h1; // @[RegFile.scala 74:20:@38041.4]
  assign regs_30_clock = clock; // @[:@38050.4]
  assign regs_30_reset = io_reset; // @[:@38051.4 RegFile.scala 76:16:@38058.4]
  assign regs_30_io_in = 64'h0; // @[RegFile.scala 75:16:@38057.4]
  assign regs_30_io_reset = reset; // @[RegFile.scala 78:19:@38061.4]
  assign regs_30_io_enable = 1'h1; // @[RegFile.scala 74:20:@38055.4]
  assign regs_31_clock = clock; // @[:@38064.4]
  assign regs_31_reset = io_reset; // @[:@38065.4 RegFile.scala 76:16:@38072.4]
  assign regs_31_io_in = 64'h0; // @[RegFile.scala 75:16:@38071.4]
  assign regs_31_io_reset = reset; // @[RegFile.scala 78:19:@38075.4]
  assign regs_31_io_enable = 1'h1; // @[RegFile.scala 74:20:@38069.4]
  assign regs_32_clock = clock; // @[:@38078.4]
  assign regs_32_reset = io_reset; // @[:@38079.4 RegFile.scala 76:16:@38086.4]
  assign regs_32_io_in = 64'h0; // @[RegFile.scala 75:16:@38085.4]
  assign regs_32_io_reset = reset; // @[RegFile.scala 78:19:@38089.4]
  assign regs_32_io_enable = 1'h1; // @[RegFile.scala 74:20:@38083.4]
  assign regs_33_clock = clock; // @[:@38092.4]
  assign regs_33_reset = io_reset; // @[:@38093.4 RegFile.scala 76:16:@38100.4]
  assign regs_33_io_in = 64'h0; // @[RegFile.scala 75:16:@38099.4]
  assign regs_33_io_reset = reset; // @[RegFile.scala 78:19:@38103.4]
  assign regs_33_io_enable = 1'h1; // @[RegFile.scala 74:20:@38097.4]
  assign regs_34_clock = clock; // @[:@38106.4]
  assign regs_34_reset = io_reset; // @[:@38107.4 RegFile.scala 76:16:@38114.4]
  assign regs_34_io_in = 64'h0; // @[RegFile.scala 75:16:@38113.4]
  assign regs_34_io_reset = reset; // @[RegFile.scala 78:19:@38117.4]
  assign regs_34_io_enable = 1'h1; // @[RegFile.scala 74:20:@38111.4]
  assign regs_35_clock = clock; // @[:@38120.4]
  assign regs_35_reset = io_reset; // @[:@38121.4 RegFile.scala 76:16:@38128.4]
  assign regs_35_io_in = 64'h0; // @[RegFile.scala 75:16:@38127.4]
  assign regs_35_io_reset = reset; // @[RegFile.scala 78:19:@38131.4]
  assign regs_35_io_enable = 1'h1; // @[RegFile.scala 74:20:@38125.4]
  assign regs_36_clock = clock; // @[:@38134.4]
  assign regs_36_reset = io_reset; // @[:@38135.4 RegFile.scala 76:16:@38142.4]
  assign regs_36_io_in = 64'h0; // @[RegFile.scala 75:16:@38141.4]
  assign regs_36_io_reset = reset; // @[RegFile.scala 78:19:@38145.4]
  assign regs_36_io_enable = 1'h1; // @[RegFile.scala 74:20:@38139.4]
  assign regs_37_clock = clock; // @[:@38148.4]
  assign regs_37_reset = io_reset; // @[:@38149.4 RegFile.scala 76:16:@38156.4]
  assign regs_37_io_in = 64'h0; // @[RegFile.scala 75:16:@38155.4]
  assign regs_37_io_reset = reset; // @[RegFile.scala 78:19:@38159.4]
  assign regs_37_io_enable = 1'h1; // @[RegFile.scala 74:20:@38153.4]
  assign regs_38_clock = clock; // @[:@38162.4]
  assign regs_38_reset = io_reset; // @[:@38163.4 RegFile.scala 76:16:@38170.4]
  assign regs_38_io_in = 64'h0; // @[RegFile.scala 75:16:@38169.4]
  assign regs_38_io_reset = reset; // @[RegFile.scala 78:19:@38173.4]
  assign regs_38_io_enable = 1'h1; // @[RegFile.scala 74:20:@38167.4]
  assign regs_39_clock = clock; // @[:@38176.4]
  assign regs_39_reset = io_reset; // @[:@38177.4 RegFile.scala 76:16:@38184.4]
  assign regs_39_io_in = 64'h0; // @[RegFile.scala 75:16:@38183.4]
  assign regs_39_io_reset = reset; // @[RegFile.scala 78:19:@38187.4]
  assign regs_39_io_enable = 1'h1; // @[RegFile.scala 74:20:@38181.4]
  assign regs_40_clock = clock; // @[:@38190.4]
  assign regs_40_reset = io_reset; // @[:@38191.4 RegFile.scala 76:16:@38198.4]
  assign regs_40_io_in = 64'h0; // @[RegFile.scala 75:16:@38197.4]
  assign regs_40_io_reset = reset; // @[RegFile.scala 78:19:@38201.4]
  assign regs_40_io_enable = 1'h1; // @[RegFile.scala 74:20:@38195.4]
  assign regs_41_clock = clock; // @[:@38204.4]
  assign regs_41_reset = io_reset; // @[:@38205.4 RegFile.scala 76:16:@38212.4]
  assign regs_41_io_in = 64'h0; // @[RegFile.scala 75:16:@38211.4]
  assign regs_41_io_reset = reset; // @[RegFile.scala 78:19:@38215.4]
  assign regs_41_io_enable = 1'h1; // @[RegFile.scala 74:20:@38209.4]
  assign regs_42_clock = clock; // @[:@38218.4]
  assign regs_42_reset = io_reset; // @[:@38219.4 RegFile.scala 76:16:@38226.4]
  assign regs_42_io_in = 64'h0; // @[RegFile.scala 75:16:@38225.4]
  assign regs_42_io_reset = reset; // @[RegFile.scala 78:19:@38229.4]
  assign regs_42_io_enable = 1'h1; // @[RegFile.scala 74:20:@38223.4]
  assign regs_43_clock = clock; // @[:@38232.4]
  assign regs_43_reset = io_reset; // @[:@38233.4 RegFile.scala 76:16:@38240.4]
  assign regs_43_io_in = 64'h0; // @[RegFile.scala 75:16:@38239.4]
  assign regs_43_io_reset = reset; // @[RegFile.scala 78:19:@38243.4]
  assign regs_43_io_enable = 1'h1; // @[RegFile.scala 74:20:@38237.4]
  assign regs_44_clock = clock; // @[:@38246.4]
  assign regs_44_reset = io_reset; // @[:@38247.4 RegFile.scala 76:16:@38254.4]
  assign regs_44_io_in = 64'h0; // @[RegFile.scala 75:16:@38253.4]
  assign regs_44_io_reset = reset; // @[RegFile.scala 78:19:@38257.4]
  assign regs_44_io_enable = 1'h1; // @[RegFile.scala 74:20:@38251.4]
  assign regs_45_clock = clock; // @[:@38260.4]
  assign regs_45_reset = io_reset; // @[:@38261.4 RegFile.scala 76:16:@38268.4]
  assign regs_45_io_in = 64'h0; // @[RegFile.scala 75:16:@38267.4]
  assign regs_45_io_reset = reset; // @[RegFile.scala 78:19:@38271.4]
  assign regs_45_io_enable = 1'h1; // @[RegFile.scala 74:20:@38265.4]
  assign regs_46_clock = clock; // @[:@38274.4]
  assign regs_46_reset = io_reset; // @[:@38275.4 RegFile.scala 76:16:@38282.4]
  assign regs_46_io_in = 64'h0; // @[RegFile.scala 75:16:@38281.4]
  assign regs_46_io_reset = reset; // @[RegFile.scala 78:19:@38285.4]
  assign regs_46_io_enable = 1'h1; // @[RegFile.scala 74:20:@38279.4]
  assign regs_47_clock = clock; // @[:@38288.4]
  assign regs_47_reset = io_reset; // @[:@38289.4 RegFile.scala 76:16:@38296.4]
  assign regs_47_io_in = 64'h0; // @[RegFile.scala 75:16:@38295.4]
  assign regs_47_io_reset = reset; // @[RegFile.scala 78:19:@38299.4]
  assign regs_47_io_enable = 1'h1; // @[RegFile.scala 74:20:@38293.4]
  assign regs_48_clock = clock; // @[:@38302.4]
  assign regs_48_reset = io_reset; // @[:@38303.4 RegFile.scala 76:16:@38310.4]
  assign regs_48_io_in = 64'h0; // @[RegFile.scala 75:16:@38309.4]
  assign regs_48_io_reset = reset; // @[RegFile.scala 78:19:@38313.4]
  assign regs_48_io_enable = 1'h1; // @[RegFile.scala 74:20:@38307.4]
  assign regs_49_clock = clock; // @[:@38316.4]
  assign regs_49_reset = io_reset; // @[:@38317.4 RegFile.scala 76:16:@38324.4]
  assign regs_49_io_in = 64'h0; // @[RegFile.scala 75:16:@38323.4]
  assign regs_49_io_reset = reset; // @[RegFile.scala 78:19:@38327.4]
  assign regs_49_io_enable = 1'h1; // @[RegFile.scala 74:20:@38321.4]
  assign regs_50_clock = clock; // @[:@38330.4]
  assign regs_50_reset = io_reset; // @[:@38331.4 RegFile.scala 76:16:@38338.4]
  assign regs_50_io_in = 64'h0; // @[RegFile.scala 75:16:@38337.4]
  assign regs_50_io_reset = reset; // @[RegFile.scala 78:19:@38341.4]
  assign regs_50_io_enable = 1'h1; // @[RegFile.scala 74:20:@38335.4]
  assign regs_51_clock = clock; // @[:@38344.4]
  assign regs_51_reset = io_reset; // @[:@38345.4 RegFile.scala 76:16:@38352.4]
  assign regs_51_io_in = 64'h0; // @[RegFile.scala 75:16:@38351.4]
  assign regs_51_io_reset = reset; // @[RegFile.scala 78:19:@38355.4]
  assign regs_51_io_enable = 1'h1; // @[RegFile.scala 74:20:@38349.4]
  assign regs_52_clock = clock; // @[:@38358.4]
  assign regs_52_reset = io_reset; // @[:@38359.4 RegFile.scala 76:16:@38366.4]
  assign regs_52_io_in = 64'h0; // @[RegFile.scala 75:16:@38365.4]
  assign regs_52_io_reset = reset; // @[RegFile.scala 78:19:@38369.4]
  assign regs_52_io_enable = 1'h1; // @[RegFile.scala 74:20:@38363.4]
  assign regs_53_clock = clock; // @[:@38372.4]
  assign regs_53_reset = io_reset; // @[:@38373.4 RegFile.scala 76:16:@38380.4]
  assign regs_53_io_in = 64'h0; // @[RegFile.scala 75:16:@38379.4]
  assign regs_53_io_reset = reset; // @[RegFile.scala 78:19:@38383.4]
  assign regs_53_io_enable = 1'h1; // @[RegFile.scala 74:20:@38377.4]
  assign regs_54_clock = clock; // @[:@38386.4]
  assign regs_54_reset = io_reset; // @[:@38387.4 RegFile.scala 76:16:@38394.4]
  assign regs_54_io_in = 64'h0; // @[RegFile.scala 75:16:@38393.4]
  assign regs_54_io_reset = reset; // @[RegFile.scala 78:19:@38397.4]
  assign regs_54_io_enable = 1'h1; // @[RegFile.scala 74:20:@38391.4]
  assign regs_55_clock = clock; // @[:@38400.4]
  assign regs_55_reset = io_reset; // @[:@38401.4 RegFile.scala 76:16:@38408.4]
  assign regs_55_io_in = 64'h0; // @[RegFile.scala 75:16:@38407.4]
  assign regs_55_io_reset = reset; // @[RegFile.scala 78:19:@38411.4]
  assign regs_55_io_enable = 1'h1; // @[RegFile.scala 74:20:@38405.4]
  assign regs_56_clock = clock; // @[:@38414.4]
  assign regs_56_reset = io_reset; // @[:@38415.4 RegFile.scala 76:16:@38422.4]
  assign regs_56_io_in = 64'h0; // @[RegFile.scala 75:16:@38421.4]
  assign regs_56_io_reset = reset; // @[RegFile.scala 78:19:@38425.4]
  assign regs_56_io_enable = 1'h1; // @[RegFile.scala 74:20:@38419.4]
  assign regs_57_clock = clock; // @[:@38428.4]
  assign regs_57_reset = io_reset; // @[:@38429.4 RegFile.scala 76:16:@38436.4]
  assign regs_57_io_in = 64'h0; // @[RegFile.scala 75:16:@38435.4]
  assign regs_57_io_reset = reset; // @[RegFile.scala 78:19:@38439.4]
  assign regs_57_io_enable = 1'h1; // @[RegFile.scala 74:20:@38433.4]
  assign regs_58_clock = clock; // @[:@38442.4]
  assign regs_58_reset = io_reset; // @[:@38443.4 RegFile.scala 76:16:@38450.4]
  assign regs_58_io_in = 64'h0; // @[RegFile.scala 75:16:@38449.4]
  assign regs_58_io_reset = reset; // @[RegFile.scala 78:19:@38453.4]
  assign regs_58_io_enable = 1'h1; // @[RegFile.scala 74:20:@38447.4]
  assign regs_59_clock = clock; // @[:@38456.4]
  assign regs_59_reset = io_reset; // @[:@38457.4 RegFile.scala 76:16:@38464.4]
  assign regs_59_io_in = 64'h0; // @[RegFile.scala 75:16:@38463.4]
  assign regs_59_io_reset = reset; // @[RegFile.scala 78:19:@38467.4]
  assign regs_59_io_enable = 1'h1; // @[RegFile.scala 74:20:@38461.4]
  assign regs_60_clock = clock; // @[:@38470.4]
  assign regs_60_reset = io_reset; // @[:@38471.4 RegFile.scala 76:16:@38478.4]
  assign regs_60_io_in = 64'h0; // @[RegFile.scala 75:16:@38477.4]
  assign regs_60_io_reset = reset; // @[RegFile.scala 78:19:@38481.4]
  assign regs_60_io_enable = 1'h1; // @[RegFile.scala 74:20:@38475.4]
  assign regs_61_clock = clock; // @[:@38484.4]
  assign regs_61_reset = io_reset; // @[:@38485.4 RegFile.scala 76:16:@38492.4]
  assign regs_61_io_in = 64'h0; // @[RegFile.scala 75:16:@38491.4]
  assign regs_61_io_reset = reset; // @[RegFile.scala 78:19:@38495.4]
  assign regs_61_io_enable = 1'h1; // @[RegFile.scala 74:20:@38489.4]
  assign regs_62_clock = clock; // @[:@38498.4]
  assign regs_62_reset = io_reset; // @[:@38499.4 RegFile.scala 76:16:@38506.4]
  assign regs_62_io_in = 64'h0; // @[RegFile.scala 75:16:@38505.4]
  assign regs_62_io_reset = reset; // @[RegFile.scala 78:19:@38509.4]
  assign regs_62_io_enable = 1'h1; // @[RegFile.scala 74:20:@38503.4]
  assign regs_63_clock = clock; // @[:@38512.4]
  assign regs_63_reset = io_reset; // @[:@38513.4 RegFile.scala 76:16:@38520.4]
  assign regs_63_io_in = 64'h0; // @[RegFile.scala 75:16:@38519.4]
  assign regs_63_io_reset = reset; // @[RegFile.scala 78:19:@38523.4]
  assign regs_63_io_enable = 1'h1; // @[RegFile.scala 74:20:@38517.4]
  assign regs_64_clock = clock; // @[:@38526.4]
  assign regs_64_reset = io_reset; // @[:@38527.4 RegFile.scala 76:16:@38534.4]
  assign regs_64_io_in = 64'h0; // @[RegFile.scala 75:16:@38533.4]
  assign regs_64_io_reset = reset; // @[RegFile.scala 78:19:@38537.4]
  assign regs_64_io_enable = 1'h1; // @[RegFile.scala 74:20:@38531.4]
  assign regs_65_clock = clock; // @[:@38540.4]
  assign regs_65_reset = io_reset; // @[:@38541.4 RegFile.scala 76:16:@38548.4]
  assign regs_65_io_in = 64'h0; // @[RegFile.scala 75:16:@38547.4]
  assign regs_65_io_reset = reset; // @[RegFile.scala 78:19:@38551.4]
  assign regs_65_io_enable = 1'h1; // @[RegFile.scala 74:20:@38545.4]
  assign regs_66_clock = clock; // @[:@38554.4]
  assign regs_66_reset = io_reset; // @[:@38555.4 RegFile.scala 76:16:@38562.4]
  assign regs_66_io_in = 64'h0; // @[RegFile.scala 75:16:@38561.4]
  assign regs_66_io_reset = reset; // @[RegFile.scala 78:19:@38565.4]
  assign regs_66_io_enable = 1'h1; // @[RegFile.scala 74:20:@38559.4]
  assign regs_67_clock = clock; // @[:@38568.4]
  assign regs_67_reset = io_reset; // @[:@38569.4 RegFile.scala 76:16:@38576.4]
  assign regs_67_io_in = 64'h0; // @[RegFile.scala 75:16:@38575.4]
  assign regs_67_io_reset = reset; // @[RegFile.scala 78:19:@38579.4]
  assign regs_67_io_enable = 1'h1; // @[RegFile.scala 74:20:@38573.4]
  assign regs_68_clock = clock; // @[:@38582.4]
  assign regs_68_reset = io_reset; // @[:@38583.4 RegFile.scala 76:16:@38590.4]
  assign regs_68_io_in = 64'h0; // @[RegFile.scala 75:16:@38589.4]
  assign regs_68_io_reset = reset; // @[RegFile.scala 78:19:@38593.4]
  assign regs_68_io_enable = 1'h1; // @[RegFile.scala 74:20:@38587.4]
  assign regs_69_clock = clock; // @[:@38596.4]
  assign regs_69_reset = io_reset; // @[:@38597.4 RegFile.scala 76:16:@38604.4]
  assign regs_69_io_in = 64'h0; // @[RegFile.scala 75:16:@38603.4]
  assign regs_69_io_reset = reset; // @[RegFile.scala 78:19:@38607.4]
  assign regs_69_io_enable = 1'h1; // @[RegFile.scala 74:20:@38601.4]
  assign regs_70_clock = clock; // @[:@38610.4]
  assign regs_70_reset = io_reset; // @[:@38611.4 RegFile.scala 76:16:@38618.4]
  assign regs_70_io_in = 64'h0; // @[RegFile.scala 75:16:@38617.4]
  assign regs_70_io_reset = reset; // @[RegFile.scala 78:19:@38621.4]
  assign regs_70_io_enable = 1'h1; // @[RegFile.scala 74:20:@38615.4]
  assign regs_71_clock = clock; // @[:@38624.4]
  assign regs_71_reset = io_reset; // @[:@38625.4 RegFile.scala 76:16:@38632.4]
  assign regs_71_io_in = 64'h0; // @[RegFile.scala 75:16:@38631.4]
  assign regs_71_io_reset = reset; // @[RegFile.scala 78:19:@38635.4]
  assign regs_71_io_enable = 1'h1; // @[RegFile.scala 74:20:@38629.4]
  assign regs_72_clock = clock; // @[:@38638.4]
  assign regs_72_reset = io_reset; // @[:@38639.4 RegFile.scala 76:16:@38646.4]
  assign regs_72_io_in = 64'h0; // @[RegFile.scala 75:16:@38645.4]
  assign regs_72_io_reset = reset; // @[RegFile.scala 78:19:@38649.4]
  assign regs_72_io_enable = 1'h1; // @[RegFile.scala 74:20:@38643.4]
  assign regs_73_clock = clock; // @[:@38652.4]
  assign regs_73_reset = io_reset; // @[:@38653.4 RegFile.scala 76:16:@38660.4]
  assign regs_73_io_in = 64'h0; // @[RegFile.scala 75:16:@38659.4]
  assign regs_73_io_reset = reset; // @[RegFile.scala 78:19:@38663.4]
  assign regs_73_io_enable = 1'h1; // @[RegFile.scala 74:20:@38657.4]
  assign regs_74_clock = clock; // @[:@38666.4]
  assign regs_74_reset = io_reset; // @[:@38667.4 RegFile.scala 76:16:@38674.4]
  assign regs_74_io_in = 64'h0; // @[RegFile.scala 75:16:@38673.4]
  assign regs_74_io_reset = reset; // @[RegFile.scala 78:19:@38677.4]
  assign regs_74_io_enable = 1'h1; // @[RegFile.scala 74:20:@38671.4]
  assign regs_75_clock = clock; // @[:@38680.4]
  assign regs_75_reset = io_reset; // @[:@38681.4 RegFile.scala 76:16:@38688.4]
  assign regs_75_io_in = 64'h0; // @[RegFile.scala 75:16:@38687.4]
  assign regs_75_io_reset = reset; // @[RegFile.scala 78:19:@38691.4]
  assign regs_75_io_enable = 1'h1; // @[RegFile.scala 74:20:@38685.4]
  assign regs_76_clock = clock; // @[:@38694.4]
  assign regs_76_reset = io_reset; // @[:@38695.4 RegFile.scala 76:16:@38702.4]
  assign regs_76_io_in = 64'h0; // @[RegFile.scala 75:16:@38701.4]
  assign regs_76_io_reset = reset; // @[RegFile.scala 78:19:@38705.4]
  assign regs_76_io_enable = 1'h1; // @[RegFile.scala 74:20:@38699.4]
  assign regs_77_clock = clock; // @[:@38708.4]
  assign regs_77_reset = io_reset; // @[:@38709.4 RegFile.scala 76:16:@38716.4]
  assign regs_77_io_in = 64'h0; // @[RegFile.scala 75:16:@38715.4]
  assign regs_77_io_reset = reset; // @[RegFile.scala 78:19:@38719.4]
  assign regs_77_io_enable = 1'h1; // @[RegFile.scala 74:20:@38713.4]
  assign regs_78_clock = clock; // @[:@38722.4]
  assign regs_78_reset = io_reset; // @[:@38723.4 RegFile.scala 76:16:@38730.4]
  assign regs_78_io_in = 64'h0; // @[RegFile.scala 75:16:@38729.4]
  assign regs_78_io_reset = reset; // @[RegFile.scala 78:19:@38733.4]
  assign regs_78_io_enable = 1'h1; // @[RegFile.scala 74:20:@38727.4]
  assign regs_79_clock = clock; // @[:@38736.4]
  assign regs_79_reset = io_reset; // @[:@38737.4 RegFile.scala 76:16:@38744.4]
  assign regs_79_io_in = 64'h0; // @[RegFile.scala 75:16:@38743.4]
  assign regs_79_io_reset = reset; // @[RegFile.scala 78:19:@38747.4]
  assign regs_79_io_enable = 1'h1; // @[RegFile.scala 74:20:@38741.4]
  assign regs_80_clock = clock; // @[:@38750.4]
  assign regs_80_reset = io_reset; // @[:@38751.4 RegFile.scala 76:16:@38758.4]
  assign regs_80_io_in = 64'h0; // @[RegFile.scala 75:16:@38757.4]
  assign regs_80_io_reset = reset; // @[RegFile.scala 78:19:@38761.4]
  assign regs_80_io_enable = 1'h1; // @[RegFile.scala 74:20:@38755.4]
  assign regs_81_clock = clock; // @[:@38764.4]
  assign regs_81_reset = io_reset; // @[:@38765.4 RegFile.scala 76:16:@38772.4]
  assign regs_81_io_in = 64'h0; // @[RegFile.scala 75:16:@38771.4]
  assign regs_81_io_reset = reset; // @[RegFile.scala 78:19:@38775.4]
  assign regs_81_io_enable = 1'h1; // @[RegFile.scala 74:20:@38769.4]
  assign regs_82_clock = clock; // @[:@38778.4]
  assign regs_82_reset = io_reset; // @[:@38779.4 RegFile.scala 76:16:@38786.4]
  assign regs_82_io_in = 64'h0; // @[RegFile.scala 75:16:@38785.4]
  assign regs_82_io_reset = reset; // @[RegFile.scala 78:19:@38789.4]
  assign regs_82_io_enable = 1'h1; // @[RegFile.scala 74:20:@38783.4]
  assign regs_83_clock = clock; // @[:@38792.4]
  assign regs_83_reset = io_reset; // @[:@38793.4 RegFile.scala 76:16:@38800.4]
  assign regs_83_io_in = 64'h0; // @[RegFile.scala 75:16:@38799.4]
  assign regs_83_io_reset = reset; // @[RegFile.scala 78:19:@38803.4]
  assign regs_83_io_enable = 1'h1; // @[RegFile.scala 74:20:@38797.4]
  assign regs_84_clock = clock; // @[:@38806.4]
  assign regs_84_reset = io_reset; // @[:@38807.4 RegFile.scala 76:16:@38814.4]
  assign regs_84_io_in = 64'h0; // @[RegFile.scala 75:16:@38813.4]
  assign regs_84_io_reset = reset; // @[RegFile.scala 78:19:@38817.4]
  assign regs_84_io_enable = 1'h1; // @[RegFile.scala 74:20:@38811.4]
  assign regs_85_clock = clock; // @[:@38820.4]
  assign regs_85_reset = io_reset; // @[:@38821.4 RegFile.scala 76:16:@38828.4]
  assign regs_85_io_in = 64'h0; // @[RegFile.scala 75:16:@38827.4]
  assign regs_85_io_reset = reset; // @[RegFile.scala 78:19:@38831.4]
  assign regs_85_io_enable = 1'h1; // @[RegFile.scala 74:20:@38825.4]
  assign regs_86_clock = clock; // @[:@38834.4]
  assign regs_86_reset = io_reset; // @[:@38835.4 RegFile.scala 76:16:@38842.4]
  assign regs_86_io_in = 64'h0; // @[RegFile.scala 75:16:@38841.4]
  assign regs_86_io_reset = reset; // @[RegFile.scala 78:19:@38845.4]
  assign regs_86_io_enable = 1'h1; // @[RegFile.scala 74:20:@38839.4]
  assign regs_87_clock = clock; // @[:@38848.4]
  assign regs_87_reset = io_reset; // @[:@38849.4 RegFile.scala 76:16:@38856.4]
  assign regs_87_io_in = 64'h0; // @[RegFile.scala 75:16:@38855.4]
  assign regs_87_io_reset = reset; // @[RegFile.scala 78:19:@38859.4]
  assign regs_87_io_enable = 1'h1; // @[RegFile.scala 74:20:@38853.4]
  assign regs_88_clock = clock; // @[:@38862.4]
  assign regs_88_reset = io_reset; // @[:@38863.4 RegFile.scala 76:16:@38870.4]
  assign regs_88_io_in = 64'h0; // @[RegFile.scala 75:16:@38869.4]
  assign regs_88_io_reset = reset; // @[RegFile.scala 78:19:@38873.4]
  assign regs_88_io_enable = 1'h1; // @[RegFile.scala 74:20:@38867.4]
  assign regs_89_clock = clock; // @[:@38876.4]
  assign regs_89_reset = io_reset; // @[:@38877.4 RegFile.scala 76:16:@38884.4]
  assign regs_89_io_in = 64'h0; // @[RegFile.scala 75:16:@38883.4]
  assign regs_89_io_reset = reset; // @[RegFile.scala 78:19:@38887.4]
  assign regs_89_io_enable = 1'h1; // @[RegFile.scala 74:20:@38881.4]
  assign regs_90_clock = clock; // @[:@38890.4]
  assign regs_90_reset = io_reset; // @[:@38891.4 RegFile.scala 76:16:@38898.4]
  assign regs_90_io_in = 64'h0; // @[RegFile.scala 75:16:@38897.4]
  assign regs_90_io_reset = reset; // @[RegFile.scala 78:19:@38901.4]
  assign regs_90_io_enable = 1'h1; // @[RegFile.scala 74:20:@38895.4]
  assign regs_91_clock = clock; // @[:@38904.4]
  assign regs_91_reset = io_reset; // @[:@38905.4 RegFile.scala 76:16:@38912.4]
  assign regs_91_io_in = 64'h0; // @[RegFile.scala 75:16:@38911.4]
  assign regs_91_io_reset = reset; // @[RegFile.scala 78:19:@38915.4]
  assign regs_91_io_enable = 1'h1; // @[RegFile.scala 74:20:@38909.4]
  assign regs_92_clock = clock; // @[:@38918.4]
  assign regs_92_reset = io_reset; // @[:@38919.4 RegFile.scala 76:16:@38926.4]
  assign regs_92_io_in = 64'h0; // @[RegFile.scala 75:16:@38925.4]
  assign regs_92_io_reset = reset; // @[RegFile.scala 78:19:@38929.4]
  assign regs_92_io_enable = 1'h1; // @[RegFile.scala 74:20:@38923.4]
  assign regs_93_clock = clock; // @[:@38932.4]
  assign regs_93_reset = io_reset; // @[:@38933.4 RegFile.scala 76:16:@38940.4]
  assign regs_93_io_in = 64'h0; // @[RegFile.scala 75:16:@38939.4]
  assign regs_93_io_reset = reset; // @[RegFile.scala 78:19:@38943.4]
  assign regs_93_io_enable = 1'h1; // @[RegFile.scala 74:20:@38937.4]
  assign regs_94_clock = clock; // @[:@38946.4]
  assign regs_94_reset = io_reset; // @[:@38947.4 RegFile.scala 76:16:@38954.4]
  assign regs_94_io_in = 64'h0; // @[RegFile.scala 75:16:@38953.4]
  assign regs_94_io_reset = reset; // @[RegFile.scala 78:19:@38957.4]
  assign regs_94_io_enable = 1'h1; // @[RegFile.scala 74:20:@38951.4]
  assign regs_95_clock = clock; // @[:@38960.4]
  assign regs_95_reset = io_reset; // @[:@38961.4 RegFile.scala 76:16:@38968.4]
  assign regs_95_io_in = 64'h0; // @[RegFile.scala 75:16:@38967.4]
  assign regs_95_io_reset = reset; // @[RegFile.scala 78:19:@38971.4]
  assign regs_95_io_enable = 1'h1; // @[RegFile.scala 74:20:@38965.4]
  assign regs_96_clock = clock; // @[:@38974.4]
  assign regs_96_reset = io_reset; // @[:@38975.4 RegFile.scala 76:16:@38982.4]
  assign regs_96_io_in = 64'h0; // @[RegFile.scala 75:16:@38981.4]
  assign regs_96_io_reset = reset; // @[RegFile.scala 78:19:@38985.4]
  assign regs_96_io_enable = 1'h1; // @[RegFile.scala 74:20:@38979.4]
  assign regs_97_clock = clock; // @[:@38988.4]
  assign regs_97_reset = io_reset; // @[:@38989.4 RegFile.scala 76:16:@38996.4]
  assign regs_97_io_in = 64'h0; // @[RegFile.scala 75:16:@38995.4]
  assign regs_97_io_reset = reset; // @[RegFile.scala 78:19:@38999.4]
  assign regs_97_io_enable = 1'h1; // @[RegFile.scala 74:20:@38993.4]
  assign regs_98_clock = clock; // @[:@39002.4]
  assign regs_98_reset = io_reset; // @[:@39003.4 RegFile.scala 76:16:@39010.4]
  assign regs_98_io_in = 64'h0; // @[RegFile.scala 75:16:@39009.4]
  assign regs_98_io_reset = reset; // @[RegFile.scala 78:19:@39013.4]
  assign regs_98_io_enable = 1'h1; // @[RegFile.scala 74:20:@39007.4]
  assign regs_99_clock = clock; // @[:@39016.4]
  assign regs_99_reset = io_reset; // @[:@39017.4 RegFile.scala 76:16:@39024.4]
  assign regs_99_io_in = 64'h0; // @[RegFile.scala 75:16:@39023.4]
  assign regs_99_io_reset = reset; // @[RegFile.scala 78:19:@39027.4]
  assign regs_99_io_enable = 1'h1; // @[RegFile.scala 74:20:@39021.4]
  assign regs_100_clock = clock; // @[:@39030.4]
  assign regs_100_reset = io_reset; // @[:@39031.4 RegFile.scala 76:16:@39038.4]
  assign regs_100_io_in = 64'h0; // @[RegFile.scala 75:16:@39037.4]
  assign regs_100_io_reset = reset; // @[RegFile.scala 78:19:@39041.4]
  assign regs_100_io_enable = 1'h1; // @[RegFile.scala 74:20:@39035.4]
  assign regs_101_clock = clock; // @[:@39044.4]
  assign regs_101_reset = io_reset; // @[:@39045.4 RegFile.scala 76:16:@39052.4]
  assign regs_101_io_in = 64'h0; // @[RegFile.scala 75:16:@39051.4]
  assign regs_101_io_reset = reset; // @[RegFile.scala 78:19:@39055.4]
  assign regs_101_io_enable = 1'h1; // @[RegFile.scala 74:20:@39049.4]
  assign regs_102_clock = clock; // @[:@39058.4]
  assign regs_102_reset = io_reset; // @[:@39059.4 RegFile.scala 76:16:@39066.4]
  assign regs_102_io_in = 64'h0; // @[RegFile.scala 75:16:@39065.4]
  assign regs_102_io_reset = reset; // @[RegFile.scala 78:19:@39069.4]
  assign regs_102_io_enable = 1'h1; // @[RegFile.scala 74:20:@39063.4]
  assign regs_103_clock = clock; // @[:@39072.4]
  assign regs_103_reset = io_reset; // @[:@39073.4 RegFile.scala 76:16:@39080.4]
  assign regs_103_io_in = 64'h0; // @[RegFile.scala 75:16:@39079.4]
  assign regs_103_io_reset = reset; // @[RegFile.scala 78:19:@39083.4]
  assign regs_103_io_enable = 1'h1; // @[RegFile.scala 74:20:@39077.4]
  assign regs_104_clock = clock; // @[:@39086.4]
  assign regs_104_reset = io_reset; // @[:@39087.4 RegFile.scala 76:16:@39094.4]
  assign regs_104_io_in = 64'h0; // @[RegFile.scala 75:16:@39093.4]
  assign regs_104_io_reset = reset; // @[RegFile.scala 78:19:@39097.4]
  assign regs_104_io_enable = 1'h1; // @[RegFile.scala 74:20:@39091.4]
  assign regs_105_clock = clock; // @[:@39100.4]
  assign regs_105_reset = io_reset; // @[:@39101.4 RegFile.scala 76:16:@39108.4]
  assign regs_105_io_in = 64'h0; // @[RegFile.scala 75:16:@39107.4]
  assign regs_105_io_reset = reset; // @[RegFile.scala 78:19:@39111.4]
  assign regs_105_io_enable = 1'h1; // @[RegFile.scala 74:20:@39105.4]
  assign regs_106_clock = clock; // @[:@39114.4]
  assign regs_106_reset = io_reset; // @[:@39115.4 RegFile.scala 76:16:@39122.4]
  assign regs_106_io_in = 64'h0; // @[RegFile.scala 75:16:@39121.4]
  assign regs_106_io_reset = reset; // @[RegFile.scala 78:19:@39125.4]
  assign regs_106_io_enable = 1'h1; // @[RegFile.scala 74:20:@39119.4]
  assign regs_107_clock = clock; // @[:@39128.4]
  assign regs_107_reset = io_reset; // @[:@39129.4 RegFile.scala 76:16:@39136.4]
  assign regs_107_io_in = 64'h0; // @[RegFile.scala 75:16:@39135.4]
  assign regs_107_io_reset = reset; // @[RegFile.scala 78:19:@39139.4]
  assign regs_107_io_enable = 1'h1; // @[RegFile.scala 74:20:@39133.4]
  assign regs_108_clock = clock; // @[:@39142.4]
  assign regs_108_reset = io_reset; // @[:@39143.4 RegFile.scala 76:16:@39150.4]
  assign regs_108_io_in = 64'h0; // @[RegFile.scala 75:16:@39149.4]
  assign regs_108_io_reset = reset; // @[RegFile.scala 78:19:@39153.4]
  assign regs_108_io_enable = 1'h1; // @[RegFile.scala 74:20:@39147.4]
  assign regs_109_clock = clock; // @[:@39156.4]
  assign regs_109_reset = io_reset; // @[:@39157.4 RegFile.scala 76:16:@39164.4]
  assign regs_109_io_in = 64'h0; // @[RegFile.scala 75:16:@39163.4]
  assign regs_109_io_reset = reset; // @[RegFile.scala 78:19:@39167.4]
  assign regs_109_io_enable = 1'h1; // @[RegFile.scala 74:20:@39161.4]
  assign regs_110_clock = clock; // @[:@39170.4]
  assign regs_110_reset = io_reset; // @[:@39171.4 RegFile.scala 76:16:@39178.4]
  assign regs_110_io_in = 64'h0; // @[RegFile.scala 75:16:@39177.4]
  assign regs_110_io_reset = reset; // @[RegFile.scala 78:19:@39181.4]
  assign regs_110_io_enable = 1'h1; // @[RegFile.scala 74:20:@39175.4]
  assign regs_111_clock = clock; // @[:@39184.4]
  assign regs_111_reset = io_reset; // @[:@39185.4 RegFile.scala 76:16:@39192.4]
  assign regs_111_io_in = 64'h0; // @[RegFile.scala 75:16:@39191.4]
  assign regs_111_io_reset = reset; // @[RegFile.scala 78:19:@39195.4]
  assign regs_111_io_enable = 1'h1; // @[RegFile.scala 74:20:@39189.4]
  assign regs_112_clock = clock; // @[:@39198.4]
  assign regs_112_reset = io_reset; // @[:@39199.4 RegFile.scala 76:16:@39206.4]
  assign regs_112_io_in = 64'h0; // @[RegFile.scala 75:16:@39205.4]
  assign regs_112_io_reset = reset; // @[RegFile.scala 78:19:@39209.4]
  assign regs_112_io_enable = 1'h1; // @[RegFile.scala 74:20:@39203.4]
  assign regs_113_clock = clock; // @[:@39212.4]
  assign regs_113_reset = io_reset; // @[:@39213.4 RegFile.scala 76:16:@39220.4]
  assign regs_113_io_in = 64'h0; // @[RegFile.scala 75:16:@39219.4]
  assign regs_113_io_reset = reset; // @[RegFile.scala 78:19:@39223.4]
  assign regs_113_io_enable = 1'h1; // @[RegFile.scala 74:20:@39217.4]
  assign regs_114_clock = clock; // @[:@39226.4]
  assign regs_114_reset = io_reset; // @[:@39227.4 RegFile.scala 76:16:@39234.4]
  assign regs_114_io_in = 64'h0; // @[RegFile.scala 75:16:@39233.4]
  assign regs_114_io_reset = reset; // @[RegFile.scala 78:19:@39237.4]
  assign regs_114_io_enable = 1'h1; // @[RegFile.scala 74:20:@39231.4]
  assign regs_115_clock = clock; // @[:@39240.4]
  assign regs_115_reset = io_reset; // @[:@39241.4 RegFile.scala 76:16:@39248.4]
  assign regs_115_io_in = 64'h0; // @[RegFile.scala 75:16:@39247.4]
  assign regs_115_io_reset = reset; // @[RegFile.scala 78:19:@39251.4]
  assign regs_115_io_enable = 1'h1; // @[RegFile.scala 74:20:@39245.4]
  assign regs_116_clock = clock; // @[:@39254.4]
  assign regs_116_reset = io_reset; // @[:@39255.4 RegFile.scala 76:16:@39262.4]
  assign regs_116_io_in = 64'h0; // @[RegFile.scala 75:16:@39261.4]
  assign regs_116_io_reset = reset; // @[RegFile.scala 78:19:@39265.4]
  assign regs_116_io_enable = 1'h1; // @[RegFile.scala 74:20:@39259.4]
  assign regs_117_clock = clock; // @[:@39268.4]
  assign regs_117_reset = io_reset; // @[:@39269.4 RegFile.scala 76:16:@39276.4]
  assign regs_117_io_in = 64'h0; // @[RegFile.scala 75:16:@39275.4]
  assign regs_117_io_reset = reset; // @[RegFile.scala 78:19:@39279.4]
  assign regs_117_io_enable = 1'h1; // @[RegFile.scala 74:20:@39273.4]
  assign regs_118_clock = clock; // @[:@39282.4]
  assign regs_118_reset = io_reset; // @[:@39283.4 RegFile.scala 76:16:@39290.4]
  assign regs_118_io_in = 64'h0; // @[RegFile.scala 75:16:@39289.4]
  assign regs_118_io_reset = reset; // @[RegFile.scala 78:19:@39293.4]
  assign regs_118_io_enable = 1'h1; // @[RegFile.scala 74:20:@39287.4]
  assign regs_119_clock = clock; // @[:@39296.4]
  assign regs_119_reset = io_reset; // @[:@39297.4 RegFile.scala 76:16:@39304.4]
  assign regs_119_io_in = 64'h0; // @[RegFile.scala 75:16:@39303.4]
  assign regs_119_io_reset = reset; // @[RegFile.scala 78:19:@39307.4]
  assign regs_119_io_enable = 1'h1; // @[RegFile.scala 74:20:@39301.4]
  assign regs_120_clock = clock; // @[:@39310.4]
  assign regs_120_reset = io_reset; // @[:@39311.4 RegFile.scala 76:16:@39318.4]
  assign regs_120_io_in = 64'h0; // @[RegFile.scala 75:16:@39317.4]
  assign regs_120_io_reset = reset; // @[RegFile.scala 78:19:@39321.4]
  assign regs_120_io_enable = 1'h1; // @[RegFile.scala 74:20:@39315.4]
  assign regs_121_clock = clock; // @[:@39324.4]
  assign regs_121_reset = io_reset; // @[:@39325.4 RegFile.scala 76:16:@39332.4]
  assign regs_121_io_in = 64'h0; // @[RegFile.scala 75:16:@39331.4]
  assign regs_121_io_reset = reset; // @[RegFile.scala 78:19:@39335.4]
  assign regs_121_io_enable = 1'h1; // @[RegFile.scala 74:20:@39329.4]
  assign regs_122_clock = clock; // @[:@39338.4]
  assign regs_122_reset = io_reset; // @[:@39339.4 RegFile.scala 76:16:@39346.4]
  assign regs_122_io_in = 64'h0; // @[RegFile.scala 75:16:@39345.4]
  assign regs_122_io_reset = reset; // @[RegFile.scala 78:19:@39349.4]
  assign regs_122_io_enable = 1'h1; // @[RegFile.scala 74:20:@39343.4]
  assign regs_123_clock = clock; // @[:@39352.4]
  assign regs_123_reset = io_reset; // @[:@39353.4 RegFile.scala 76:16:@39360.4]
  assign regs_123_io_in = 64'h0; // @[RegFile.scala 75:16:@39359.4]
  assign regs_123_io_reset = reset; // @[RegFile.scala 78:19:@39363.4]
  assign regs_123_io_enable = 1'h1; // @[RegFile.scala 74:20:@39357.4]
  assign regs_124_clock = clock; // @[:@39366.4]
  assign regs_124_reset = io_reset; // @[:@39367.4 RegFile.scala 76:16:@39374.4]
  assign regs_124_io_in = 64'h0; // @[RegFile.scala 75:16:@39373.4]
  assign regs_124_io_reset = reset; // @[RegFile.scala 78:19:@39377.4]
  assign regs_124_io_enable = 1'h1; // @[RegFile.scala 74:20:@39371.4]
  assign regs_125_clock = clock; // @[:@39380.4]
  assign regs_125_reset = io_reset; // @[:@39381.4 RegFile.scala 76:16:@39388.4]
  assign regs_125_io_in = 64'h0; // @[RegFile.scala 75:16:@39387.4]
  assign regs_125_io_reset = reset; // @[RegFile.scala 78:19:@39391.4]
  assign regs_125_io_enable = 1'h1; // @[RegFile.scala 74:20:@39385.4]
  assign regs_126_clock = clock; // @[:@39394.4]
  assign regs_126_reset = io_reset; // @[:@39395.4 RegFile.scala 76:16:@39402.4]
  assign regs_126_io_in = 64'h0; // @[RegFile.scala 75:16:@39401.4]
  assign regs_126_io_reset = reset; // @[RegFile.scala 78:19:@39405.4]
  assign regs_126_io_enable = 1'h1; // @[RegFile.scala 74:20:@39399.4]
  assign regs_127_clock = clock; // @[:@39408.4]
  assign regs_127_reset = io_reset; // @[:@39409.4 RegFile.scala 76:16:@39416.4]
  assign regs_127_io_in = 64'h0; // @[RegFile.scala 75:16:@39415.4]
  assign regs_127_io_reset = reset; // @[RegFile.scala 78:19:@39419.4]
  assign regs_127_io_enable = 1'h1; // @[RegFile.scala 74:20:@39413.4]
  assign regs_128_clock = clock; // @[:@39422.4]
  assign regs_128_reset = io_reset; // @[:@39423.4 RegFile.scala 76:16:@39430.4]
  assign regs_128_io_in = 64'h0; // @[RegFile.scala 75:16:@39429.4]
  assign regs_128_io_reset = reset; // @[RegFile.scala 78:19:@39433.4]
  assign regs_128_io_enable = 1'h1; // @[RegFile.scala 74:20:@39427.4]
  assign regs_129_clock = clock; // @[:@39436.4]
  assign regs_129_reset = io_reset; // @[:@39437.4 RegFile.scala 76:16:@39444.4]
  assign regs_129_io_in = 64'h0; // @[RegFile.scala 75:16:@39443.4]
  assign regs_129_io_reset = reset; // @[RegFile.scala 78:19:@39447.4]
  assign regs_129_io_enable = 1'h1; // @[RegFile.scala 74:20:@39441.4]
  assign regs_130_clock = clock; // @[:@39450.4]
  assign regs_130_reset = io_reset; // @[:@39451.4 RegFile.scala 76:16:@39458.4]
  assign regs_130_io_in = 64'h0; // @[RegFile.scala 75:16:@39457.4]
  assign regs_130_io_reset = reset; // @[RegFile.scala 78:19:@39461.4]
  assign regs_130_io_enable = 1'h1; // @[RegFile.scala 74:20:@39455.4]
  assign regs_131_clock = clock; // @[:@39464.4]
  assign regs_131_reset = io_reset; // @[:@39465.4 RegFile.scala 76:16:@39472.4]
  assign regs_131_io_in = 64'h0; // @[RegFile.scala 75:16:@39471.4]
  assign regs_131_io_reset = reset; // @[RegFile.scala 78:19:@39475.4]
  assign regs_131_io_enable = 1'h1; // @[RegFile.scala 74:20:@39469.4]
  assign regs_132_clock = clock; // @[:@39478.4]
  assign regs_132_reset = io_reset; // @[:@39479.4 RegFile.scala 76:16:@39486.4]
  assign regs_132_io_in = 64'h0; // @[RegFile.scala 75:16:@39485.4]
  assign regs_132_io_reset = reset; // @[RegFile.scala 78:19:@39489.4]
  assign regs_132_io_enable = 1'h1; // @[RegFile.scala 74:20:@39483.4]
  assign regs_133_clock = clock; // @[:@39492.4]
  assign regs_133_reset = io_reset; // @[:@39493.4 RegFile.scala 76:16:@39500.4]
  assign regs_133_io_in = 64'h0; // @[RegFile.scala 75:16:@39499.4]
  assign regs_133_io_reset = reset; // @[RegFile.scala 78:19:@39503.4]
  assign regs_133_io_enable = 1'h1; // @[RegFile.scala 74:20:@39497.4]
  assign regs_134_clock = clock; // @[:@39506.4]
  assign regs_134_reset = io_reset; // @[:@39507.4 RegFile.scala 76:16:@39514.4]
  assign regs_134_io_in = 64'h0; // @[RegFile.scala 75:16:@39513.4]
  assign regs_134_io_reset = reset; // @[RegFile.scala 78:19:@39517.4]
  assign regs_134_io_enable = 1'h1; // @[RegFile.scala 74:20:@39511.4]
  assign regs_135_clock = clock; // @[:@39520.4]
  assign regs_135_reset = io_reset; // @[:@39521.4 RegFile.scala 76:16:@39528.4]
  assign regs_135_io_in = 64'h0; // @[RegFile.scala 75:16:@39527.4]
  assign regs_135_io_reset = reset; // @[RegFile.scala 78:19:@39531.4]
  assign regs_135_io_enable = 1'h1; // @[RegFile.scala 74:20:@39525.4]
  assign regs_136_clock = clock; // @[:@39534.4]
  assign regs_136_reset = io_reset; // @[:@39535.4 RegFile.scala 76:16:@39542.4]
  assign regs_136_io_in = 64'h0; // @[RegFile.scala 75:16:@39541.4]
  assign regs_136_io_reset = reset; // @[RegFile.scala 78:19:@39545.4]
  assign regs_136_io_enable = 1'h1; // @[RegFile.scala 74:20:@39539.4]
  assign regs_137_clock = clock; // @[:@39548.4]
  assign regs_137_reset = io_reset; // @[:@39549.4 RegFile.scala 76:16:@39556.4]
  assign regs_137_io_in = 64'h0; // @[RegFile.scala 75:16:@39555.4]
  assign regs_137_io_reset = reset; // @[RegFile.scala 78:19:@39559.4]
  assign regs_137_io_enable = 1'h1; // @[RegFile.scala 74:20:@39553.4]
  assign regs_138_clock = clock; // @[:@39562.4]
  assign regs_138_reset = io_reset; // @[:@39563.4 RegFile.scala 76:16:@39570.4]
  assign regs_138_io_in = 64'h0; // @[RegFile.scala 75:16:@39569.4]
  assign regs_138_io_reset = reset; // @[RegFile.scala 78:19:@39573.4]
  assign regs_138_io_enable = 1'h1; // @[RegFile.scala 74:20:@39567.4]
  assign regs_139_clock = clock; // @[:@39576.4]
  assign regs_139_reset = io_reset; // @[:@39577.4 RegFile.scala 76:16:@39584.4]
  assign regs_139_io_in = 64'h0; // @[RegFile.scala 75:16:@39583.4]
  assign regs_139_io_reset = reset; // @[RegFile.scala 78:19:@39587.4]
  assign regs_139_io_enable = 1'h1; // @[RegFile.scala 74:20:@39581.4]
  assign regs_140_clock = clock; // @[:@39590.4]
  assign regs_140_reset = io_reset; // @[:@39591.4 RegFile.scala 76:16:@39598.4]
  assign regs_140_io_in = 64'h0; // @[RegFile.scala 75:16:@39597.4]
  assign regs_140_io_reset = reset; // @[RegFile.scala 78:19:@39601.4]
  assign regs_140_io_enable = 1'h1; // @[RegFile.scala 74:20:@39595.4]
  assign regs_141_clock = clock; // @[:@39604.4]
  assign regs_141_reset = io_reset; // @[:@39605.4 RegFile.scala 76:16:@39612.4]
  assign regs_141_io_in = 64'h0; // @[RegFile.scala 75:16:@39611.4]
  assign regs_141_io_reset = reset; // @[RegFile.scala 78:19:@39615.4]
  assign regs_141_io_enable = 1'h1; // @[RegFile.scala 74:20:@39609.4]
  assign regs_142_clock = clock; // @[:@39618.4]
  assign regs_142_reset = io_reset; // @[:@39619.4 RegFile.scala 76:16:@39626.4]
  assign regs_142_io_in = 64'h0; // @[RegFile.scala 75:16:@39625.4]
  assign regs_142_io_reset = reset; // @[RegFile.scala 78:19:@39629.4]
  assign regs_142_io_enable = 1'h1; // @[RegFile.scala 74:20:@39623.4]
  assign regs_143_clock = clock; // @[:@39632.4]
  assign regs_143_reset = io_reset; // @[:@39633.4 RegFile.scala 76:16:@39640.4]
  assign regs_143_io_in = 64'h0; // @[RegFile.scala 75:16:@39639.4]
  assign regs_143_io_reset = reset; // @[RegFile.scala 78:19:@39643.4]
  assign regs_143_io_enable = 1'h1; // @[RegFile.scala 74:20:@39637.4]
  assign regs_144_clock = clock; // @[:@39646.4]
  assign regs_144_reset = io_reset; // @[:@39647.4 RegFile.scala 76:16:@39654.4]
  assign regs_144_io_in = 64'h0; // @[RegFile.scala 75:16:@39653.4]
  assign regs_144_io_reset = reset; // @[RegFile.scala 78:19:@39657.4]
  assign regs_144_io_enable = 1'h1; // @[RegFile.scala 74:20:@39651.4]
  assign regs_145_clock = clock; // @[:@39660.4]
  assign regs_145_reset = io_reset; // @[:@39661.4 RegFile.scala 76:16:@39668.4]
  assign regs_145_io_in = 64'h0; // @[RegFile.scala 75:16:@39667.4]
  assign regs_145_io_reset = reset; // @[RegFile.scala 78:19:@39671.4]
  assign regs_145_io_enable = 1'h1; // @[RegFile.scala 74:20:@39665.4]
  assign regs_146_clock = clock; // @[:@39674.4]
  assign regs_146_reset = io_reset; // @[:@39675.4 RegFile.scala 76:16:@39682.4]
  assign regs_146_io_in = 64'h0; // @[RegFile.scala 75:16:@39681.4]
  assign regs_146_io_reset = reset; // @[RegFile.scala 78:19:@39685.4]
  assign regs_146_io_enable = 1'h1; // @[RegFile.scala 74:20:@39679.4]
  assign regs_147_clock = clock; // @[:@39688.4]
  assign regs_147_reset = io_reset; // @[:@39689.4 RegFile.scala 76:16:@39696.4]
  assign regs_147_io_in = 64'h0; // @[RegFile.scala 75:16:@39695.4]
  assign regs_147_io_reset = reset; // @[RegFile.scala 78:19:@39699.4]
  assign regs_147_io_enable = 1'h1; // @[RegFile.scala 74:20:@39693.4]
  assign regs_148_clock = clock; // @[:@39702.4]
  assign regs_148_reset = io_reset; // @[:@39703.4 RegFile.scala 76:16:@39710.4]
  assign regs_148_io_in = 64'h0; // @[RegFile.scala 75:16:@39709.4]
  assign regs_148_io_reset = reset; // @[RegFile.scala 78:19:@39713.4]
  assign regs_148_io_enable = 1'h1; // @[RegFile.scala 74:20:@39707.4]
  assign regs_149_clock = clock; // @[:@39716.4]
  assign regs_149_reset = io_reset; // @[:@39717.4 RegFile.scala 76:16:@39724.4]
  assign regs_149_io_in = 64'h0; // @[RegFile.scala 75:16:@39723.4]
  assign regs_149_io_reset = reset; // @[RegFile.scala 78:19:@39727.4]
  assign regs_149_io_enable = 1'h1; // @[RegFile.scala 74:20:@39721.4]
  assign regs_150_clock = clock; // @[:@39730.4]
  assign regs_150_reset = io_reset; // @[:@39731.4 RegFile.scala 76:16:@39738.4]
  assign regs_150_io_in = 64'h0; // @[RegFile.scala 75:16:@39737.4]
  assign regs_150_io_reset = reset; // @[RegFile.scala 78:19:@39741.4]
  assign regs_150_io_enable = 1'h1; // @[RegFile.scala 74:20:@39735.4]
  assign regs_151_clock = clock; // @[:@39744.4]
  assign regs_151_reset = io_reset; // @[:@39745.4 RegFile.scala 76:16:@39752.4]
  assign regs_151_io_in = 64'h0; // @[RegFile.scala 75:16:@39751.4]
  assign regs_151_io_reset = reset; // @[RegFile.scala 78:19:@39755.4]
  assign regs_151_io_enable = 1'h1; // @[RegFile.scala 74:20:@39749.4]
  assign regs_152_clock = clock; // @[:@39758.4]
  assign regs_152_reset = io_reset; // @[:@39759.4 RegFile.scala 76:16:@39766.4]
  assign regs_152_io_in = 64'h0; // @[RegFile.scala 75:16:@39765.4]
  assign regs_152_io_reset = reset; // @[RegFile.scala 78:19:@39769.4]
  assign regs_152_io_enable = 1'h1; // @[RegFile.scala 74:20:@39763.4]
  assign regs_153_clock = clock; // @[:@39772.4]
  assign regs_153_reset = io_reset; // @[:@39773.4 RegFile.scala 76:16:@39780.4]
  assign regs_153_io_in = 64'h0; // @[RegFile.scala 75:16:@39779.4]
  assign regs_153_io_reset = reset; // @[RegFile.scala 78:19:@39783.4]
  assign regs_153_io_enable = 1'h1; // @[RegFile.scala 74:20:@39777.4]
  assign regs_154_clock = clock; // @[:@39786.4]
  assign regs_154_reset = io_reset; // @[:@39787.4 RegFile.scala 76:16:@39794.4]
  assign regs_154_io_in = 64'h0; // @[RegFile.scala 75:16:@39793.4]
  assign regs_154_io_reset = reset; // @[RegFile.scala 78:19:@39797.4]
  assign regs_154_io_enable = 1'h1; // @[RegFile.scala 74:20:@39791.4]
  assign regs_155_clock = clock; // @[:@39800.4]
  assign regs_155_reset = io_reset; // @[:@39801.4 RegFile.scala 76:16:@39808.4]
  assign regs_155_io_in = 64'h0; // @[RegFile.scala 75:16:@39807.4]
  assign regs_155_io_reset = reset; // @[RegFile.scala 78:19:@39811.4]
  assign regs_155_io_enable = 1'h1; // @[RegFile.scala 74:20:@39805.4]
  assign regs_156_clock = clock; // @[:@39814.4]
  assign regs_156_reset = io_reset; // @[:@39815.4 RegFile.scala 76:16:@39822.4]
  assign regs_156_io_in = 64'h0; // @[RegFile.scala 75:16:@39821.4]
  assign regs_156_io_reset = reset; // @[RegFile.scala 78:19:@39825.4]
  assign regs_156_io_enable = 1'h1; // @[RegFile.scala 74:20:@39819.4]
  assign regs_157_clock = clock; // @[:@39828.4]
  assign regs_157_reset = io_reset; // @[:@39829.4 RegFile.scala 76:16:@39836.4]
  assign regs_157_io_in = 64'h0; // @[RegFile.scala 75:16:@39835.4]
  assign regs_157_io_reset = reset; // @[RegFile.scala 78:19:@39839.4]
  assign regs_157_io_enable = 1'h1; // @[RegFile.scala 74:20:@39833.4]
  assign regs_158_clock = clock; // @[:@39842.4]
  assign regs_158_reset = io_reset; // @[:@39843.4 RegFile.scala 76:16:@39850.4]
  assign regs_158_io_in = 64'h0; // @[RegFile.scala 75:16:@39849.4]
  assign regs_158_io_reset = reset; // @[RegFile.scala 78:19:@39853.4]
  assign regs_158_io_enable = 1'h1; // @[RegFile.scala 74:20:@39847.4]
  assign regs_159_clock = clock; // @[:@39856.4]
  assign regs_159_reset = io_reset; // @[:@39857.4 RegFile.scala 76:16:@39864.4]
  assign regs_159_io_in = 64'h0; // @[RegFile.scala 75:16:@39863.4]
  assign regs_159_io_reset = reset; // @[RegFile.scala 78:19:@39867.4]
  assign regs_159_io_enable = 1'h1; // @[RegFile.scala 74:20:@39861.4]
  assign regs_160_clock = clock; // @[:@39870.4]
  assign regs_160_reset = io_reset; // @[:@39871.4 RegFile.scala 76:16:@39878.4]
  assign regs_160_io_in = 64'h0; // @[RegFile.scala 75:16:@39877.4]
  assign regs_160_io_reset = reset; // @[RegFile.scala 78:19:@39881.4]
  assign regs_160_io_enable = 1'h1; // @[RegFile.scala 74:20:@39875.4]
  assign regs_161_clock = clock; // @[:@39884.4]
  assign regs_161_reset = io_reset; // @[:@39885.4 RegFile.scala 76:16:@39892.4]
  assign regs_161_io_in = 64'h0; // @[RegFile.scala 75:16:@39891.4]
  assign regs_161_io_reset = reset; // @[RegFile.scala 78:19:@39895.4]
  assign regs_161_io_enable = 1'h1; // @[RegFile.scala 74:20:@39889.4]
  assign regs_162_clock = clock; // @[:@39898.4]
  assign regs_162_reset = io_reset; // @[:@39899.4 RegFile.scala 76:16:@39906.4]
  assign regs_162_io_in = 64'h0; // @[RegFile.scala 75:16:@39905.4]
  assign regs_162_io_reset = reset; // @[RegFile.scala 78:19:@39909.4]
  assign regs_162_io_enable = 1'h1; // @[RegFile.scala 74:20:@39903.4]
  assign regs_163_clock = clock; // @[:@39912.4]
  assign regs_163_reset = io_reset; // @[:@39913.4 RegFile.scala 76:16:@39920.4]
  assign regs_163_io_in = 64'h0; // @[RegFile.scala 75:16:@39919.4]
  assign regs_163_io_reset = reset; // @[RegFile.scala 78:19:@39923.4]
  assign regs_163_io_enable = 1'h1; // @[RegFile.scala 74:20:@39917.4]
  assign regs_164_clock = clock; // @[:@39926.4]
  assign regs_164_reset = io_reset; // @[:@39927.4 RegFile.scala 76:16:@39934.4]
  assign regs_164_io_in = 64'h0; // @[RegFile.scala 75:16:@39933.4]
  assign regs_164_io_reset = reset; // @[RegFile.scala 78:19:@39937.4]
  assign regs_164_io_enable = 1'h1; // @[RegFile.scala 74:20:@39931.4]
  assign regs_165_clock = clock; // @[:@39940.4]
  assign regs_165_reset = io_reset; // @[:@39941.4 RegFile.scala 76:16:@39948.4]
  assign regs_165_io_in = 64'h0; // @[RegFile.scala 75:16:@39947.4]
  assign regs_165_io_reset = reset; // @[RegFile.scala 78:19:@39951.4]
  assign regs_165_io_enable = 1'h1; // @[RegFile.scala 74:20:@39945.4]
  assign regs_166_clock = clock; // @[:@39954.4]
  assign regs_166_reset = io_reset; // @[:@39955.4 RegFile.scala 76:16:@39962.4]
  assign regs_166_io_in = 64'h0; // @[RegFile.scala 75:16:@39961.4]
  assign regs_166_io_reset = reset; // @[RegFile.scala 78:19:@39965.4]
  assign regs_166_io_enable = 1'h1; // @[RegFile.scala 74:20:@39959.4]
  assign regs_167_clock = clock; // @[:@39968.4]
  assign regs_167_reset = io_reset; // @[:@39969.4 RegFile.scala 76:16:@39976.4]
  assign regs_167_io_in = 64'h0; // @[RegFile.scala 75:16:@39975.4]
  assign regs_167_io_reset = reset; // @[RegFile.scala 78:19:@39979.4]
  assign regs_167_io_enable = 1'h1; // @[RegFile.scala 74:20:@39973.4]
  assign regs_168_clock = clock; // @[:@39982.4]
  assign regs_168_reset = io_reset; // @[:@39983.4 RegFile.scala 76:16:@39990.4]
  assign regs_168_io_in = 64'h0; // @[RegFile.scala 75:16:@39989.4]
  assign regs_168_io_reset = reset; // @[RegFile.scala 78:19:@39993.4]
  assign regs_168_io_enable = 1'h1; // @[RegFile.scala 74:20:@39987.4]
  assign regs_169_clock = clock; // @[:@39996.4]
  assign regs_169_reset = io_reset; // @[:@39997.4 RegFile.scala 76:16:@40004.4]
  assign regs_169_io_in = 64'h0; // @[RegFile.scala 75:16:@40003.4]
  assign regs_169_io_reset = reset; // @[RegFile.scala 78:19:@40007.4]
  assign regs_169_io_enable = 1'h1; // @[RegFile.scala 74:20:@40001.4]
  assign regs_170_clock = clock; // @[:@40010.4]
  assign regs_170_reset = io_reset; // @[:@40011.4 RegFile.scala 76:16:@40018.4]
  assign regs_170_io_in = 64'h0; // @[RegFile.scala 75:16:@40017.4]
  assign regs_170_io_reset = reset; // @[RegFile.scala 78:19:@40021.4]
  assign regs_170_io_enable = 1'h1; // @[RegFile.scala 74:20:@40015.4]
  assign regs_171_clock = clock; // @[:@40024.4]
  assign regs_171_reset = io_reset; // @[:@40025.4 RegFile.scala 76:16:@40032.4]
  assign regs_171_io_in = 64'h0; // @[RegFile.scala 75:16:@40031.4]
  assign regs_171_io_reset = reset; // @[RegFile.scala 78:19:@40035.4]
  assign regs_171_io_enable = 1'h1; // @[RegFile.scala 74:20:@40029.4]
  assign regs_172_clock = clock; // @[:@40038.4]
  assign regs_172_reset = io_reset; // @[:@40039.4 RegFile.scala 76:16:@40046.4]
  assign regs_172_io_in = 64'h0; // @[RegFile.scala 75:16:@40045.4]
  assign regs_172_io_reset = reset; // @[RegFile.scala 78:19:@40049.4]
  assign regs_172_io_enable = 1'h1; // @[RegFile.scala 74:20:@40043.4]
  assign regs_173_clock = clock; // @[:@40052.4]
  assign regs_173_reset = io_reset; // @[:@40053.4 RegFile.scala 76:16:@40060.4]
  assign regs_173_io_in = 64'h0; // @[RegFile.scala 75:16:@40059.4]
  assign regs_173_io_reset = reset; // @[RegFile.scala 78:19:@40063.4]
  assign regs_173_io_enable = 1'h1; // @[RegFile.scala 74:20:@40057.4]
  assign regs_174_clock = clock; // @[:@40066.4]
  assign regs_174_reset = io_reset; // @[:@40067.4 RegFile.scala 76:16:@40074.4]
  assign regs_174_io_in = 64'h0; // @[RegFile.scala 75:16:@40073.4]
  assign regs_174_io_reset = reset; // @[RegFile.scala 78:19:@40077.4]
  assign regs_174_io_enable = 1'h1; // @[RegFile.scala 74:20:@40071.4]
  assign regs_175_clock = clock; // @[:@40080.4]
  assign regs_175_reset = io_reset; // @[:@40081.4 RegFile.scala 76:16:@40088.4]
  assign regs_175_io_in = 64'h0; // @[RegFile.scala 75:16:@40087.4]
  assign regs_175_io_reset = reset; // @[RegFile.scala 78:19:@40091.4]
  assign regs_175_io_enable = 1'h1; // @[RegFile.scala 74:20:@40085.4]
  assign regs_176_clock = clock; // @[:@40094.4]
  assign regs_176_reset = io_reset; // @[:@40095.4 RegFile.scala 76:16:@40102.4]
  assign regs_176_io_in = 64'h0; // @[RegFile.scala 75:16:@40101.4]
  assign regs_176_io_reset = reset; // @[RegFile.scala 78:19:@40105.4]
  assign regs_176_io_enable = 1'h1; // @[RegFile.scala 74:20:@40099.4]
  assign regs_177_clock = clock; // @[:@40108.4]
  assign regs_177_reset = io_reset; // @[:@40109.4 RegFile.scala 76:16:@40116.4]
  assign regs_177_io_in = 64'h0; // @[RegFile.scala 75:16:@40115.4]
  assign regs_177_io_reset = reset; // @[RegFile.scala 78:19:@40119.4]
  assign regs_177_io_enable = 1'h1; // @[RegFile.scala 74:20:@40113.4]
  assign regs_178_clock = clock; // @[:@40122.4]
  assign regs_178_reset = io_reset; // @[:@40123.4 RegFile.scala 76:16:@40130.4]
  assign regs_178_io_in = 64'h0; // @[RegFile.scala 75:16:@40129.4]
  assign regs_178_io_reset = reset; // @[RegFile.scala 78:19:@40133.4]
  assign regs_178_io_enable = 1'h1; // @[RegFile.scala 74:20:@40127.4]
  assign regs_179_clock = clock; // @[:@40136.4]
  assign regs_179_reset = io_reset; // @[:@40137.4 RegFile.scala 76:16:@40144.4]
  assign regs_179_io_in = 64'h0; // @[RegFile.scala 75:16:@40143.4]
  assign regs_179_io_reset = reset; // @[RegFile.scala 78:19:@40147.4]
  assign regs_179_io_enable = 1'h1; // @[RegFile.scala 74:20:@40141.4]
  assign regs_180_clock = clock; // @[:@40150.4]
  assign regs_180_reset = io_reset; // @[:@40151.4 RegFile.scala 76:16:@40158.4]
  assign regs_180_io_in = 64'h0; // @[RegFile.scala 75:16:@40157.4]
  assign regs_180_io_reset = reset; // @[RegFile.scala 78:19:@40161.4]
  assign regs_180_io_enable = 1'h1; // @[RegFile.scala 74:20:@40155.4]
  assign regs_181_clock = clock; // @[:@40164.4]
  assign regs_181_reset = io_reset; // @[:@40165.4 RegFile.scala 76:16:@40172.4]
  assign regs_181_io_in = 64'h0; // @[RegFile.scala 75:16:@40171.4]
  assign regs_181_io_reset = reset; // @[RegFile.scala 78:19:@40175.4]
  assign regs_181_io_enable = 1'h1; // @[RegFile.scala 74:20:@40169.4]
  assign regs_182_clock = clock; // @[:@40178.4]
  assign regs_182_reset = io_reset; // @[:@40179.4 RegFile.scala 76:16:@40186.4]
  assign regs_182_io_in = 64'h0; // @[RegFile.scala 75:16:@40185.4]
  assign regs_182_io_reset = reset; // @[RegFile.scala 78:19:@40189.4]
  assign regs_182_io_enable = 1'h1; // @[RegFile.scala 74:20:@40183.4]
  assign regs_183_clock = clock; // @[:@40192.4]
  assign regs_183_reset = io_reset; // @[:@40193.4 RegFile.scala 76:16:@40200.4]
  assign regs_183_io_in = 64'h0; // @[RegFile.scala 75:16:@40199.4]
  assign regs_183_io_reset = reset; // @[RegFile.scala 78:19:@40203.4]
  assign regs_183_io_enable = 1'h1; // @[RegFile.scala 74:20:@40197.4]
  assign regs_184_clock = clock; // @[:@40206.4]
  assign regs_184_reset = io_reset; // @[:@40207.4 RegFile.scala 76:16:@40214.4]
  assign regs_184_io_in = 64'h0; // @[RegFile.scala 75:16:@40213.4]
  assign regs_184_io_reset = reset; // @[RegFile.scala 78:19:@40217.4]
  assign regs_184_io_enable = 1'h1; // @[RegFile.scala 74:20:@40211.4]
  assign regs_185_clock = clock; // @[:@40220.4]
  assign regs_185_reset = io_reset; // @[:@40221.4 RegFile.scala 76:16:@40228.4]
  assign regs_185_io_in = 64'h0; // @[RegFile.scala 75:16:@40227.4]
  assign regs_185_io_reset = reset; // @[RegFile.scala 78:19:@40231.4]
  assign regs_185_io_enable = 1'h1; // @[RegFile.scala 74:20:@40225.4]
  assign regs_186_clock = clock; // @[:@40234.4]
  assign regs_186_reset = io_reset; // @[:@40235.4 RegFile.scala 76:16:@40242.4]
  assign regs_186_io_in = 64'h0; // @[RegFile.scala 75:16:@40241.4]
  assign regs_186_io_reset = reset; // @[RegFile.scala 78:19:@40245.4]
  assign regs_186_io_enable = 1'h1; // @[RegFile.scala 74:20:@40239.4]
  assign regs_187_clock = clock; // @[:@40248.4]
  assign regs_187_reset = io_reset; // @[:@40249.4 RegFile.scala 76:16:@40256.4]
  assign regs_187_io_in = 64'h0; // @[RegFile.scala 75:16:@40255.4]
  assign regs_187_io_reset = reset; // @[RegFile.scala 78:19:@40259.4]
  assign regs_187_io_enable = 1'h1; // @[RegFile.scala 74:20:@40253.4]
  assign regs_188_clock = clock; // @[:@40262.4]
  assign regs_188_reset = io_reset; // @[:@40263.4 RegFile.scala 76:16:@40270.4]
  assign regs_188_io_in = 64'h0; // @[RegFile.scala 75:16:@40269.4]
  assign regs_188_io_reset = reset; // @[RegFile.scala 78:19:@40273.4]
  assign regs_188_io_enable = 1'h1; // @[RegFile.scala 74:20:@40267.4]
  assign regs_189_clock = clock; // @[:@40276.4]
  assign regs_189_reset = io_reset; // @[:@40277.4 RegFile.scala 76:16:@40284.4]
  assign regs_189_io_in = 64'h0; // @[RegFile.scala 75:16:@40283.4]
  assign regs_189_io_reset = reset; // @[RegFile.scala 78:19:@40287.4]
  assign regs_189_io_enable = 1'h1; // @[RegFile.scala 74:20:@40281.4]
  assign regs_190_clock = clock; // @[:@40290.4]
  assign regs_190_reset = io_reset; // @[:@40291.4 RegFile.scala 76:16:@40298.4]
  assign regs_190_io_in = 64'h0; // @[RegFile.scala 75:16:@40297.4]
  assign regs_190_io_reset = reset; // @[RegFile.scala 78:19:@40301.4]
  assign regs_190_io_enable = 1'h1; // @[RegFile.scala 74:20:@40295.4]
  assign regs_191_clock = clock; // @[:@40304.4]
  assign regs_191_reset = io_reset; // @[:@40305.4 RegFile.scala 76:16:@40312.4]
  assign regs_191_io_in = 64'h0; // @[RegFile.scala 75:16:@40311.4]
  assign regs_191_io_reset = reset; // @[RegFile.scala 78:19:@40315.4]
  assign regs_191_io_enable = 1'h1; // @[RegFile.scala 74:20:@40309.4]
  assign regs_192_clock = clock; // @[:@40318.4]
  assign regs_192_reset = io_reset; // @[:@40319.4 RegFile.scala 76:16:@40326.4]
  assign regs_192_io_in = 64'h0; // @[RegFile.scala 75:16:@40325.4]
  assign regs_192_io_reset = reset; // @[RegFile.scala 78:19:@40329.4]
  assign regs_192_io_enable = 1'h1; // @[RegFile.scala 74:20:@40323.4]
  assign regs_193_clock = clock; // @[:@40332.4]
  assign regs_193_reset = io_reset; // @[:@40333.4 RegFile.scala 76:16:@40340.4]
  assign regs_193_io_in = 64'h0; // @[RegFile.scala 75:16:@40339.4]
  assign regs_193_io_reset = reset; // @[RegFile.scala 78:19:@40343.4]
  assign regs_193_io_enable = 1'h1; // @[RegFile.scala 74:20:@40337.4]
  assign regs_194_clock = clock; // @[:@40346.4]
  assign regs_194_reset = io_reset; // @[:@40347.4 RegFile.scala 76:16:@40354.4]
  assign regs_194_io_in = 64'h0; // @[RegFile.scala 75:16:@40353.4]
  assign regs_194_io_reset = reset; // @[RegFile.scala 78:19:@40357.4]
  assign regs_194_io_enable = 1'h1; // @[RegFile.scala 74:20:@40351.4]
  assign regs_195_clock = clock; // @[:@40360.4]
  assign regs_195_reset = io_reset; // @[:@40361.4 RegFile.scala 76:16:@40368.4]
  assign regs_195_io_in = 64'h0; // @[RegFile.scala 75:16:@40367.4]
  assign regs_195_io_reset = reset; // @[RegFile.scala 78:19:@40371.4]
  assign regs_195_io_enable = 1'h1; // @[RegFile.scala 74:20:@40365.4]
  assign regs_196_clock = clock; // @[:@40374.4]
  assign regs_196_reset = io_reset; // @[:@40375.4 RegFile.scala 76:16:@40382.4]
  assign regs_196_io_in = 64'h0; // @[RegFile.scala 75:16:@40381.4]
  assign regs_196_io_reset = reset; // @[RegFile.scala 78:19:@40385.4]
  assign regs_196_io_enable = 1'h1; // @[RegFile.scala 74:20:@40379.4]
  assign regs_197_clock = clock; // @[:@40388.4]
  assign regs_197_reset = io_reset; // @[:@40389.4 RegFile.scala 76:16:@40396.4]
  assign regs_197_io_in = 64'h0; // @[RegFile.scala 75:16:@40395.4]
  assign regs_197_io_reset = reset; // @[RegFile.scala 78:19:@40399.4]
  assign regs_197_io_enable = 1'h1; // @[RegFile.scala 74:20:@40393.4]
  assign regs_198_clock = clock; // @[:@40402.4]
  assign regs_198_reset = io_reset; // @[:@40403.4 RegFile.scala 76:16:@40410.4]
  assign regs_198_io_in = 64'h0; // @[RegFile.scala 75:16:@40409.4]
  assign regs_198_io_reset = reset; // @[RegFile.scala 78:19:@40413.4]
  assign regs_198_io_enable = 1'h1; // @[RegFile.scala 74:20:@40407.4]
  assign regs_199_clock = clock; // @[:@40416.4]
  assign regs_199_reset = io_reset; // @[:@40417.4 RegFile.scala 76:16:@40424.4]
  assign regs_199_io_in = 64'h0; // @[RegFile.scala 75:16:@40423.4]
  assign regs_199_io_reset = reset; // @[RegFile.scala 78:19:@40427.4]
  assign regs_199_io_enable = 1'h1; // @[RegFile.scala 74:20:@40421.4]
  assign regs_200_clock = clock; // @[:@40430.4]
  assign regs_200_reset = io_reset; // @[:@40431.4 RegFile.scala 76:16:@40438.4]
  assign regs_200_io_in = 64'h0; // @[RegFile.scala 75:16:@40437.4]
  assign regs_200_io_reset = reset; // @[RegFile.scala 78:19:@40441.4]
  assign regs_200_io_enable = 1'h1; // @[RegFile.scala 74:20:@40435.4]
  assign regs_201_clock = clock; // @[:@40444.4]
  assign regs_201_reset = io_reset; // @[:@40445.4 RegFile.scala 76:16:@40452.4]
  assign regs_201_io_in = 64'h0; // @[RegFile.scala 75:16:@40451.4]
  assign regs_201_io_reset = reset; // @[RegFile.scala 78:19:@40455.4]
  assign regs_201_io_enable = 1'h1; // @[RegFile.scala 74:20:@40449.4]
  assign regs_202_clock = clock; // @[:@40458.4]
  assign regs_202_reset = io_reset; // @[:@40459.4 RegFile.scala 76:16:@40466.4]
  assign regs_202_io_in = 64'h0; // @[RegFile.scala 75:16:@40465.4]
  assign regs_202_io_reset = reset; // @[RegFile.scala 78:19:@40469.4]
  assign regs_202_io_enable = 1'h1; // @[RegFile.scala 74:20:@40463.4]
  assign regs_203_clock = clock; // @[:@40472.4]
  assign regs_203_reset = io_reset; // @[:@40473.4 RegFile.scala 76:16:@40480.4]
  assign regs_203_io_in = 64'h0; // @[RegFile.scala 75:16:@40479.4]
  assign regs_203_io_reset = reset; // @[RegFile.scala 78:19:@40483.4]
  assign regs_203_io_enable = 1'h1; // @[RegFile.scala 74:20:@40477.4]
  assign regs_204_clock = clock; // @[:@40486.4]
  assign regs_204_reset = io_reset; // @[:@40487.4 RegFile.scala 76:16:@40494.4]
  assign regs_204_io_in = 64'h0; // @[RegFile.scala 75:16:@40493.4]
  assign regs_204_io_reset = reset; // @[RegFile.scala 78:19:@40497.4]
  assign regs_204_io_enable = 1'h1; // @[RegFile.scala 74:20:@40491.4]
  assign regs_205_clock = clock; // @[:@40500.4]
  assign regs_205_reset = io_reset; // @[:@40501.4 RegFile.scala 76:16:@40508.4]
  assign regs_205_io_in = 64'h0; // @[RegFile.scala 75:16:@40507.4]
  assign regs_205_io_reset = reset; // @[RegFile.scala 78:19:@40511.4]
  assign regs_205_io_enable = 1'h1; // @[RegFile.scala 74:20:@40505.4]
  assign regs_206_clock = clock; // @[:@40514.4]
  assign regs_206_reset = io_reset; // @[:@40515.4 RegFile.scala 76:16:@40522.4]
  assign regs_206_io_in = 64'h0; // @[RegFile.scala 75:16:@40521.4]
  assign regs_206_io_reset = reset; // @[RegFile.scala 78:19:@40525.4]
  assign regs_206_io_enable = 1'h1; // @[RegFile.scala 74:20:@40519.4]
  assign regs_207_clock = clock; // @[:@40528.4]
  assign regs_207_reset = io_reset; // @[:@40529.4 RegFile.scala 76:16:@40536.4]
  assign regs_207_io_in = 64'h0; // @[RegFile.scala 75:16:@40535.4]
  assign regs_207_io_reset = reset; // @[RegFile.scala 78:19:@40539.4]
  assign regs_207_io_enable = 1'h1; // @[RegFile.scala 74:20:@40533.4]
  assign regs_208_clock = clock; // @[:@40542.4]
  assign regs_208_reset = io_reset; // @[:@40543.4 RegFile.scala 76:16:@40550.4]
  assign regs_208_io_in = 64'h0; // @[RegFile.scala 75:16:@40549.4]
  assign regs_208_io_reset = reset; // @[RegFile.scala 78:19:@40553.4]
  assign regs_208_io_enable = 1'h1; // @[RegFile.scala 74:20:@40547.4]
  assign regs_209_clock = clock; // @[:@40556.4]
  assign regs_209_reset = io_reset; // @[:@40557.4 RegFile.scala 76:16:@40564.4]
  assign regs_209_io_in = 64'h0; // @[RegFile.scala 75:16:@40563.4]
  assign regs_209_io_reset = reset; // @[RegFile.scala 78:19:@40567.4]
  assign regs_209_io_enable = 1'h1; // @[RegFile.scala 74:20:@40561.4]
  assign regs_210_clock = clock; // @[:@40570.4]
  assign regs_210_reset = io_reset; // @[:@40571.4 RegFile.scala 76:16:@40578.4]
  assign regs_210_io_in = 64'h0; // @[RegFile.scala 75:16:@40577.4]
  assign regs_210_io_reset = reset; // @[RegFile.scala 78:19:@40581.4]
  assign regs_210_io_enable = 1'h1; // @[RegFile.scala 74:20:@40575.4]
  assign regs_211_clock = clock; // @[:@40584.4]
  assign regs_211_reset = io_reset; // @[:@40585.4 RegFile.scala 76:16:@40592.4]
  assign regs_211_io_in = 64'h0; // @[RegFile.scala 75:16:@40591.4]
  assign regs_211_io_reset = reset; // @[RegFile.scala 78:19:@40595.4]
  assign regs_211_io_enable = 1'h1; // @[RegFile.scala 74:20:@40589.4]
  assign regs_212_clock = clock; // @[:@40598.4]
  assign regs_212_reset = io_reset; // @[:@40599.4 RegFile.scala 76:16:@40606.4]
  assign regs_212_io_in = 64'h0; // @[RegFile.scala 75:16:@40605.4]
  assign regs_212_io_reset = reset; // @[RegFile.scala 78:19:@40609.4]
  assign regs_212_io_enable = 1'h1; // @[RegFile.scala 74:20:@40603.4]
  assign regs_213_clock = clock; // @[:@40612.4]
  assign regs_213_reset = io_reset; // @[:@40613.4 RegFile.scala 76:16:@40620.4]
  assign regs_213_io_in = 64'h0; // @[RegFile.scala 75:16:@40619.4]
  assign regs_213_io_reset = reset; // @[RegFile.scala 78:19:@40623.4]
  assign regs_213_io_enable = 1'h1; // @[RegFile.scala 74:20:@40617.4]
  assign regs_214_clock = clock; // @[:@40626.4]
  assign regs_214_reset = io_reset; // @[:@40627.4 RegFile.scala 76:16:@40634.4]
  assign regs_214_io_in = 64'h0; // @[RegFile.scala 75:16:@40633.4]
  assign regs_214_io_reset = reset; // @[RegFile.scala 78:19:@40637.4]
  assign regs_214_io_enable = 1'h1; // @[RegFile.scala 74:20:@40631.4]
  assign regs_215_clock = clock; // @[:@40640.4]
  assign regs_215_reset = io_reset; // @[:@40641.4 RegFile.scala 76:16:@40648.4]
  assign regs_215_io_in = 64'h0; // @[RegFile.scala 75:16:@40647.4]
  assign regs_215_io_reset = reset; // @[RegFile.scala 78:19:@40651.4]
  assign regs_215_io_enable = 1'h1; // @[RegFile.scala 74:20:@40645.4]
  assign regs_216_clock = clock; // @[:@40654.4]
  assign regs_216_reset = io_reset; // @[:@40655.4 RegFile.scala 76:16:@40662.4]
  assign regs_216_io_in = 64'h0; // @[RegFile.scala 75:16:@40661.4]
  assign regs_216_io_reset = reset; // @[RegFile.scala 78:19:@40665.4]
  assign regs_216_io_enable = 1'h1; // @[RegFile.scala 74:20:@40659.4]
  assign regs_217_clock = clock; // @[:@40668.4]
  assign regs_217_reset = io_reset; // @[:@40669.4 RegFile.scala 76:16:@40676.4]
  assign regs_217_io_in = 64'h0; // @[RegFile.scala 75:16:@40675.4]
  assign regs_217_io_reset = reset; // @[RegFile.scala 78:19:@40679.4]
  assign regs_217_io_enable = 1'h1; // @[RegFile.scala 74:20:@40673.4]
  assign regs_218_clock = clock; // @[:@40682.4]
  assign regs_218_reset = io_reset; // @[:@40683.4 RegFile.scala 76:16:@40690.4]
  assign regs_218_io_in = 64'h0; // @[RegFile.scala 75:16:@40689.4]
  assign regs_218_io_reset = reset; // @[RegFile.scala 78:19:@40693.4]
  assign regs_218_io_enable = 1'h1; // @[RegFile.scala 74:20:@40687.4]
  assign regs_219_clock = clock; // @[:@40696.4]
  assign regs_219_reset = io_reset; // @[:@40697.4 RegFile.scala 76:16:@40704.4]
  assign regs_219_io_in = 64'h0; // @[RegFile.scala 75:16:@40703.4]
  assign regs_219_io_reset = reset; // @[RegFile.scala 78:19:@40707.4]
  assign regs_219_io_enable = 1'h1; // @[RegFile.scala 74:20:@40701.4]
  assign regs_220_clock = clock; // @[:@40710.4]
  assign regs_220_reset = io_reset; // @[:@40711.4 RegFile.scala 76:16:@40718.4]
  assign regs_220_io_in = 64'h0; // @[RegFile.scala 75:16:@40717.4]
  assign regs_220_io_reset = reset; // @[RegFile.scala 78:19:@40721.4]
  assign regs_220_io_enable = 1'h1; // @[RegFile.scala 74:20:@40715.4]
  assign regs_221_clock = clock; // @[:@40724.4]
  assign regs_221_reset = io_reset; // @[:@40725.4 RegFile.scala 76:16:@40732.4]
  assign regs_221_io_in = 64'h0; // @[RegFile.scala 75:16:@40731.4]
  assign regs_221_io_reset = reset; // @[RegFile.scala 78:19:@40735.4]
  assign regs_221_io_enable = 1'h1; // @[RegFile.scala 74:20:@40729.4]
  assign regs_222_clock = clock; // @[:@40738.4]
  assign regs_222_reset = io_reset; // @[:@40739.4 RegFile.scala 76:16:@40746.4]
  assign regs_222_io_in = 64'h0; // @[RegFile.scala 75:16:@40745.4]
  assign regs_222_io_reset = reset; // @[RegFile.scala 78:19:@40749.4]
  assign regs_222_io_enable = 1'h1; // @[RegFile.scala 74:20:@40743.4]
  assign regs_223_clock = clock; // @[:@40752.4]
  assign regs_223_reset = io_reset; // @[:@40753.4 RegFile.scala 76:16:@40760.4]
  assign regs_223_io_in = 64'h0; // @[RegFile.scala 75:16:@40759.4]
  assign regs_223_io_reset = reset; // @[RegFile.scala 78:19:@40763.4]
  assign regs_223_io_enable = 1'h1; // @[RegFile.scala 74:20:@40757.4]
  assign regs_224_clock = clock; // @[:@40766.4]
  assign regs_224_reset = io_reset; // @[:@40767.4 RegFile.scala 76:16:@40774.4]
  assign regs_224_io_in = 64'h0; // @[RegFile.scala 75:16:@40773.4]
  assign regs_224_io_reset = reset; // @[RegFile.scala 78:19:@40777.4]
  assign regs_224_io_enable = 1'h1; // @[RegFile.scala 74:20:@40771.4]
  assign regs_225_clock = clock; // @[:@40780.4]
  assign regs_225_reset = io_reset; // @[:@40781.4 RegFile.scala 76:16:@40788.4]
  assign regs_225_io_in = 64'h0; // @[RegFile.scala 75:16:@40787.4]
  assign regs_225_io_reset = reset; // @[RegFile.scala 78:19:@40791.4]
  assign regs_225_io_enable = 1'h1; // @[RegFile.scala 74:20:@40785.4]
  assign regs_226_clock = clock; // @[:@40794.4]
  assign regs_226_reset = io_reset; // @[:@40795.4 RegFile.scala 76:16:@40802.4]
  assign regs_226_io_in = 64'h0; // @[RegFile.scala 75:16:@40801.4]
  assign regs_226_io_reset = reset; // @[RegFile.scala 78:19:@40805.4]
  assign regs_226_io_enable = 1'h1; // @[RegFile.scala 74:20:@40799.4]
  assign regs_227_clock = clock; // @[:@40808.4]
  assign regs_227_reset = io_reset; // @[:@40809.4 RegFile.scala 76:16:@40816.4]
  assign regs_227_io_in = 64'h0; // @[RegFile.scala 75:16:@40815.4]
  assign regs_227_io_reset = reset; // @[RegFile.scala 78:19:@40819.4]
  assign regs_227_io_enable = 1'h1; // @[RegFile.scala 74:20:@40813.4]
  assign regs_228_clock = clock; // @[:@40822.4]
  assign regs_228_reset = io_reset; // @[:@40823.4 RegFile.scala 76:16:@40830.4]
  assign regs_228_io_in = 64'h0; // @[RegFile.scala 75:16:@40829.4]
  assign regs_228_io_reset = reset; // @[RegFile.scala 78:19:@40833.4]
  assign regs_228_io_enable = 1'h1; // @[RegFile.scala 74:20:@40827.4]
  assign regs_229_clock = clock; // @[:@40836.4]
  assign regs_229_reset = io_reset; // @[:@40837.4 RegFile.scala 76:16:@40844.4]
  assign regs_229_io_in = 64'h0; // @[RegFile.scala 75:16:@40843.4]
  assign regs_229_io_reset = reset; // @[RegFile.scala 78:19:@40847.4]
  assign regs_229_io_enable = 1'h1; // @[RegFile.scala 74:20:@40841.4]
  assign regs_230_clock = clock; // @[:@40850.4]
  assign regs_230_reset = io_reset; // @[:@40851.4 RegFile.scala 76:16:@40858.4]
  assign regs_230_io_in = 64'h0; // @[RegFile.scala 75:16:@40857.4]
  assign regs_230_io_reset = reset; // @[RegFile.scala 78:19:@40861.4]
  assign regs_230_io_enable = 1'h1; // @[RegFile.scala 74:20:@40855.4]
  assign regs_231_clock = clock; // @[:@40864.4]
  assign regs_231_reset = io_reset; // @[:@40865.4 RegFile.scala 76:16:@40872.4]
  assign regs_231_io_in = 64'h0; // @[RegFile.scala 75:16:@40871.4]
  assign regs_231_io_reset = reset; // @[RegFile.scala 78:19:@40875.4]
  assign regs_231_io_enable = 1'h1; // @[RegFile.scala 74:20:@40869.4]
  assign regs_232_clock = clock; // @[:@40878.4]
  assign regs_232_reset = io_reset; // @[:@40879.4 RegFile.scala 76:16:@40886.4]
  assign regs_232_io_in = 64'h0; // @[RegFile.scala 75:16:@40885.4]
  assign regs_232_io_reset = reset; // @[RegFile.scala 78:19:@40889.4]
  assign regs_232_io_enable = 1'h1; // @[RegFile.scala 74:20:@40883.4]
  assign regs_233_clock = clock; // @[:@40892.4]
  assign regs_233_reset = io_reset; // @[:@40893.4 RegFile.scala 76:16:@40900.4]
  assign regs_233_io_in = 64'h0; // @[RegFile.scala 75:16:@40899.4]
  assign regs_233_io_reset = reset; // @[RegFile.scala 78:19:@40903.4]
  assign regs_233_io_enable = 1'h1; // @[RegFile.scala 74:20:@40897.4]
  assign regs_234_clock = clock; // @[:@40906.4]
  assign regs_234_reset = io_reset; // @[:@40907.4 RegFile.scala 76:16:@40914.4]
  assign regs_234_io_in = 64'h0; // @[RegFile.scala 75:16:@40913.4]
  assign regs_234_io_reset = reset; // @[RegFile.scala 78:19:@40917.4]
  assign regs_234_io_enable = 1'h1; // @[RegFile.scala 74:20:@40911.4]
  assign regs_235_clock = clock; // @[:@40920.4]
  assign regs_235_reset = io_reset; // @[:@40921.4 RegFile.scala 76:16:@40928.4]
  assign regs_235_io_in = 64'h0; // @[RegFile.scala 75:16:@40927.4]
  assign regs_235_io_reset = reset; // @[RegFile.scala 78:19:@40931.4]
  assign regs_235_io_enable = 1'h1; // @[RegFile.scala 74:20:@40925.4]
  assign regs_236_clock = clock; // @[:@40934.4]
  assign regs_236_reset = io_reset; // @[:@40935.4 RegFile.scala 76:16:@40942.4]
  assign regs_236_io_in = 64'h0; // @[RegFile.scala 75:16:@40941.4]
  assign regs_236_io_reset = reset; // @[RegFile.scala 78:19:@40945.4]
  assign regs_236_io_enable = 1'h1; // @[RegFile.scala 74:20:@40939.4]
  assign regs_237_clock = clock; // @[:@40948.4]
  assign regs_237_reset = io_reset; // @[:@40949.4 RegFile.scala 76:16:@40956.4]
  assign regs_237_io_in = 64'h0; // @[RegFile.scala 75:16:@40955.4]
  assign regs_237_io_reset = reset; // @[RegFile.scala 78:19:@40959.4]
  assign regs_237_io_enable = 1'h1; // @[RegFile.scala 74:20:@40953.4]
  assign regs_238_clock = clock; // @[:@40962.4]
  assign regs_238_reset = io_reset; // @[:@40963.4 RegFile.scala 76:16:@40970.4]
  assign regs_238_io_in = 64'h0; // @[RegFile.scala 75:16:@40969.4]
  assign regs_238_io_reset = reset; // @[RegFile.scala 78:19:@40973.4]
  assign regs_238_io_enable = 1'h1; // @[RegFile.scala 74:20:@40967.4]
  assign regs_239_clock = clock; // @[:@40976.4]
  assign regs_239_reset = io_reset; // @[:@40977.4 RegFile.scala 76:16:@40984.4]
  assign regs_239_io_in = 64'h0; // @[RegFile.scala 75:16:@40983.4]
  assign regs_239_io_reset = reset; // @[RegFile.scala 78:19:@40987.4]
  assign regs_239_io_enable = 1'h1; // @[RegFile.scala 74:20:@40981.4]
  assign regs_240_clock = clock; // @[:@40990.4]
  assign regs_240_reset = io_reset; // @[:@40991.4 RegFile.scala 76:16:@40998.4]
  assign regs_240_io_in = 64'h0; // @[RegFile.scala 75:16:@40997.4]
  assign regs_240_io_reset = reset; // @[RegFile.scala 78:19:@41001.4]
  assign regs_240_io_enable = 1'h1; // @[RegFile.scala 74:20:@40995.4]
  assign regs_241_clock = clock; // @[:@41004.4]
  assign regs_241_reset = io_reset; // @[:@41005.4 RegFile.scala 76:16:@41012.4]
  assign regs_241_io_in = 64'h0; // @[RegFile.scala 75:16:@41011.4]
  assign regs_241_io_reset = reset; // @[RegFile.scala 78:19:@41015.4]
  assign regs_241_io_enable = 1'h1; // @[RegFile.scala 74:20:@41009.4]
  assign regs_242_clock = clock; // @[:@41018.4]
  assign regs_242_reset = io_reset; // @[:@41019.4 RegFile.scala 76:16:@41026.4]
  assign regs_242_io_in = 64'h0; // @[RegFile.scala 75:16:@41025.4]
  assign regs_242_io_reset = reset; // @[RegFile.scala 78:19:@41029.4]
  assign regs_242_io_enable = 1'h1; // @[RegFile.scala 74:20:@41023.4]
  assign regs_243_clock = clock; // @[:@41032.4]
  assign regs_243_reset = io_reset; // @[:@41033.4 RegFile.scala 76:16:@41040.4]
  assign regs_243_io_in = 64'h0; // @[RegFile.scala 75:16:@41039.4]
  assign regs_243_io_reset = reset; // @[RegFile.scala 78:19:@41043.4]
  assign regs_243_io_enable = 1'h1; // @[RegFile.scala 74:20:@41037.4]
  assign regs_244_clock = clock; // @[:@41046.4]
  assign regs_244_reset = io_reset; // @[:@41047.4 RegFile.scala 76:16:@41054.4]
  assign regs_244_io_in = 64'h0; // @[RegFile.scala 75:16:@41053.4]
  assign regs_244_io_reset = reset; // @[RegFile.scala 78:19:@41057.4]
  assign regs_244_io_enable = 1'h1; // @[RegFile.scala 74:20:@41051.4]
  assign regs_245_clock = clock; // @[:@41060.4]
  assign regs_245_reset = io_reset; // @[:@41061.4 RegFile.scala 76:16:@41068.4]
  assign regs_245_io_in = 64'h0; // @[RegFile.scala 75:16:@41067.4]
  assign regs_245_io_reset = reset; // @[RegFile.scala 78:19:@41071.4]
  assign regs_245_io_enable = 1'h1; // @[RegFile.scala 74:20:@41065.4]
  assign regs_246_clock = clock; // @[:@41074.4]
  assign regs_246_reset = io_reset; // @[:@41075.4 RegFile.scala 76:16:@41082.4]
  assign regs_246_io_in = 64'h0; // @[RegFile.scala 75:16:@41081.4]
  assign regs_246_io_reset = reset; // @[RegFile.scala 78:19:@41085.4]
  assign regs_246_io_enable = 1'h1; // @[RegFile.scala 74:20:@41079.4]
  assign regs_247_clock = clock; // @[:@41088.4]
  assign regs_247_reset = io_reset; // @[:@41089.4 RegFile.scala 76:16:@41096.4]
  assign regs_247_io_in = 64'h0; // @[RegFile.scala 75:16:@41095.4]
  assign regs_247_io_reset = reset; // @[RegFile.scala 78:19:@41099.4]
  assign regs_247_io_enable = 1'h1; // @[RegFile.scala 74:20:@41093.4]
  assign regs_248_clock = clock; // @[:@41102.4]
  assign regs_248_reset = io_reset; // @[:@41103.4 RegFile.scala 76:16:@41110.4]
  assign regs_248_io_in = 64'h0; // @[RegFile.scala 75:16:@41109.4]
  assign regs_248_io_reset = reset; // @[RegFile.scala 78:19:@41113.4]
  assign regs_248_io_enable = 1'h1; // @[RegFile.scala 74:20:@41107.4]
  assign regs_249_clock = clock; // @[:@41116.4]
  assign regs_249_reset = io_reset; // @[:@41117.4 RegFile.scala 76:16:@41124.4]
  assign regs_249_io_in = 64'h0; // @[RegFile.scala 75:16:@41123.4]
  assign regs_249_io_reset = reset; // @[RegFile.scala 78:19:@41127.4]
  assign regs_249_io_enable = 1'h1; // @[RegFile.scala 74:20:@41121.4]
  assign regs_250_clock = clock; // @[:@41130.4]
  assign regs_250_reset = io_reset; // @[:@41131.4 RegFile.scala 76:16:@41138.4]
  assign regs_250_io_in = 64'h0; // @[RegFile.scala 75:16:@41137.4]
  assign regs_250_io_reset = reset; // @[RegFile.scala 78:19:@41141.4]
  assign regs_250_io_enable = 1'h1; // @[RegFile.scala 74:20:@41135.4]
  assign regs_251_clock = clock; // @[:@41144.4]
  assign regs_251_reset = io_reset; // @[:@41145.4 RegFile.scala 76:16:@41152.4]
  assign regs_251_io_in = 64'h0; // @[RegFile.scala 75:16:@41151.4]
  assign regs_251_io_reset = reset; // @[RegFile.scala 78:19:@41155.4]
  assign regs_251_io_enable = 1'h1; // @[RegFile.scala 74:20:@41149.4]
  assign regs_252_clock = clock; // @[:@41158.4]
  assign regs_252_reset = io_reset; // @[:@41159.4 RegFile.scala 76:16:@41166.4]
  assign regs_252_io_in = 64'h0; // @[RegFile.scala 75:16:@41165.4]
  assign regs_252_io_reset = reset; // @[RegFile.scala 78:19:@41169.4]
  assign regs_252_io_enable = 1'h1; // @[RegFile.scala 74:20:@41163.4]
  assign regs_253_clock = clock; // @[:@41172.4]
  assign regs_253_reset = io_reset; // @[:@41173.4 RegFile.scala 76:16:@41180.4]
  assign regs_253_io_in = 64'h0; // @[RegFile.scala 75:16:@41179.4]
  assign regs_253_io_reset = reset; // @[RegFile.scala 78:19:@41183.4]
  assign regs_253_io_enable = 1'h1; // @[RegFile.scala 74:20:@41177.4]
  assign regs_254_clock = clock; // @[:@41186.4]
  assign regs_254_reset = io_reset; // @[:@41187.4 RegFile.scala 76:16:@41194.4]
  assign regs_254_io_in = 64'h0; // @[RegFile.scala 75:16:@41193.4]
  assign regs_254_io_reset = reset; // @[RegFile.scala 78:19:@41197.4]
  assign regs_254_io_enable = 1'h1; // @[RegFile.scala 74:20:@41191.4]
  assign regs_255_clock = clock; // @[:@41200.4]
  assign regs_255_reset = io_reset; // @[:@41201.4 RegFile.scala 76:16:@41208.4]
  assign regs_255_io_in = 64'h0; // @[RegFile.scala 75:16:@41207.4]
  assign regs_255_io_reset = reset; // @[RegFile.scala 78:19:@41211.4]
  assign regs_255_io_enable = 1'h1; // @[RegFile.scala 74:20:@41205.4]
  assign regs_256_clock = clock; // @[:@41214.4]
  assign regs_256_reset = io_reset; // @[:@41215.4 RegFile.scala 76:16:@41222.4]
  assign regs_256_io_in = 64'h0; // @[RegFile.scala 75:16:@41221.4]
  assign regs_256_io_reset = reset; // @[RegFile.scala 78:19:@41225.4]
  assign regs_256_io_enable = 1'h1; // @[RegFile.scala 74:20:@41219.4]
  assign regs_257_clock = clock; // @[:@41228.4]
  assign regs_257_reset = io_reset; // @[:@41229.4 RegFile.scala 76:16:@41236.4]
  assign regs_257_io_in = 64'h0; // @[RegFile.scala 75:16:@41235.4]
  assign regs_257_io_reset = reset; // @[RegFile.scala 78:19:@41239.4]
  assign regs_257_io_enable = 1'h1; // @[RegFile.scala 74:20:@41233.4]
  assign regs_258_clock = clock; // @[:@41242.4]
  assign regs_258_reset = io_reset; // @[:@41243.4 RegFile.scala 76:16:@41250.4]
  assign regs_258_io_in = 64'h0; // @[RegFile.scala 75:16:@41249.4]
  assign regs_258_io_reset = reset; // @[RegFile.scala 78:19:@41253.4]
  assign regs_258_io_enable = 1'h1; // @[RegFile.scala 74:20:@41247.4]
  assign regs_259_clock = clock; // @[:@41256.4]
  assign regs_259_reset = io_reset; // @[:@41257.4 RegFile.scala 76:16:@41264.4]
  assign regs_259_io_in = 64'h0; // @[RegFile.scala 75:16:@41263.4]
  assign regs_259_io_reset = reset; // @[RegFile.scala 78:19:@41267.4]
  assign regs_259_io_enable = 1'h1; // @[RegFile.scala 74:20:@41261.4]
  assign regs_260_clock = clock; // @[:@41270.4]
  assign regs_260_reset = io_reset; // @[:@41271.4 RegFile.scala 76:16:@41278.4]
  assign regs_260_io_in = 64'h0; // @[RegFile.scala 75:16:@41277.4]
  assign regs_260_io_reset = reset; // @[RegFile.scala 78:19:@41281.4]
  assign regs_260_io_enable = 1'h1; // @[RegFile.scala 74:20:@41275.4]
  assign regs_261_clock = clock; // @[:@41284.4]
  assign regs_261_reset = io_reset; // @[:@41285.4 RegFile.scala 76:16:@41292.4]
  assign regs_261_io_in = 64'h0; // @[RegFile.scala 75:16:@41291.4]
  assign regs_261_io_reset = reset; // @[RegFile.scala 78:19:@41295.4]
  assign regs_261_io_enable = 1'h1; // @[RegFile.scala 74:20:@41289.4]
  assign regs_262_clock = clock; // @[:@41298.4]
  assign regs_262_reset = io_reset; // @[:@41299.4 RegFile.scala 76:16:@41306.4]
  assign regs_262_io_in = 64'h0; // @[RegFile.scala 75:16:@41305.4]
  assign regs_262_io_reset = reset; // @[RegFile.scala 78:19:@41309.4]
  assign regs_262_io_enable = 1'h1; // @[RegFile.scala 74:20:@41303.4]
  assign regs_263_clock = clock; // @[:@41312.4]
  assign regs_263_reset = io_reset; // @[:@41313.4 RegFile.scala 76:16:@41320.4]
  assign regs_263_io_in = 64'h0; // @[RegFile.scala 75:16:@41319.4]
  assign regs_263_io_reset = reset; // @[RegFile.scala 78:19:@41323.4]
  assign regs_263_io_enable = 1'h1; // @[RegFile.scala 74:20:@41317.4]
  assign regs_264_clock = clock; // @[:@41326.4]
  assign regs_264_reset = io_reset; // @[:@41327.4 RegFile.scala 76:16:@41334.4]
  assign regs_264_io_in = 64'h0; // @[RegFile.scala 75:16:@41333.4]
  assign regs_264_io_reset = reset; // @[RegFile.scala 78:19:@41337.4]
  assign regs_264_io_enable = 1'h1; // @[RegFile.scala 74:20:@41331.4]
  assign regs_265_clock = clock; // @[:@41340.4]
  assign regs_265_reset = io_reset; // @[:@41341.4 RegFile.scala 76:16:@41348.4]
  assign regs_265_io_in = 64'h0; // @[RegFile.scala 75:16:@41347.4]
  assign regs_265_io_reset = reset; // @[RegFile.scala 78:19:@41351.4]
  assign regs_265_io_enable = 1'h1; // @[RegFile.scala 74:20:@41345.4]
  assign regs_266_clock = clock; // @[:@41354.4]
  assign regs_266_reset = io_reset; // @[:@41355.4 RegFile.scala 76:16:@41362.4]
  assign regs_266_io_in = 64'h0; // @[RegFile.scala 75:16:@41361.4]
  assign regs_266_io_reset = reset; // @[RegFile.scala 78:19:@41365.4]
  assign regs_266_io_enable = 1'h1; // @[RegFile.scala 74:20:@41359.4]
  assign regs_267_clock = clock; // @[:@41368.4]
  assign regs_267_reset = io_reset; // @[:@41369.4 RegFile.scala 76:16:@41376.4]
  assign regs_267_io_in = 64'h0; // @[RegFile.scala 75:16:@41375.4]
  assign regs_267_io_reset = reset; // @[RegFile.scala 78:19:@41379.4]
  assign regs_267_io_enable = 1'h1; // @[RegFile.scala 74:20:@41373.4]
  assign regs_268_clock = clock; // @[:@41382.4]
  assign regs_268_reset = io_reset; // @[:@41383.4 RegFile.scala 76:16:@41390.4]
  assign regs_268_io_in = 64'h0; // @[RegFile.scala 75:16:@41389.4]
  assign regs_268_io_reset = reset; // @[RegFile.scala 78:19:@41393.4]
  assign regs_268_io_enable = 1'h1; // @[RegFile.scala 74:20:@41387.4]
  assign regs_269_clock = clock; // @[:@41396.4]
  assign regs_269_reset = io_reset; // @[:@41397.4 RegFile.scala 76:16:@41404.4]
  assign regs_269_io_in = 64'h0; // @[RegFile.scala 75:16:@41403.4]
  assign regs_269_io_reset = reset; // @[RegFile.scala 78:19:@41407.4]
  assign regs_269_io_enable = 1'h1; // @[RegFile.scala 74:20:@41401.4]
  assign regs_270_clock = clock; // @[:@41410.4]
  assign regs_270_reset = io_reset; // @[:@41411.4 RegFile.scala 76:16:@41418.4]
  assign regs_270_io_in = 64'h0; // @[RegFile.scala 75:16:@41417.4]
  assign regs_270_io_reset = reset; // @[RegFile.scala 78:19:@41421.4]
  assign regs_270_io_enable = 1'h1; // @[RegFile.scala 74:20:@41415.4]
  assign regs_271_clock = clock; // @[:@41424.4]
  assign regs_271_reset = io_reset; // @[:@41425.4 RegFile.scala 76:16:@41432.4]
  assign regs_271_io_in = 64'h0; // @[RegFile.scala 75:16:@41431.4]
  assign regs_271_io_reset = reset; // @[RegFile.scala 78:19:@41435.4]
  assign regs_271_io_enable = 1'h1; // @[RegFile.scala 74:20:@41429.4]
  assign regs_272_clock = clock; // @[:@41438.4]
  assign regs_272_reset = io_reset; // @[:@41439.4 RegFile.scala 76:16:@41446.4]
  assign regs_272_io_in = 64'h0; // @[RegFile.scala 75:16:@41445.4]
  assign regs_272_io_reset = reset; // @[RegFile.scala 78:19:@41449.4]
  assign regs_272_io_enable = 1'h1; // @[RegFile.scala 74:20:@41443.4]
  assign regs_273_clock = clock; // @[:@41452.4]
  assign regs_273_reset = io_reset; // @[:@41453.4 RegFile.scala 76:16:@41460.4]
  assign regs_273_io_in = 64'h0; // @[RegFile.scala 75:16:@41459.4]
  assign regs_273_io_reset = reset; // @[RegFile.scala 78:19:@41463.4]
  assign regs_273_io_enable = 1'h1; // @[RegFile.scala 74:20:@41457.4]
  assign regs_274_clock = clock; // @[:@41466.4]
  assign regs_274_reset = io_reset; // @[:@41467.4 RegFile.scala 76:16:@41474.4]
  assign regs_274_io_in = 64'h0; // @[RegFile.scala 75:16:@41473.4]
  assign regs_274_io_reset = reset; // @[RegFile.scala 78:19:@41477.4]
  assign regs_274_io_enable = 1'h1; // @[RegFile.scala 74:20:@41471.4]
  assign regs_275_clock = clock; // @[:@41480.4]
  assign regs_275_reset = io_reset; // @[:@41481.4 RegFile.scala 76:16:@41488.4]
  assign regs_275_io_in = 64'h0; // @[RegFile.scala 75:16:@41487.4]
  assign regs_275_io_reset = reset; // @[RegFile.scala 78:19:@41491.4]
  assign regs_275_io_enable = 1'h1; // @[RegFile.scala 74:20:@41485.4]
  assign regs_276_clock = clock; // @[:@41494.4]
  assign regs_276_reset = io_reset; // @[:@41495.4 RegFile.scala 76:16:@41502.4]
  assign regs_276_io_in = 64'h0; // @[RegFile.scala 75:16:@41501.4]
  assign regs_276_io_reset = reset; // @[RegFile.scala 78:19:@41505.4]
  assign regs_276_io_enable = 1'h1; // @[RegFile.scala 74:20:@41499.4]
  assign regs_277_clock = clock; // @[:@41508.4]
  assign regs_277_reset = io_reset; // @[:@41509.4 RegFile.scala 76:16:@41516.4]
  assign regs_277_io_in = 64'h0; // @[RegFile.scala 75:16:@41515.4]
  assign regs_277_io_reset = reset; // @[RegFile.scala 78:19:@41519.4]
  assign regs_277_io_enable = 1'h1; // @[RegFile.scala 74:20:@41513.4]
  assign regs_278_clock = clock; // @[:@41522.4]
  assign regs_278_reset = io_reset; // @[:@41523.4 RegFile.scala 76:16:@41530.4]
  assign regs_278_io_in = 64'h0; // @[RegFile.scala 75:16:@41529.4]
  assign regs_278_io_reset = reset; // @[RegFile.scala 78:19:@41533.4]
  assign regs_278_io_enable = 1'h1; // @[RegFile.scala 74:20:@41527.4]
  assign regs_279_clock = clock; // @[:@41536.4]
  assign regs_279_reset = io_reset; // @[:@41537.4 RegFile.scala 76:16:@41544.4]
  assign regs_279_io_in = 64'h0; // @[RegFile.scala 75:16:@41543.4]
  assign regs_279_io_reset = reset; // @[RegFile.scala 78:19:@41547.4]
  assign regs_279_io_enable = 1'h1; // @[RegFile.scala 74:20:@41541.4]
  assign regs_280_clock = clock; // @[:@41550.4]
  assign regs_280_reset = io_reset; // @[:@41551.4 RegFile.scala 76:16:@41558.4]
  assign regs_280_io_in = 64'h0; // @[RegFile.scala 75:16:@41557.4]
  assign regs_280_io_reset = reset; // @[RegFile.scala 78:19:@41561.4]
  assign regs_280_io_enable = 1'h1; // @[RegFile.scala 74:20:@41555.4]
  assign regs_281_clock = clock; // @[:@41564.4]
  assign regs_281_reset = io_reset; // @[:@41565.4 RegFile.scala 76:16:@41572.4]
  assign regs_281_io_in = 64'h0; // @[RegFile.scala 75:16:@41571.4]
  assign regs_281_io_reset = reset; // @[RegFile.scala 78:19:@41575.4]
  assign regs_281_io_enable = 1'h1; // @[RegFile.scala 74:20:@41569.4]
  assign regs_282_clock = clock; // @[:@41578.4]
  assign regs_282_reset = io_reset; // @[:@41579.4 RegFile.scala 76:16:@41586.4]
  assign regs_282_io_in = 64'h0; // @[RegFile.scala 75:16:@41585.4]
  assign regs_282_io_reset = reset; // @[RegFile.scala 78:19:@41589.4]
  assign regs_282_io_enable = 1'h1; // @[RegFile.scala 74:20:@41583.4]
  assign regs_283_clock = clock; // @[:@41592.4]
  assign regs_283_reset = io_reset; // @[:@41593.4 RegFile.scala 76:16:@41600.4]
  assign regs_283_io_in = 64'h0; // @[RegFile.scala 75:16:@41599.4]
  assign regs_283_io_reset = reset; // @[RegFile.scala 78:19:@41603.4]
  assign regs_283_io_enable = 1'h1; // @[RegFile.scala 74:20:@41597.4]
  assign regs_284_clock = clock; // @[:@41606.4]
  assign regs_284_reset = io_reset; // @[:@41607.4 RegFile.scala 76:16:@41614.4]
  assign regs_284_io_in = 64'h0; // @[RegFile.scala 75:16:@41613.4]
  assign regs_284_io_reset = reset; // @[RegFile.scala 78:19:@41617.4]
  assign regs_284_io_enable = 1'h1; // @[RegFile.scala 74:20:@41611.4]
  assign regs_285_clock = clock; // @[:@41620.4]
  assign regs_285_reset = io_reset; // @[:@41621.4 RegFile.scala 76:16:@41628.4]
  assign regs_285_io_in = 64'h0; // @[RegFile.scala 75:16:@41627.4]
  assign regs_285_io_reset = reset; // @[RegFile.scala 78:19:@41631.4]
  assign regs_285_io_enable = 1'h1; // @[RegFile.scala 74:20:@41625.4]
  assign regs_286_clock = clock; // @[:@41634.4]
  assign regs_286_reset = io_reset; // @[:@41635.4 RegFile.scala 76:16:@41642.4]
  assign regs_286_io_in = 64'h0; // @[RegFile.scala 75:16:@41641.4]
  assign regs_286_io_reset = reset; // @[RegFile.scala 78:19:@41645.4]
  assign regs_286_io_enable = 1'h1; // @[RegFile.scala 74:20:@41639.4]
  assign regs_287_clock = clock; // @[:@41648.4]
  assign regs_287_reset = io_reset; // @[:@41649.4 RegFile.scala 76:16:@41656.4]
  assign regs_287_io_in = 64'h0; // @[RegFile.scala 75:16:@41655.4]
  assign regs_287_io_reset = reset; // @[RegFile.scala 78:19:@41659.4]
  assign regs_287_io_enable = 1'h1; // @[RegFile.scala 74:20:@41653.4]
  assign regs_288_clock = clock; // @[:@41662.4]
  assign regs_288_reset = io_reset; // @[:@41663.4 RegFile.scala 76:16:@41670.4]
  assign regs_288_io_in = 64'h0; // @[RegFile.scala 75:16:@41669.4]
  assign regs_288_io_reset = reset; // @[RegFile.scala 78:19:@41673.4]
  assign regs_288_io_enable = 1'h1; // @[RegFile.scala 74:20:@41667.4]
  assign regs_289_clock = clock; // @[:@41676.4]
  assign regs_289_reset = io_reset; // @[:@41677.4 RegFile.scala 76:16:@41684.4]
  assign regs_289_io_in = 64'h0; // @[RegFile.scala 75:16:@41683.4]
  assign regs_289_io_reset = reset; // @[RegFile.scala 78:19:@41687.4]
  assign regs_289_io_enable = 1'h1; // @[RegFile.scala 74:20:@41681.4]
  assign regs_290_clock = clock; // @[:@41690.4]
  assign regs_290_reset = io_reset; // @[:@41691.4 RegFile.scala 76:16:@41698.4]
  assign regs_290_io_in = 64'h0; // @[RegFile.scala 75:16:@41697.4]
  assign regs_290_io_reset = reset; // @[RegFile.scala 78:19:@41701.4]
  assign regs_290_io_enable = 1'h1; // @[RegFile.scala 74:20:@41695.4]
  assign regs_291_clock = clock; // @[:@41704.4]
  assign regs_291_reset = io_reset; // @[:@41705.4 RegFile.scala 76:16:@41712.4]
  assign regs_291_io_in = 64'h0; // @[RegFile.scala 75:16:@41711.4]
  assign regs_291_io_reset = reset; // @[RegFile.scala 78:19:@41715.4]
  assign regs_291_io_enable = 1'h1; // @[RegFile.scala 74:20:@41709.4]
  assign regs_292_clock = clock; // @[:@41718.4]
  assign regs_292_reset = io_reset; // @[:@41719.4 RegFile.scala 76:16:@41726.4]
  assign regs_292_io_in = 64'h0; // @[RegFile.scala 75:16:@41725.4]
  assign regs_292_io_reset = reset; // @[RegFile.scala 78:19:@41729.4]
  assign regs_292_io_enable = 1'h1; // @[RegFile.scala 74:20:@41723.4]
  assign regs_293_clock = clock; // @[:@41732.4]
  assign regs_293_reset = io_reset; // @[:@41733.4 RegFile.scala 76:16:@41740.4]
  assign regs_293_io_in = 64'h0; // @[RegFile.scala 75:16:@41739.4]
  assign regs_293_io_reset = reset; // @[RegFile.scala 78:19:@41743.4]
  assign regs_293_io_enable = 1'h1; // @[RegFile.scala 74:20:@41737.4]
  assign regs_294_clock = clock; // @[:@41746.4]
  assign regs_294_reset = io_reset; // @[:@41747.4 RegFile.scala 76:16:@41754.4]
  assign regs_294_io_in = 64'h0; // @[RegFile.scala 75:16:@41753.4]
  assign regs_294_io_reset = reset; // @[RegFile.scala 78:19:@41757.4]
  assign regs_294_io_enable = 1'h1; // @[RegFile.scala 74:20:@41751.4]
  assign regs_295_clock = clock; // @[:@41760.4]
  assign regs_295_reset = io_reset; // @[:@41761.4 RegFile.scala 76:16:@41768.4]
  assign regs_295_io_in = 64'h0; // @[RegFile.scala 75:16:@41767.4]
  assign regs_295_io_reset = reset; // @[RegFile.scala 78:19:@41771.4]
  assign regs_295_io_enable = 1'h1; // @[RegFile.scala 74:20:@41765.4]
  assign regs_296_clock = clock; // @[:@41774.4]
  assign regs_296_reset = io_reset; // @[:@41775.4 RegFile.scala 76:16:@41782.4]
  assign regs_296_io_in = 64'h0; // @[RegFile.scala 75:16:@41781.4]
  assign regs_296_io_reset = reset; // @[RegFile.scala 78:19:@41785.4]
  assign regs_296_io_enable = 1'h1; // @[RegFile.scala 74:20:@41779.4]
  assign regs_297_clock = clock; // @[:@41788.4]
  assign regs_297_reset = io_reset; // @[:@41789.4 RegFile.scala 76:16:@41796.4]
  assign regs_297_io_in = 64'h0; // @[RegFile.scala 75:16:@41795.4]
  assign regs_297_io_reset = reset; // @[RegFile.scala 78:19:@41799.4]
  assign regs_297_io_enable = 1'h1; // @[RegFile.scala 74:20:@41793.4]
  assign regs_298_clock = clock; // @[:@41802.4]
  assign regs_298_reset = io_reset; // @[:@41803.4 RegFile.scala 76:16:@41810.4]
  assign regs_298_io_in = 64'h0; // @[RegFile.scala 75:16:@41809.4]
  assign regs_298_io_reset = reset; // @[RegFile.scala 78:19:@41813.4]
  assign regs_298_io_enable = 1'h1; // @[RegFile.scala 74:20:@41807.4]
  assign regs_299_clock = clock; // @[:@41816.4]
  assign regs_299_reset = io_reset; // @[:@41817.4 RegFile.scala 76:16:@41824.4]
  assign regs_299_io_in = 64'h0; // @[RegFile.scala 75:16:@41823.4]
  assign regs_299_io_reset = reset; // @[RegFile.scala 78:19:@41827.4]
  assign regs_299_io_enable = 1'h1; // @[RegFile.scala 74:20:@41821.4]
  assign regs_300_clock = clock; // @[:@41830.4]
  assign regs_300_reset = io_reset; // @[:@41831.4 RegFile.scala 76:16:@41838.4]
  assign regs_300_io_in = 64'h0; // @[RegFile.scala 75:16:@41837.4]
  assign regs_300_io_reset = reset; // @[RegFile.scala 78:19:@41841.4]
  assign regs_300_io_enable = 1'h1; // @[RegFile.scala 74:20:@41835.4]
  assign regs_301_clock = clock; // @[:@41844.4]
  assign regs_301_reset = io_reset; // @[:@41845.4 RegFile.scala 76:16:@41852.4]
  assign regs_301_io_in = 64'h0; // @[RegFile.scala 75:16:@41851.4]
  assign regs_301_io_reset = reset; // @[RegFile.scala 78:19:@41855.4]
  assign regs_301_io_enable = 1'h1; // @[RegFile.scala 74:20:@41849.4]
  assign regs_302_clock = clock; // @[:@41858.4]
  assign regs_302_reset = io_reset; // @[:@41859.4 RegFile.scala 76:16:@41866.4]
  assign regs_302_io_in = 64'h0; // @[RegFile.scala 75:16:@41865.4]
  assign regs_302_io_reset = reset; // @[RegFile.scala 78:19:@41869.4]
  assign regs_302_io_enable = 1'h1; // @[RegFile.scala 74:20:@41863.4]
  assign regs_303_clock = clock; // @[:@41872.4]
  assign regs_303_reset = io_reset; // @[:@41873.4 RegFile.scala 76:16:@41880.4]
  assign regs_303_io_in = 64'h0; // @[RegFile.scala 75:16:@41879.4]
  assign regs_303_io_reset = reset; // @[RegFile.scala 78:19:@41883.4]
  assign regs_303_io_enable = 1'h1; // @[RegFile.scala 74:20:@41877.4]
  assign regs_304_clock = clock; // @[:@41886.4]
  assign regs_304_reset = io_reset; // @[:@41887.4 RegFile.scala 76:16:@41894.4]
  assign regs_304_io_in = 64'h0; // @[RegFile.scala 75:16:@41893.4]
  assign regs_304_io_reset = reset; // @[RegFile.scala 78:19:@41897.4]
  assign regs_304_io_enable = 1'h1; // @[RegFile.scala 74:20:@41891.4]
  assign regs_305_clock = clock; // @[:@41900.4]
  assign regs_305_reset = io_reset; // @[:@41901.4 RegFile.scala 76:16:@41908.4]
  assign regs_305_io_in = 64'h0; // @[RegFile.scala 75:16:@41907.4]
  assign regs_305_io_reset = reset; // @[RegFile.scala 78:19:@41911.4]
  assign regs_305_io_enable = 1'h1; // @[RegFile.scala 74:20:@41905.4]
  assign regs_306_clock = clock; // @[:@41914.4]
  assign regs_306_reset = io_reset; // @[:@41915.4 RegFile.scala 76:16:@41922.4]
  assign regs_306_io_in = 64'h0; // @[RegFile.scala 75:16:@41921.4]
  assign regs_306_io_reset = reset; // @[RegFile.scala 78:19:@41925.4]
  assign regs_306_io_enable = 1'h1; // @[RegFile.scala 74:20:@41919.4]
  assign regs_307_clock = clock; // @[:@41928.4]
  assign regs_307_reset = io_reset; // @[:@41929.4 RegFile.scala 76:16:@41936.4]
  assign regs_307_io_in = 64'h0; // @[RegFile.scala 75:16:@41935.4]
  assign regs_307_io_reset = reset; // @[RegFile.scala 78:19:@41939.4]
  assign regs_307_io_enable = 1'h1; // @[RegFile.scala 74:20:@41933.4]
  assign regs_308_clock = clock; // @[:@41942.4]
  assign regs_308_reset = io_reset; // @[:@41943.4 RegFile.scala 76:16:@41950.4]
  assign regs_308_io_in = 64'h0; // @[RegFile.scala 75:16:@41949.4]
  assign regs_308_io_reset = reset; // @[RegFile.scala 78:19:@41953.4]
  assign regs_308_io_enable = 1'h1; // @[RegFile.scala 74:20:@41947.4]
  assign regs_309_clock = clock; // @[:@41956.4]
  assign regs_309_reset = io_reset; // @[:@41957.4 RegFile.scala 76:16:@41964.4]
  assign regs_309_io_in = 64'h0; // @[RegFile.scala 75:16:@41963.4]
  assign regs_309_io_reset = reset; // @[RegFile.scala 78:19:@41967.4]
  assign regs_309_io_enable = 1'h1; // @[RegFile.scala 74:20:@41961.4]
  assign regs_310_clock = clock; // @[:@41970.4]
  assign regs_310_reset = io_reset; // @[:@41971.4 RegFile.scala 76:16:@41978.4]
  assign regs_310_io_in = 64'h0; // @[RegFile.scala 75:16:@41977.4]
  assign regs_310_io_reset = reset; // @[RegFile.scala 78:19:@41981.4]
  assign regs_310_io_enable = 1'h1; // @[RegFile.scala 74:20:@41975.4]
  assign regs_311_clock = clock; // @[:@41984.4]
  assign regs_311_reset = io_reset; // @[:@41985.4 RegFile.scala 76:16:@41992.4]
  assign regs_311_io_in = 64'h0; // @[RegFile.scala 75:16:@41991.4]
  assign regs_311_io_reset = reset; // @[RegFile.scala 78:19:@41995.4]
  assign regs_311_io_enable = 1'h1; // @[RegFile.scala 74:20:@41989.4]
  assign regs_312_clock = clock; // @[:@41998.4]
  assign regs_312_reset = io_reset; // @[:@41999.4 RegFile.scala 76:16:@42006.4]
  assign regs_312_io_in = 64'h0; // @[RegFile.scala 75:16:@42005.4]
  assign regs_312_io_reset = reset; // @[RegFile.scala 78:19:@42009.4]
  assign regs_312_io_enable = 1'h1; // @[RegFile.scala 74:20:@42003.4]
  assign regs_313_clock = clock; // @[:@42012.4]
  assign regs_313_reset = io_reset; // @[:@42013.4 RegFile.scala 76:16:@42020.4]
  assign regs_313_io_in = 64'h0; // @[RegFile.scala 75:16:@42019.4]
  assign regs_313_io_reset = reset; // @[RegFile.scala 78:19:@42023.4]
  assign regs_313_io_enable = 1'h1; // @[RegFile.scala 74:20:@42017.4]
  assign regs_314_clock = clock; // @[:@42026.4]
  assign regs_314_reset = io_reset; // @[:@42027.4 RegFile.scala 76:16:@42034.4]
  assign regs_314_io_in = 64'h0; // @[RegFile.scala 75:16:@42033.4]
  assign regs_314_io_reset = reset; // @[RegFile.scala 78:19:@42037.4]
  assign regs_314_io_enable = 1'h1; // @[RegFile.scala 74:20:@42031.4]
  assign regs_315_clock = clock; // @[:@42040.4]
  assign regs_315_reset = io_reset; // @[:@42041.4 RegFile.scala 76:16:@42048.4]
  assign regs_315_io_in = 64'h0; // @[RegFile.scala 75:16:@42047.4]
  assign regs_315_io_reset = reset; // @[RegFile.scala 78:19:@42051.4]
  assign regs_315_io_enable = 1'h1; // @[RegFile.scala 74:20:@42045.4]
  assign regs_316_clock = clock; // @[:@42054.4]
  assign regs_316_reset = io_reset; // @[:@42055.4 RegFile.scala 76:16:@42062.4]
  assign regs_316_io_in = 64'h0; // @[RegFile.scala 75:16:@42061.4]
  assign regs_316_io_reset = reset; // @[RegFile.scala 78:19:@42065.4]
  assign regs_316_io_enable = 1'h1; // @[RegFile.scala 74:20:@42059.4]
  assign regs_317_clock = clock; // @[:@42068.4]
  assign regs_317_reset = io_reset; // @[:@42069.4 RegFile.scala 76:16:@42076.4]
  assign regs_317_io_in = 64'h0; // @[RegFile.scala 75:16:@42075.4]
  assign regs_317_io_reset = reset; // @[RegFile.scala 78:19:@42079.4]
  assign regs_317_io_enable = 1'h1; // @[RegFile.scala 74:20:@42073.4]
  assign regs_318_clock = clock; // @[:@42082.4]
  assign regs_318_reset = io_reset; // @[:@42083.4 RegFile.scala 76:16:@42090.4]
  assign regs_318_io_in = 64'h0; // @[RegFile.scala 75:16:@42089.4]
  assign regs_318_io_reset = reset; // @[RegFile.scala 78:19:@42093.4]
  assign regs_318_io_enable = 1'h1; // @[RegFile.scala 74:20:@42087.4]
  assign regs_319_clock = clock; // @[:@42096.4]
  assign regs_319_reset = io_reset; // @[:@42097.4 RegFile.scala 76:16:@42104.4]
  assign regs_319_io_in = 64'h0; // @[RegFile.scala 75:16:@42103.4]
  assign regs_319_io_reset = reset; // @[RegFile.scala 78:19:@42107.4]
  assign regs_319_io_enable = 1'h1; // @[RegFile.scala 74:20:@42101.4]
  assign regs_320_clock = clock; // @[:@42110.4]
  assign regs_320_reset = io_reset; // @[:@42111.4 RegFile.scala 76:16:@42118.4]
  assign regs_320_io_in = 64'h0; // @[RegFile.scala 75:16:@42117.4]
  assign regs_320_io_reset = reset; // @[RegFile.scala 78:19:@42121.4]
  assign regs_320_io_enable = 1'h1; // @[RegFile.scala 74:20:@42115.4]
  assign regs_321_clock = clock; // @[:@42124.4]
  assign regs_321_reset = io_reset; // @[:@42125.4 RegFile.scala 76:16:@42132.4]
  assign regs_321_io_in = 64'h0; // @[RegFile.scala 75:16:@42131.4]
  assign regs_321_io_reset = reset; // @[RegFile.scala 78:19:@42135.4]
  assign regs_321_io_enable = 1'h1; // @[RegFile.scala 74:20:@42129.4]
  assign regs_322_clock = clock; // @[:@42138.4]
  assign regs_322_reset = io_reset; // @[:@42139.4 RegFile.scala 76:16:@42146.4]
  assign regs_322_io_in = 64'h0; // @[RegFile.scala 75:16:@42145.4]
  assign regs_322_io_reset = reset; // @[RegFile.scala 78:19:@42149.4]
  assign regs_322_io_enable = 1'h1; // @[RegFile.scala 74:20:@42143.4]
  assign regs_323_clock = clock; // @[:@42152.4]
  assign regs_323_reset = io_reset; // @[:@42153.4 RegFile.scala 76:16:@42160.4]
  assign regs_323_io_in = 64'h0; // @[RegFile.scala 75:16:@42159.4]
  assign regs_323_io_reset = reset; // @[RegFile.scala 78:19:@42163.4]
  assign regs_323_io_enable = 1'h1; // @[RegFile.scala 74:20:@42157.4]
  assign regs_324_clock = clock; // @[:@42166.4]
  assign regs_324_reset = io_reset; // @[:@42167.4 RegFile.scala 76:16:@42174.4]
  assign regs_324_io_in = 64'h0; // @[RegFile.scala 75:16:@42173.4]
  assign regs_324_io_reset = reset; // @[RegFile.scala 78:19:@42177.4]
  assign regs_324_io_enable = 1'h1; // @[RegFile.scala 74:20:@42171.4]
  assign regs_325_clock = clock; // @[:@42180.4]
  assign regs_325_reset = io_reset; // @[:@42181.4 RegFile.scala 76:16:@42188.4]
  assign regs_325_io_in = 64'h0; // @[RegFile.scala 75:16:@42187.4]
  assign regs_325_io_reset = reset; // @[RegFile.scala 78:19:@42191.4]
  assign regs_325_io_enable = 1'h1; // @[RegFile.scala 74:20:@42185.4]
  assign regs_326_clock = clock; // @[:@42194.4]
  assign regs_326_reset = io_reset; // @[:@42195.4 RegFile.scala 76:16:@42202.4]
  assign regs_326_io_in = 64'h0; // @[RegFile.scala 75:16:@42201.4]
  assign regs_326_io_reset = reset; // @[RegFile.scala 78:19:@42205.4]
  assign regs_326_io_enable = 1'h1; // @[RegFile.scala 74:20:@42199.4]
  assign regs_327_clock = clock; // @[:@42208.4]
  assign regs_327_reset = io_reset; // @[:@42209.4 RegFile.scala 76:16:@42216.4]
  assign regs_327_io_in = 64'h0; // @[RegFile.scala 75:16:@42215.4]
  assign regs_327_io_reset = reset; // @[RegFile.scala 78:19:@42219.4]
  assign regs_327_io_enable = 1'h1; // @[RegFile.scala 74:20:@42213.4]
  assign regs_328_clock = clock; // @[:@42222.4]
  assign regs_328_reset = io_reset; // @[:@42223.4 RegFile.scala 76:16:@42230.4]
  assign regs_328_io_in = 64'h0; // @[RegFile.scala 75:16:@42229.4]
  assign regs_328_io_reset = reset; // @[RegFile.scala 78:19:@42233.4]
  assign regs_328_io_enable = 1'h1; // @[RegFile.scala 74:20:@42227.4]
  assign regs_329_clock = clock; // @[:@42236.4]
  assign regs_329_reset = io_reset; // @[:@42237.4 RegFile.scala 76:16:@42244.4]
  assign regs_329_io_in = 64'h0; // @[RegFile.scala 75:16:@42243.4]
  assign regs_329_io_reset = reset; // @[RegFile.scala 78:19:@42247.4]
  assign regs_329_io_enable = 1'h1; // @[RegFile.scala 74:20:@42241.4]
  assign regs_330_clock = clock; // @[:@42250.4]
  assign regs_330_reset = io_reset; // @[:@42251.4 RegFile.scala 76:16:@42258.4]
  assign regs_330_io_in = 64'h0; // @[RegFile.scala 75:16:@42257.4]
  assign regs_330_io_reset = reset; // @[RegFile.scala 78:19:@42261.4]
  assign regs_330_io_enable = 1'h1; // @[RegFile.scala 74:20:@42255.4]
  assign regs_331_clock = clock; // @[:@42264.4]
  assign regs_331_reset = io_reset; // @[:@42265.4 RegFile.scala 76:16:@42272.4]
  assign regs_331_io_in = 64'h0; // @[RegFile.scala 75:16:@42271.4]
  assign regs_331_io_reset = reset; // @[RegFile.scala 78:19:@42275.4]
  assign regs_331_io_enable = 1'h1; // @[RegFile.scala 74:20:@42269.4]
  assign regs_332_clock = clock; // @[:@42278.4]
  assign regs_332_reset = io_reset; // @[:@42279.4 RegFile.scala 76:16:@42286.4]
  assign regs_332_io_in = 64'h0; // @[RegFile.scala 75:16:@42285.4]
  assign regs_332_io_reset = reset; // @[RegFile.scala 78:19:@42289.4]
  assign regs_332_io_enable = 1'h1; // @[RegFile.scala 74:20:@42283.4]
  assign regs_333_clock = clock; // @[:@42292.4]
  assign regs_333_reset = io_reset; // @[:@42293.4 RegFile.scala 76:16:@42300.4]
  assign regs_333_io_in = 64'h0; // @[RegFile.scala 75:16:@42299.4]
  assign regs_333_io_reset = reset; // @[RegFile.scala 78:19:@42303.4]
  assign regs_333_io_enable = 1'h1; // @[RegFile.scala 74:20:@42297.4]
  assign regs_334_clock = clock; // @[:@42306.4]
  assign regs_334_reset = io_reset; // @[:@42307.4 RegFile.scala 76:16:@42314.4]
  assign regs_334_io_in = 64'h0; // @[RegFile.scala 75:16:@42313.4]
  assign regs_334_io_reset = reset; // @[RegFile.scala 78:19:@42317.4]
  assign regs_334_io_enable = 1'h1; // @[RegFile.scala 74:20:@42311.4]
  assign regs_335_clock = clock; // @[:@42320.4]
  assign regs_335_reset = io_reset; // @[:@42321.4 RegFile.scala 76:16:@42328.4]
  assign regs_335_io_in = 64'h0; // @[RegFile.scala 75:16:@42327.4]
  assign regs_335_io_reset = reset; // @[RegFile.scala 78:19:@42331.4]
  assign regs_335_io_enable = 1'h1; // @[RegFile.scala 74:20:@42325.4]
  assign regs_336_clock = clock; // @[:@42334.4]
  assign regs_336_reset = io_reset; // @[:@42335.4 RegFile.scala 76:16:@42342.4]
  assign regs_336_io_in = 64'h0; // @[RegFile.scala 75:16:@42341.4]
  assign regs_336_io_reset = reset; // @[RegFile.scala 78:19:@42345.4]
  assign regs_336_io_enable = 1'h1; // @[RegFile.scala 74:20:@42339.4]
  assign regs_337_clock = clock; // @[:@42348.4]
  assign regs_337_reset = io_reset; // @[:@42349.4 RegFile.scala 76:16:@42356.4]
  assign regs_337_io_in = 64'h0; // @[RegFile.scala 75:16:@42355.4]
  assign regs_337_io_reset = reset; // @[RegFile.scala 78:19:@42359.4]
  assign regs_337_io_enable = 1'h1; // @[RegFile.scala 74:20:@42353.4]
  assign regs_338_clock = clock; // @[:@42362.4]
  assign regs_338_reset = io_reset; // @[:@42363.4 RegFile.scala 76:16:@42370.4]
  assign regs_338_io_in = 64'h0; // @[RegFile.scala 75:16:@42369.4]
  assign regs_338_io_reset = reset; // @[RegFile.scala 78:19:@42373.4]
  assign regs_338_io_enable = 1'h1; // @[RegFile.scala 74:20:@42367.4]
  assign regs_339_clock = clock; // @[:@42376.4]
  assign regs_339_reset = io_reset; // @[:@42377.4 RegFile.scala 76:16:@42384.4]
  assign regs_339_io_in = 64'h0; // @[RegFile.scala 75:16:@42383.4]
  assign regs_339_io_reset = reset; // @[RegFile.scala 78:19:@42387.4]
  assign regs_339_io_enable = 1'h1; // @[RegFile.scala 74:20:@42381.4]
  assign regs_340_clock = clock; // @[:@42390.4]
  assign regs_340_reset = io_reset; // @[:@42391.4 RegFile.scala 76:16:@42398.4]
  assign regs_340_io_in = 64'h0; // @[RegFile.scala 75:16:@42397.4]
  assign regs_340_io_reset = reset; // @[RegFile.scala 78:19:@42401.4]
  assign regs_340_io_enable = 1'h1; // @[RegFile.scala 74:20:@42395.4]
  assign regs_341_clock = clock; // @[:@42404.4]
  assign regs_341_reset = io_reset; // @[:@42405.4 RegFile.scala 76:16:@42412.4]
  assign regs_341_io_in = 64'h0; // @[RegFile.scala 75:16:@42411.4]
  assign regs_341_io_reset = reset; // @[RegFile.scala 78:19:@42415.4]
  assign regs_341_io_enable = 1'h1; // @[RegFile.scala 74:20:@42409.4]
  assign regs_342_clock = clock; // @[:@42418.4]
  assign regs_342_reset = io_reset; // @[:@42419.4 RegFile.scala 76:16:@42426.4]
  assign regs_342_io_in = 64'h0; // @[RegFile.scala 75:16:@42425.4]
  assign regs_342_io_reset = reset; // @[RegFile.scala 78:19:@42429.4]
  assign regs_342_io_enable = 1'h1; // @[RegFile.scala 74:20:@42423.4]
  assign regs_343_clock = clock; // @[:@42432.4]
  assign regs_343_reset = io_reset; // @[:@42433.4 RegFile.scala 76:16:@42440.4]
  assign regs_343_io_in = 64'h0; // @[RegFile.scala 75:16:@42439.4]
  assign regs_343_io_reset = reset; // @[RegFile.scala 78:19:@42443.4]
  assign regs_343_io_enable = 1'h1; // @[RegFile.scala 74:20:@42437.4]
  assign regs_344_clock = clock; // @[:@42446.4]
  assign regs_344_reset = io_reset; // @[:@42447.4 RegFile.scala 76:16:@42454.4]
  assign regs_344_io_in = 64'h0; // @[RegFile.scala 75:16:@42453.4]
  assign regs_344_io_reset = reset; // @[RegFile.scala 78:19:@42457.4]
  assign regs_344_io_enable = 1'h1; // @[RegFile.scala 74:20:@42451.4]
  assign regs_345_clock = clock; // @[:@42460.4]
  assign regs_345_reset = io_reset; // @[:@42461.4 RegFile.scala 76:16:@42468.4]
  assign regs_345_io_in = 64'h0; // @[RegFile.scala 75:16:@42467.4]
  assign regs_345_io_reset = reset; // @[RegFile.scala 78:19:@42471.4]
  assign regs_345_io_enable = 1'h1; // @[RegFile.scala 74:20:@42465.4]
  assign regs_346_clock = clock; // @[:@42474.4]
  assign regs_346_reset = io_reset; // @[:@42475.4 RegFile.scala 76:16:@42482.4]
  assign regs_346_io_in = 64'h0; // @[RegFile.scala 75:16:@42481.4]
  assign regs_346_io_reset = reset; // @[RegFile.scala 78:19:@42485.4]
  assign regs_346_io_enable = 1'h1; // @[RegFile.scala 74:20:@42479.4]
  assign regs_347_clock = clock; // @[:@42488.4]
  assign regs_347_reset = io_reset; // @[:@42489.4 RegFile.scala 76:16:@42496.4]
  assign regs_347_io_in = 64'h0; // @[RegFile.scala 75:16:@42495.4]
  assign regs_347_io_reset = reset; // @[RegFile.scala 78:19:@42499.4]
  assign regs_347_io_enable = 1'h1; // @[RegFile.scala 74:20:@42493.4]
  assign regs_348_clock = clock; // @[:@42502.4]
  assign regs_348_reset = io_reset; // @[:@42503.4 RegFile.scala 76:16:@42510.4]
  assign regs_348_io_in = 64'h0; // @[RegFile.scala 75:16:@42509.4]
  assign regs_348_io_reset = reset; // @[RegFile.scala 78:19:@42513.4]
  assign regs_348_io_enable = 1'h1; // @[RegFile.scala 74:20:@42507.4]
  assign regs_349_clock = clock; // @[:@42516.4]
  assign regs_349_reset = io_reset; // @[:@42517.4 RegFile.scala 76:16:@42524.4]
  assign regs_349_io_in = 64'h0; // @[RegFile.scala 75:16:@42523.4]
  assign regs_349_io_reset = reset; // @[RegFile.scala 78:19:@42527.4]
  assign regs_349_io_enable = 1'h1; // @[RegFile.scala 74:20:@42521.4]
  assign regs_350_clock = clock; // @[:@42530.4]
  assign regs_350_reset = io_reset; // @[:@42531.4 RegFile.scala 76:16:@42538.4]
  assign regs_350_io_in = 64'h0; // @[RegFile.scala 75:16:@42537.4]
  assign regs_350_io_reset = reset; // @[RegFile.scala 78:19:@42541.4]
  assign regs_350_io_enable = 1'h1; // @[RegFile.scala 74:20:@42535.4]
  assign regs_351_clock = clock; // @[:@42544.4]
  assign regs_351_reset = io_reset; // @[:@42545.4 RegFile.scala 76:16:@42552.4]
  assign regs_351_io_in = 64'h0; // @[RegFile.scala 75:16:@42551.4]
  assign regs_351_io_reset = reset; // @[RegFile.scala 78:19:@42555.4]
  assign regs_351_io_enable = 1'h1; // @[RegFile.scala 74:20:@42549.4]
  assign regs_352_clock = clock; // @[:@42558.4]
  assign regs_352_reset = io_reset; // @[:@42559.4 RegFile.scala 76:16:@42566.4]
  assign regs_352_io_in = 64'h0; // @[RegFile.scala 75:16:@42565.4]
  assign regs_352_io_reset = reset; // @[RegFile.scala 78:19:@42569.4]
  assign regs_352_io_enable = 1'h1; // @[RegFile.scala 74:20:@42563.4]
  assign regs_353_clock = clock; // @[:@42572.4]
  assign regs_353_reset = io_reset; // @[:@42573.4 RegFile.scala 76:16:@42580.4]
  assign regs_353_io_in = 64'h0; // @[RegFile.scala 75:16:@42579.4]
  assign regs_353_io_reset = reset; // @[RegFile.scala 78:19:@42583.4]
  assign regs_353_io_enable = 1'h1; // @[RegFile.scala 74:20:@42577.4]
  assign regs_354_clock = clock; // @[:@42586.4]
  assign regs_354_reset = io_reset; // @[:@42587.4 RegFile.scala 76:16:@42594.4]
  assign regs_354_io_in = 64'h0; // @[RegFile.scala 75:16:@42593.4]
  assign regs_354_io_reset = reset; // @[RegFile.scala 78:19:@42597.4]
  assign regs_354_io_enable = 1'h1; // @[RegFile.scala 74:20:@42591.4]
  assign regs_355_clock = clock; // @[:@42600.4]
  assign regs_355_reset = io_reset; // @[:@42601.4 RegFile.scala 76:16:@42608.4]
  assign regs_355_io_in = 64'h0; // @[RegFile.scala 75:16:@42607.4]
  assign regs_355_io_reset = reset; // @[RegFile.scala 78:19:@42611.4]
  assign regs_355_io_enable = 1'h1; // @[RegFile.scala 74:20:@42605.4]
  assign regs_356_clock = clock; // @[:@42614.4]
  assign regs_356_reset = io_reset; // @[:@42615.4 RegFile.scala 76:16:@42622.4]
  assign regs_356_io_in = 64'h0; // @[RegFile.scala 75:16:@42621.4]
  assign regs_356_io_reset = reset; // @[RegFile.scala 78:19:@42625.4]
  assign regs_356_io_enable = 1'h1; // @[RegFile.scala 74:20:@42619.4]
  assign regs_357_clock = clock; // @[:@42628.4]
  assign regs_357_reset = io_reset; // @[:@42629.4 RegFile.scala 76:16:@42636.4]
  assign regs_357_io_in = 64'h0; // @[RegFile.scala 75:16:@42635.4]
  assign regs_357_io_reset = reset; // @[RegFile.scala 78:19:@42639.4]
  assign regs_357_io_enable = 1'h1; // @[RegFile.scala 74:20:@42633.4]
  assign regs_358_clock = clock; // @[:@42642.4]
  assign regs_358_reset = io_reset; // @[:@42643.4 RegFile.scala 76:16:@42650.4]
  assign regs_358_io_in = 64'h0; // @[RegFile.scala 75:16:@42649.4]
  assign regs_358_io_reset = reset; // @[RegFile.scala 78:19:@42653.4]
  assign regs_358_io_enable = 1'h1; // @[RegFile.scala 74:20:@42647.4]
  assign regs_359_clock = clock; // @[:@42656.4]
  assign regs_359_reset = io_reset; // @[:@42657.4 RegFile.scala 76:16:@42664.4]
  assign regs_359_io_in = 64'h0; // @[RegFile.scala 75:16:@42663.4]
  assign regs_359_io_reset = reset; // @[RegFile.scala 78:19:@42667.4]
  assign regs_359_io_enable = 1'h1; // @[RegFile.scala 74:20:@42661.4]
  assign regs_360_clock = clock; // @[:@42670.4]
  assign regs_360_reset = io_reset; // @[:@42671.4 RegFile.scala 76:16:@42678.4]
  assign regs_360_io_in = 64'h0; // @[RegFile.scala 75:16:@42677.4]
  assign regs_360_io_reset = reset; // @[RegFile.scala 78:19:@42681.4]
  assign regs_360_io_enable = 1'h1; // @[RegFile.scala 74:20:@42675.4]
  assign regs_361_clock = clock; // @[:@42684.4]
  assign regs_361_reset = io_reset; // @[:@42685.4 RegFile.scala 76:16:@42692.4]
  assign regs_361_io_in = 64'h0; // @[RegFile.scala 75:16:@42691.4]
  assign regs_361_io_reset = reset; // @[RegFile.scala 78:19:@42695.4]
  assign regs_361_io_enable = 1'h1; // @[RegFile.scala 74:20:@42689.4]
  assign regs_362_clock = clock; // @[:@42698.4]
  assign regs_362_reset = io_reset; // @[:@42699.4 RegFile.scala 76:16:@42706.4]
  assign regs_362_io_in = 64'h0; // @[RegFile.scala 75:16:@42705.4]
  assign regs_362_io_reset = reset; // @[RegFile.scala 78:19:@42709.4]
  assign regs_362_io_enable = 1'h1; // @[RegFile.scala 74:20:@42703.4]
  assign regs_363_clock = clock; // @[:@42712.4]
  assign regs_363_reset = io_reset; // @[:@42713.4 RegFile.scala 76:16:@42720.4]
  assign regs_363_io_in = 64'h0; // @[RegFile.scala 75:16:@42719.4]
  assign regs_363_io_reset = reset; // @[RegFile.scala 78:19:@42723.4]
  assign regs_363_io_enable = 1'h1; // @[RegFile.scala 74:20:@42717.4]
  assign regs_364_clock = clock; // @[:@42726.4]
  assign regs_364_reset = io_reset; // @[:@42727.4 RegFile.scala 76:16:@42734.4]
  assign regs_364_io_in = 64'h0; // @[RegFile.scala 75:16:@42733.4]
  assign regs_364_io_reset = reset; // @[RegFile.scala 78:19:@42737.4]
  assign regs_364_io_enable = 1'h1; // @[RegFile.scala 74:20:@42731.4]
  assign regs_365_clock = clock; // @[:@42740.4]
  assign regs_365_reset = io_reset; // @[:@42741.4 RegFile.scala 76:16:@42748.4]
  assign regs_365_io_in = 64'h0; // @[RegFile.scala 75:16:@42747.4]
  assign regs_365_io_reset = reset; // @[RegFile.scala 78:19:@42751.4]
  assign regs_365_io_enable = 1'h1; // @[RegFile.scala 74:20:@42745.4]
  assign regs_366_clock = clock; // @[:@42754.4]
  assign regs_366_reset = io_reset; // @[:@42755.4 RegFile.scala 76:16:@42762.4]
  assign regs_366_io_in = 64'h0; // @[RegFile.scala 75:16:@42761.4]
  assign regs_366_io_reset = reset; // @[RegFile.scala 78:19:@42765.4]
  assign regs_366_io_enable = 1'h1; // @[RegFile.scala 74:20:@42759.4]
  assign regs_367_clock = clock; // @[:@42768.4]
  assign regs_367_reset = io_reset; // @[:@42769.4 RegFile.scala 76:16:@42776.4]
  assign regs_367_io_in = 64'h0; // @[RegFile.scala 75:16:@42775.4]
  assign regs_367_io_reset = reset; // @[RegFile.scala 78:19:@42779.4]
  assign regs_367_io_enable = 1'h1; // @[RegFile.scala 74:20:@42773.4]
  assign regs_368_clock = clock; // @[:@42782.4]
  assign regs_368_reset = io_reset; // @[:@42783.4 RegFile.scala 76:16:@42790.4]
  assign regs_368_io_in = 64'h0; // @[RegFile.scala 75:16:@42789.4]
  assign regs_368_io_reset = reset; // @[RegFile.scala 78:19:@42793.4]
  assign regs_368_io_enable = 1'h1; // @[RegFile.scala 74:20:@42787.4]
  assign regs_369_clock = clock; // @[:@42796.4]
  assign regs_369_reset = io_reset; // @[:@42797.4 RegFile.scala 76:16:@42804.4]
  assign regs_369_io_in = 64'h0; // @[RegFile.scala 75:16:@42803.4]
  assign regs_369_io_reset = reset; // @[RegFile.scala 78:19:@42807.4]
  assign regs_369_io_enable = 1'h1; // @[RegFile.scala 74:20:@42801.4]
  assign regs_370_clock = clock; // @[:@42810.4]
  assign regs_370_reset = io_reset; // @[:@42811.4 RegFile.scala 76:16:@42818.4]
  assign regs_370_io_in = 64'h0; // @[RegFile.scala 75:16:@42817.4]
  assign regs_370_io_reset = reset; // @[RegFile.scala 78:19:@42821.4]
  assign regs_370_io_enable = 1'h1; // @[RegFile.scala 74:20:@42815.4]
  assign regs_371_clock = clock; // @[:@42824.4]
  assign regs_371_reset = io_reset; // @[:@42825.4 RegFile.scala 76:16:@42832.4]
  assign regs_371_io_in = 64'h0; // @[RegFile.scala 75:16:@42831.4]
  assign regs_371_io_reset = reset; // @[RegFile.scala 78:19:@42835.4]
  assign regs_371_io_enable = 1'h1; // @[RegFile.scala 74:20:@42829.4]
  assign regs_372_clock = clock; // @[:@42838.4]
  assign regs_372_reset = io_reset; // @[:@42839.4 RegFile.scala 76:16:@42846.4]
  assign regs_372_io_in = 64'h0; // @[RegFile.scala 75:16:@42845.4]
  assign regs_372_io_reset = reset; // @[RegFile.scala 78:19:@42849.4]
  assign regs_372_io_enable = 1'h1; // @[RegFile.scala 74:20:@42843.4]
  assign regs_373_clock = clock; // @[:@42852.4]
  assign regs_373_reset = io_reset; // @[:@42853.4 RegFile.scala 76:16:@42860.4]
  assign regs_373_io_in = 64'h0; // @[RegFile.scala 75:16:@42859.4]
  assign regs_373_io_reset = reset; // @[RegFile.scala 78:19:@42863.4]
  assign regs_373_io_enable = 1'h1; // @[RegFile.scala 74:20:@42857.4]
  assign regs_374_clock = clock; // @[:@42866.4]
  assign regs_374_reset = io_reset; // @[:@42867.4 RegFile.scala 76:16:@42874.4]
  assign regs_374_io_in = 64'h0; // @[RegFile.scala 75:16:@42873.4]
  assign regs_374_io_reset = reset; // @[RegFile.scala 78:19:@42877.4]
  assign regs_374_io_enable = 1'h1; // @[RegFile.scala 74:20:@42871.4]
  assign regs_375_clock = clock; // @[:@42880.4]
  assign regs_375_reset = io_reset; // @[:@42881.4 RegFile.scala 76:16:@42888.4]
  assign regs_375_io_in = 64'h0; // @[RegFile.scala 75:16:@42887.4]
  assign regs_375_io_reset = reset; // @[RegFile.scala 78:19:@42891.4]
  assign regs_375_io_enable = 1'h1; // @[RegFile.scala 74:20:@42885.4]
  assign regs_376_clock = clock; // @[:@42894.4]
  assign regs_376_reset = io_reset; // @[:@42895.4 RegFile.scala 76:16:@42902.4]
  assign regs_376_io_in = 64'h0; // @[RegFile.scala 75:16:@42901.4]
  assign regs_376_io_reset = reset; // @[RegFile.scala 78:19:@42905.4]
  assign regs_376_io_enable = 1'h1; // @[RegFile.scala 74:20:@42899.4]
  assign regs_377_clock = clock; // @[:@42908.4]
  assign regs_377_reset = io_reset; // @[:@42909.4 RegFile.scala 76:16:@42916.4]
  assign regs_377_io_in = 64'h0; // @[RegFile.scala 75:16:@42915.4]
  assign regs_377_io_reset = reset; // @[RegFile.scala 78:19:@42919.4]
  assign regs_377_io_enable = 1'h1; // @[RegFile.scala 74:20:@42913.4]
  assign regs_378_clock = clock; // @[:@42922.4]
  assign regs_378_reset = io_reset; // @[:@42923.4 RegFile.scala 76:16:@42930.4]
  assign regs_378_io_in = 64'h0; // @[RegFile.scala 75:16:@42929.4]
  assign regs_378_io_reset = reset; // @[RegFile.scala 78:19:@42933.4]
  assign regs_378_io_enable = 1'h1; // @[RegFile.scala 74:20:@42927.4]
  assign regs_379_clock = clock; // @[:@42936.4]
  assign regs_379_reset = io_reset; // @[:@42937.4 RegFile.scala 76:16:@42944.4]
  assign regs_379_io_in = 64'h0; // @[RegFile.scala 75:16:@42943.4]
  assign regs_379_io_reset = reset; // @[RegFile.scala 78:19:@42947.4]
  assign regs_379_io_enable = 1'h1; // @[RegFile.scala 74:20:@42941.4]
  assign regs_380_clock = clock; // @[:@42950.4]
  assign regs_380_reset = io_reset; // @[:@42951.4 RegFile.scala 76:16:@42958.4]
  assign regs_380_io_in = 64'h0; // @[RegFile.scala 75:16:@42957.4]
  assign regs_380_io_reset = reset; // @[RegFile.scala 78:19:@42961.4]
  assign regs_380_io_enable = 1'h1; // @[RegFile.scala 74:20:@42955.4]
  assign regs_381_clock = clock; // @[:@42964.4]
  assign regs_381_reset = io_reset; // @[:@42965.4 RegFile.scala 76:16:@42972.4]
  assign regs_381_io_in = 64'h0; // @[RegFile.scala 75:16:@42971.4]
  assign regs_381_io_reset = reset; // @[RegFile.scala 78:19:@42975.4]
  assign regs_381_io_enable = 1'h1; // @[RegFile.scala 74:20:@42969.4]
  assign regs_382_clock = clock; // @[:@42978.4]
  assign regs_382_reset = io_reset; // @[:@42979.4 RegFile.scala 76:16:@42986.4]
  assign regs_382_io_in = 64'h0; // @[RegFile.scala 75:16:@42985.4]
  assign regs_382_io_reset = reset; // @[RegFile.scala 78:19:@42989.4]
  assign regs_382_io_enable = 1'h1; // @[RegFile.scala 74:20:@42983.4]
  assign regs_383_clock = clock; // @[:@42992.4]
  assign regs_383_reset = io_reset; // @[:@42993.4 RegFile.scala 76:16:@43000.4]
  assign regs_383_io_in = 64'h0; // @[RegFile.scala 75:16:@42999.4]
  assign regs_383_io_reset = reset; // @[RegFile.scala 78:19:@43003.4]
  assign regs_383_io_enable = 1'h1; // @[RegFile.scala 74:20:@42997.4]
  assign regs_384_clock = clock; // @[:@43006.4]
  assign regs_384_reset = io_reset; // @[:@43007.4 RegFile.scala 76:16:@43014.4]
  assign regs_384_io_in = 64'h0; // @[RegFile.scala 75:16:@43013.4]
  assign regs_384_io_reset = reset; // @[RegFile.scala 78:19:@43017.4]
  assign regs_384_io_enable = 1'h1; // @[RegFile.scala 74:20:@43011.4]
  assign regs_385_clock = clock; // @[:@43020.4]
  assign regs_385_reset = io_reset; // @[:@43021.4 RegFile.scala 76:16:@43028.4]
  assign regs_385_io_in = 64'h0; // @[RegFile.scala 75:16:@43027.4]
  assign regs_385_io_reset = reset; // @[RegFile.scala 78:19:@43031.4]
  assign regs_385_io_enable = 1'h1; // @[RegFile.scala 74:20:@43025.4]
  assign regs_386_clock = clock; // @[:@43034.4]
  assign regs_386_reset = io_reset; // @[:@43035.4 RegFile.scala 76:16:@43042.4]
  assign regs_386_io_in = 64'h0; // @[RegFile.scala 75:16:@43041.4]
  assign regs_386_io_reset = reset; // @[RegFile.scala 78:19:@43045.4]
  assign regs_386_io_enable = 1'h1; // @[RegFile.scala 74:20:@43039.4]
  assign regs_387_clock = clock; // @[:@43048.4]
  assign regs_387_reset = io_reset; // @[:@43049.4 RegFile.scala 76:16:@43056.4]
  assign regs_387_io_in = 64'h0; // @[RegFile.scala 75:16:@43055.4]
  assign regs_387_io_reset = reset; // @[RegFile.scala 78:19:@43059.4]
  assign regs_387_io_enable = 1'h1; // @[RegFile.scala 74:20:@43053.4]
  assign regs_388_clock = clock; // @[:@43062.4]
  assign regs_388_reset = io_reset; // @[:@43063.4 RegFile.scala 76:16:@43070.4]
  assign regs_388_io_in = 64'h0; // @[RegFile.scala 75:16:@43069.4]
  assign regs_388_io_reset = reset; // @[RegFile.scala 78:19:@43073.4]
  assign regs_388_io_enable = 1'h1; // @[RegFile.scala 74:20:@43067.4]
  assign regs_389_clock = clock; // @[:@43076.4]
  assign regs_389_reset = io_reset; // @[:@43077.4 RegFile.scala 76:16:@43084.4]
  assign regs_389_io_in = 64'h0; // @[RegFile.scala 75:16:@43083.4]
  assign regs_389_io_reset = reset; // @[RegFile.scala 78:19:@43087.4]
  assign regs_389_io_enable = 1'h1; // @[RegFile.scala 74:20:@43081.4]
  assign regs_390_clock = clock; // @[:@43090.4]
  assign regs_390_reset = io_reset; // @[:@43091.4 RegFile.scala 76:16:@43098.4]
  assign regs_390_io_in = 64'h0; // @[RegFile.scala 75:16:@43097.4]
  assign regs_390_io_reset = reset; // @[RegFile.scala 78:19:@43101.4]
  assign regs_390_io_enable = 1'h1; // @[RegFile.scala 74:20:@43095.4]
  assign regs_391_clock = clock; // @[:@43104.4]
  assign regs_391_reset = io_reset; // @[:@43105.4 RegFile.scala 76:16:@43112.4]
  assign regs_391_io_in = 64'h0; // @[RegFile.scala 75:16:@43111.4]
  assign regs_391_io_reset = reset; // @[RegFile.scala 78:19:@43115.4]
  assign regs_391_io_enable = 1'h1; // @[RegFile.scala 74:20:@43109.4]
  assign regs_392_clock = clock; // @[:@43118.4]
  assign regs_392_reset = io_reset; // @[:@43119.4 RegFile.scala 76:16:@43126.4]
  assign regs_392_io_in = 64'h0; // @[RegFile.scala 75:16:@43125.4]
  assign regs_392_io_reset = reset; // @[RegFile.scala 78:19:@43129.4]
  assign regs_392_io_enable = 1'h1; // @[RegFile.scala 74:20:@43123.4]
  assign regs_393_clock = clock; // @[:@43132.4]
  assign regs_393_reset = io_reset; // @[:@43133.4 RegFile.scala 76:16:@43140.4]
  assign regs_393_io_in = 64'h0; // @[RegFile.scala 75:16:@43139.4]
  assign regs_393_io_reset = reset; // @[RegFile.scala 78:19:@43143.4]
  assign regs_393_io_enable = 1'h1; // @[RegFile.scala 74:20:@43137.4]
  assign regs_394_clock = clock; // @[:@43146.4]
  assign regs_394_reset = io_reset; // @[:@43147.4 RegFile.scala 76:16:@43154.4]
  assign regs_394_io_in = 64'h0; // @[RegFile.scala 75:16:@43153.4]
  assign regs_394_io_reset = reset; // @[RegFile.scala 78:19:@43157.4]
  assign regs_394_io_enable = 1'h1; // @[RegFile.scala 74:20:@43151.4]
  assign regs_395_clock = clock; // @[:@43160.4]
  assign regs_395_reset = io_reset; // @[:@43161.4 RegFile.scala 76:16:@43168.4]
  assign regs_395_io_in = 64'h0; // @[RegFile.scala 75:16:@43167.4]
  assign regs_395_io_reset = reset; // @[RegFile.scala 78:19:@43171.4]
  assign regs_395_io_enable = 1'h1; // @[RegFile.scala 74:20:@43165.4]
  assign regs_396_clock = clock; // @[:@43174.4]
  assign regs_396_reset = io_reset; // @[:@43175.4 RegFile.scala 76:16:@43182.4]
  assign regs_396_io_in = 64'h0; // @[RegFile.scala 75:16:@43181.4]
  assign regs_396_io_reset = reset; // @[RegFile.scala 78:19:@43185.4]
  assign regs_396_io_enable = 1'h1; // @[RegFile.scala 74:20:@43179.4]
  assign regs_397_clock = clock; // @[:@43188.4]
  assign regs_397_reset = io_reset; // @[:@43189.4 RegFile.scala 76:16:@43196.4]
  assign regs_397_io_in = 64'h0; // @[RegFile.scala 75:16:@43195.4]
  assign regs_397_io_reset = reset; // @[RegFile.scala 78:19:@43199.4]
  assign regs_397_io_enable = 1'h1; // @[RegFile.scala 74:20:@43193.4]
  assign regs_398_clock = clock; // @[:@43202.4]
  assign regs_398_reset = io_reset; // @[:@43203.4 RegFile.scala 76:16:@43210.4]
  assign regs_398_io_in = 64'h0; // @[RegFile.scala 75:16:@43209.4]
  assign regs_398_io_reset = reset; // @[RegFile.scala 78:19:@43213.4]
  assign regs_398_io_enable = 1'h1; // @[RegFile.scala 74:20:@43207.4]
  assign regs_399_clock = clock; // @[:@43216.4]
  assign regs_399_reset = io_reset; // @[:@43217.4 RegFile.scala 76:16:@43224.4]
  assign regs_399_io_in = 64'h0; // @[RegFile.scala 75:16:@43223.4]
  assign regs_399_io_reset = reset; // @[RegFile.scala 78:19:@43227.4]
  assign regs_399_io_enable = 1'h1; // @[RegFile.scala 74:20:@43221.4]
  assign regs_400_clock = clock; // @[:@43230.4]
  assign regs_400_reset = io_reset; // @[:@43231.4 RegFile.scala 76:16:@43238.4]
  assign regs_400_io_in = 64'h0; // @[RegFile.scala 75:16:@43237.4]
  assign regs_400_io_reset = reset; // @[RegFile.scala 78:19:@43241.4]
  assign regs_400_io_enable = 1'h1; // @[RegFile.scala 74:20:@43235.4]
  assign regs_401_clock = clock; // @[:@43244.4]
  assign regs_401_reset = io_reset; // @[:@43245.4 RegFile.scala 76:16:@43252.4]
  assign regs_401_io_in = 64'h0; // @[RegFile.scala 75:16:@43251.4]
  assign regs_401_io_reset = reset; // @[RegFile.scala 78:19:@43255.4]
  assign regs_401_io_enable = 1'h1; // @[RegFile.scala 74:20:@43249.4]
  assign regs_402_clock = clock; // @[:@43258.4]
  assign regs_402_reset = io_reset; // @[:@43259.4 RegFile.scala 76:16:@43266.4]
  assign regs_402_io_in = 64'h0; // @[RegFile.scala 75:16:@43265.4]
  assign regs_402_io_reset = reset; // @[RegFile.scala 78:19:@43269.4]
  assign regs_402_io_enable = 1'h1; // @[RegFile.scala 74:20:@43263.4]
  assign regs_403_clock = clock; // @[:@43272.4]
  assign regs_403_reset = io_reset; // @[:@43273.4 RegFile.scala 76:16:@43280.4]
  assign regs_403_io_in = 64'h0; // @[RegFile.scala 75:16:@43279.4]
  assign regs_403_io_reset = reset; // @[RegFile.scala 78:19:@43283.4]
  assign regs_403_io_enable = 1'h1; // @[RegFile.scala 74:20:@43277.4]
  assign regs_404_clock = clock; // @[:@43286.4]
  assign regs_404_reset = io_reset; // @[:@43287.4 RegFile.scala 76:16:@43294.4]
  assign regs_404_io_in = 64'h0; // @[RegFile.scala 75:16:@43293.4]
  assign regs_404_io_reset = reset; // @[RegFile.scala 78:19:@43297.4]
  assign regs_404_io_enable = 1'h1; // @[RegFile.scala 74:20:@43291.4]
  assign regs_405_clock = clock; // @[:@43300.4]
  assign regs_405_reset = io_reset; // @[:@43301.4 RegFile.scala 76:16:@43308.4]
  assign regs_405_io_in = 64'h0; // @[RegFile.scala 75:16:@43307.4]
  assign regs_405_io_reset = reset; // @[RegFile.scala 78:19:@43311.4]
  assign regs_405_io_enable = 1'h1; // @[RegFile.scala 74:20:@43305.4]
  assign regs_406_clock = clock; // @[:@43314.4]
  assign regs_406_reset = io_reset; // @[:@43315.4 RegFile.scala 76:16:@43322.4]
  assign regs_406_io_in = 64'h0; // @[RegFile.scala 75:16:@43321.4]
  assign regs_406_io_reset = reset; // @[RegFile.scala 78:19:@43325.4]
  assign regs_406_io_enable = 1'h1; // @[RegFile.scala 74:20:@43319.4]
  assign regs_407_clock = clock; // @[:@43328.4]
  assign regs_407_reset = io_reset; // @[:@43329.4 RegFile.scala 76:16:@43336.4]
  assign regs_407_io_in = 64'h0; // @[RegFile.scala 75:16:@43335.4]
  assign regs_407_io_reset = reset; // @[RegFile.scala 78:19:@43339.4]
  assign regs_407_io_enable = 1'h1; // @[RegFile.scala 74:20:@43333.4]
  assign regs_408_clock = clock; // @[:@43342.4]
  assign regs_408_reset = io_reset; // @[:@43343.4 RegFile.scala 76:16:@43350.4]
  assign regs_408_io_in = 64'h0; // @[RegFile.scala 75:16:@43349.4]
  assign regs_408_io_reset = reset; // @[RegFile.scala 78:19:@43353.4]
  assign regs_408_io_enable = 1'h1; // @[RegFile.scala 74:20:@43347.4]
  assign regs_409_clock = clock; // @[:@43356.4]
  assign regs_409_reset = io_reset; // @[:@43357.4 RegFile.scala 76:16:@43364.4]
  assign regs_409_io_in = 64'h0; // @[RegFile.scala 75:16:@43363.4]
  assign regs_409_io_reset = reset; // @[RegFile.scala 78:19:@43367.4]
  assign regs_409_io_enable = 1'h1; // @[RegFile.scala 74:20:@43361.4]
  assign regs_410_clock = clock; // @[:@43370.4]
  assign regs_410_reset = io_reset; // @[:@43371.4 RegFile.scala 76:16:@43378.4]
  assign regs_410_io_in = 64'h0; // @[RegFile.scala 75:16:@43377.4]
  assign regs_410_io_reset = reset; // @[RegFile.scala 78:19:@43381.4]
  assign regs_410_io_enable = 1'h1; // @[RegFile.scala 74:20:@43375.4]
  assign regs_411_clock = clock; // @[:@43384.4]
  assign regs_411_reset = io_reset; // @[:@43385.4 RegFile.scala 76:16:@43392.4]
  assign regs_411_io_in = 64'h0; // @[RegFile.scala 75:16:@43391.4]
  assign regs_411_io_reset = reset; // @[RegFile.scala 78:19:@43395.4]
  assign regs_411_io_enable = 1'h1; // @[RegFile.scala 74:20:@43389.4]
  assign regs_412_clock = clock; // @[:@43398.4]
  assign regs_412_reset = io_reset; // @[:@43399.4 RegFile.scala 76:16:@43406.4]
  assign regs_412_io_in = 64'h0; // @[RegFile.scala 75:16:@43405.4]
  assign regs_412_io_reset = reset; // @[RegFile.scala 78:19:@43409.4]
  assign regs_412_io_enable = 1'h1; // @[RegFile.scala 74:20:@43403.4]
  assign regs_413_clock = clock; // @[:@43412.4]
  assign regs_413_reset = io_reset; // @[:@43413.4 RegFile.scala 76:16:@43420.4]
  assign regs_413_io_in = 64'h0; // @[RegFile.scala 75:16:@43419.4]
  assign regs_413_io_reset = reset; // @[RegFile.scala 78:19:@43423.4]
  assign regs_413_io_enable = 1'h1; // @[RegFile.scala 74:20:@43417.4]
  assign regs_414_clock = clock; // @[:@43426.4]
  assign regs_414_reset = io_reset; // @[:@43427.4 RegFile.scala 76:16:@43434.4]
  assign regs_414_io_in = 64'h0; // @[RegFile.scala 75:16:@43433.4]
  assign regs_414_io_reset = reset; // @[RegFile.scala 78:19:@43437.4]
  assign regs_414_io_enable = 1'h1; // @[RegFile.scala 74:20:@43431.4]
  assign regs_415_clock = clock; // @[:@43440.4]
  assign regs_415_reset = io_reset; // @[:@43441.4 RegFile.scala 76:16:@43448.4]
  assign regs_415_io_in = 64'h0; // @[RegFile.scala 75:16:@43447.4]
  assign regs_415_io_reset = reset; // @[RegFile.scala 78:19:@43451.4]
  assign regs_415_io_enable = 1'h1; // @[RegFile.scala 74:20:@43445.4]
  assign regs_416_clock = clock; // @[:@43454.4]
  assign regs_416_reset = io_reset; // @[:@43455.4 RegFile.scala 76:16:@43462.4]
  assign regs_416_io_in = 64'h0; // @[RegFile.scala 75:16:@43461.4]
  assign regs_416_io_reset = reset; // @[RegFile.scala 78:19:@43465.4]
  assign regs_416_io_enable = 1'h1; // @[RegFile.scala 74:20:@43459.4]
  assign regs_417_clock = clock; // @[:@43468.4]
  assign regs_417_reset = io_reset; // @[:@43469.4 RegFile.scala 76:16:@43476.4]
  assign regs_417_io_in = 64'h0; // @[RegFile.scala 75:16:@43475.4]
  assign regs_417_io_reset = reset; // @[RegFile.scala 78:19:@43479.4]
  assign regs_417_io_enable = 1'h1; // @[RegFile.scala 74:20:@43473.4]
  assign regs_418_clock = clock; // @[:@43482.4]
  assign regs_418_reset = io_reset; // @[:@43483.4 RegFile.scala 76:16:@43490.4]
  assign regs_418_io_in = 64'h0; // @[RegFile.scala 75:16:@43489.4]
  assign regs_418_io_reset = reset; // @[RegFile.scala 78:19:@43493.4]
  assign regs_418_io_enable = 1'h1; // @[RegFile.scala 74:20:@43487.4]
  assign regs_419_clock = clock; // @[:@43496.4]
  assign regs_419_reset = io_reset; // @[:@43497.4 RegFile.scala 76:16:@43504.4]
  assign regs_419_io_in = 64'h0; // @[RegFile.scala 75:16:@43503.4]
  assign regs_419_io_reset = reset; // @[RegFile.scala 78:19:@43507.4]
  assign regs_419_io_enable = 1'h1; // @[RegFile.scala 74:20:@43501.4]
  assign regs_420_clock = clock; // @[:@43510.4]
  assign regs_420_reset = io_reset; // @[:@43511.4 RegFile.scala 76:16:@43518.4]
  assign regs_420_io_in = 64'h0; // @[RegFile.scala 75:16:@43517.4]
  assign regs_420_io_reset = reset; // @[RegFile.scala 78:19:@43521.4]
  assign regs_420_io_enable = 1'h1; // @[RegFile.scala 74:20:@43515.4]
  assign regs_421_clock = clock; // @[:@43524.4]
  assign regs_421_reset = io_reset; // @[:@43525.4 RegFile.scala 76:16:@43532.4]
  assign regs_421_io_in = 64'h0; // @[RegFile.scala 75:16:@43531.4]
  assign regs_421_io_reset = reset; // @[RegFile.scala 78:19:@43535.4]
  assign regs_421_io_enable = 1'h1; // @[RegFile.scala 74:20:@43529.4]
  assign regs_422_clock = clock; // @[:@43538.4]
  assign regs_422_reset = io_reset; // @[:@43539.4 RegFile.scala 76:16:@43546.4]
  assign regs_422_io_in = 64'h0; // @[RegFile.scala 75:16:@43545.4]
  assign regs_422_io_reset = reset; // @[RegFile.scala 78:19:@43549.4]
  assign regs_422_io_enable = 1'h1; // @[RegFile.scala 74:20:@43543.4]
  assign regs_423_clock = clock; // @[:@43552.4]
  assign regs_423_reset = io_reset; // @[:@43553.4 RegFile.scala 76:16:@43560.4]
  assign regs_423_io_in = 64'h0; // @[RegFile.scala 75:16:@43559.4]
  assign regs_423_io_reset = reset; // @[RegFile.scala 78:19:@43563.4]
  assign regs_423_io_enable = 1'h1; // @[RegFile.scala 74:20:@43557.4]
  assign regs_424_clock = clock; // @[:@43566.4]
  assign regs_424_reset = io_reset; // @[:@43567.4 RegFile.scala 76:16:@43574.4]
  assign regs_424_io_in = 64'h0; // @[RegFile.scala 75:16:@43573.4]
  assign regs_424_io_reset = reset; // @[RegFile.scala 78:19:@43577.4]
  assign regs_424_io_enable = 1'h1; // @[RegFile.scala 74:20:@43571.4]
  assign regs_425_clock = clock; // @[:@43580.4]
  assign regs_425_reset = io_reset; // @[:@43581.4 RegFile.scala 76:16:@43588.4]
  assign regs_425_io_in = 64'h0; // @[RegFile.scala 75:16:@43587.4]
  assign regs_425_io_reset = reset; // @[RegFile.scala 78:19:@43591.4]
  assign regs_425_io_enable = 1'h1; // @[RegFile.scala 74:20:@43585.4]
  assign regs_426_clock = clock; // @[:@43594.4]
  assign regs_426_reset = io_reset; // @[:@43595.4 RegFile.scala 76:16:@43602.4]
  assign regs_426_io_in = 64'h0; // @[RegFile.scala 75:16:@43601.4]
  assign regs_426_io_reset = reset; // @[RegFile.scala 78:19:@43605.4]
  assign regs_426_io_enable = 1'h1; // @[RegFile.scala 74:20:@43599.4]
  assign regs_427_clock = clock; // @[:@43608.4]
  assign regs_427_reset = io_reset; // @[:@43609.4 RegFile.scala 76:16:@43616.4]
  assign regs_427_io_in = 64'h0; // @[RegFile.scala 75:16:@43615.4]
  assign regs_427_io_reset = reset; // @[RegFile.scala 78:19:@43619.4]
  assign regs_427_io_enable = 1'h1; // @[RegFile.scala 74:20:@43613.4]
  assign regs_428_clock = clock; // @[:@43622.4]
  assign regs_428_reset = io_reset; // @[:@43623.4 RegFile.scala 76:16:@43630.4]
  assign regs_428_io_in = 64'h0; // @[RegFile.scala 75:16:@43629.4]
  assign regs_428_io_reset = reset; // @[RegFile.scala 78:19:@43633.4]
  assign regs_428_io_enable = 1'h1; // @[RegFile.scala 74:20:@43627.4]
  assign regs_429_clock = clock; // @[:@43636.4]
  assign regs_429_reset = io_reset; // @[:@43637.4 RegFile.scala 76:16:@43644.4]
  assign regs_429_io_in = 64'h0; // @[RegFile.scala 75:16:@43643.4]
  assign regs_429_io_reset = reset; // @[RegFile.scala 78:19:@43647.4]
  assign regs_429_io_enable = 1'h1; // @[RegFile.scala 74:20:@43641.4]
  assign regs_430_clock = clock; // @[:@43650.4]
  assign regs_430_reset = io_reset; // @[:@43651.4 RegFile.scala 76:16:@43658.4]
  assign regs_430_io_in = 64'h0; // @[RegFile.scala 75:16:@43657.4]
  assign regs_430_io_reset = reset; // @[RegFile.scala 78:19:@43661.4]
  assign regs_430_io_enable = 1'h1; // @[RegFile.scala 74:20:@43655.4]
  assign regs_431_clock = clock; // @[:@43664.4]
  assign regs_431_reset = io_reset; // @[:@43665.4 RegFile.scala 76:16:@43672.4]
  assign regs_431_io_in = 64'h0; // @[RegFile.scala 75:16:@43671.4]
  assign regs_431_io_reset = reset; // @[RegFile.scala 78:19:@43675.4]
  assign regs_431_io_enable = 1'h1; // @[RegFile.scala 74:20:@43669.4]
  assign regs_432_clock = clock; // @[:@43678.4]
  assign regs_432_reset = io_reset; // @[:@43679.4 RegFile.scala 76:16:@43686.4]
  assign regs_432_io_in = 64'h0; // @[RegFile.scala 75:16:@43685.4]
  assign regs_432_io_reset = reset; // @[RegFile.scala 78:19:@43689.4]
  assign regs_432_io_enable = 1'h1; // @[RegFile.scala 74:20:@43683.4]
  assign regs_433_clock = clock; // @[:@43692.4]
  assign regs_433_reset = io_reset; // @[:@43693.4 RegFile.scala 76:16:@43700.4]
  assign regs_433_io_in = 64'h0; // @[RegFile.scala 75:16:@43699.4]
  assign regs_433_io_reset = reset; // @[RegFile.scala 78:19:@43703.4]
  assign regs_433_io_enable = 1'h1; // @[RegFile.scala 74:20:@43697.4]
  assign regs_434_clock = clock; // @[:@43706.4]
  assign regs_434_reset = io_reset; // @[:@43707.4 RegFile.scala 76:16:@43714.4]
  assign regs_434_io_in = 64'h0; // @[RegFile.scala 75:16:@43713.4]
  assign regs_434_io_reset = reset; // @[RegFile.scala 78:19:@43717.4]
  assign regs_434_io_enable = 1'h1; // @[RegFile.scala 74:20:@43711.4]
  assign regs_435_clock = clock; // @[:@43720.4]
  assign regs_435_reset = io_reset; // @[:@43721.4 RegFile.scala 76:16:@43728.4]
  assign regs_435_io_in = 64'h0; // @[RegFile.scala 75:16:@43727.4]
  assign regs_435_io_reset = reset; // @[RegFile.scala 78:19:@43731.4]
  assign regs_435_io_enable = 1'h1; // @[RegFile.scala 74:20:@43725.4]
  assign regs_436_clock = clock; // @[:@43734.4]
  assign regs_436_reset = io_reset; // @[:@43735.4 RegFile.scala 76:16:@43742.4]
  assign regs_436_io_in = 64'h0; // @[RegFile.scala 75:16:@43741.4]
  assign regs_436_io_reset = reset; // @[RegFile.scala 78:19:@43745.4]
  assign regs_436_io_enable = 1'h1; // @[RegFile.scala 74:20:@43739.4]
  assign regs_437_clock = clock; // @[:@43748.4]
  assign regs_437_reset = io_reset; // @[:@43749.4 RegFile.scala 76:16:@43756.4]
  assign regs_437_io_in = 64'h0; // @[RegFile.scala 75:16:@43755.4]
  assign regs_437_io_reset = reset; // @[RegFile.scala 78:19:@43759.4]
  assign regs_437_io_enable = 1'h1; // @[RegFile.scala 74:20:@43753.4]
  assign regs_438_clock = clock; // @[:@43762.4]
  assign regs_438_reset = io_reset; // @[:@43763.4 RegFile.scala 76:16:@43770.4]
  assign regs_438_io_in = 64'h0; // @[RegFile.scala 75:16:@43769.4]
  assign regs_438_io_reset = reset; // @[RegFile.scala 78:19:@43773.4]
  assign regs_438_io_enable = 1'h1; // @[RegFile.scala 74:20:@43767.4]
  assign regs_439_clock = clock; // @[:@43776.4]
  assign regs_439_reset = io_reset; // @[:@43777.4 RegFile.scala 76:16:@43784.4]
  assign regs_439_io_in = 64'h0; // @[RegFile.scala 75:16:@43783.4]
  assign regs_439_io_reset = reset; // @[RegFile.scala 78:19:@43787.4]
  assign regs_439_io_enable = 1'h1; // @[RegFile.scala 74:20:@43781.4]
  assign regs_440_clock = clock; // @[:@43790.4]
  assign regs_440_reset = io_reset; // @[:@43791.4 RegFile.scala 76:16:@43798.4]
  assign regs_440_io_in = 64'h0; // @[RegFile.scala 75:16:@43797.4]
  assign regs_440_io_reset = reset; // @[RegFile.scala 78:19:@43801.4]
  assign regs_440_io_enable = 1'h1; // @[RegFile.scala 74:20:@43795.4]
  assign regs_441_clock = clock; // @[:@43804.4]
  assign regs_441_reset = io_reset; // @[:@43805.4 RegFile.scala 76:16:@43812.4]
  assign regs_441_io_in = 64'h0; // @[RegFile.scala 75:16:@43811.4]
  assign regs_441_io_reset = reset; // @[RegFile.scala 78:19:@43815.4]
  assign regs_441_io_enable = 1'h1; // @[RegFile.scala 74:20:@43809.4]
  assign regs_442_clock = clock; // @[:@43818.4]
  assign regs_442_reset = io_reset; // @[:@43819.4 RegFile.scala 76:16:@43826.4]
  assign regs_442_io_in = 64'h0; // @[RegFile.scala 75:16:@43825.4]
  assign regs_442_io_reset = reset; // @[RegFile.scala 78:19:@43829.4]
  assign regs_442_io_enable = 1'h1; // @[RegFile.scala 74:20:@43823.4]
  assign regs_443_clock = clock; // @[:@43832.4]
  assign regs_443_reset = io_reset; // @[:@43833.4 RegFile.scala 76:16:@43840.4]
  assign regs_443_io_in = 64'h0; // @[RegFile.scala 75:16:@43839.4]
  assign regs_443_io_reset = reset; // @[RegFile.scala 78:19:@43843.4]
  assign regs_443_io_enable = 1'h1; // @[RegFile.scala 74:20:@43837.4]
  assign regs_444_clock = clock; // @[:@43846.4]
  assign regs_444_reset = io_reset; // @[:@43847.4 RegFile.scala 76:16:@43854.4]
  assign regs_444_io_in = 64'h0; // @[RegFile.scala 75:16:@43853.4]
  assign regs_444_io_reset = reset; // @[RegFile.scala 78:19:@43857.4]
  assign regs_444_io_enable = 1'h1; // @[RegFile.scala 74:20:@43851.4]
  assign regs_445_clock = clock; // @[:@43860.4]
  assign regs_445_reset = io_reset; // @[:@43861.4 RegFile.scala 76:16:@43868.4]
  assign regs_445_io_in = 64'h0; // @[RegFile.scala 75:16:@43867.4]
  assign regs_445_io_reset = reset; // @[RegFile.scala 78:19:@43871.4]
  assign regs_445_io_enable = 1'h1; // @[RegFile.scala 74:20:@43865.4]
  assign regs_446_clock = clock; // @[:@43874.4]
  assign regs_446_reset = io_reset; // @[:@43875.4 RegFile.scala 76:16:@43882.4]
  assign regs_446_io_in = 64'h0; // @[RegFile.scala 75:16:@43881.4]
  assign regs_446_io_reset = reset; // @[RegFile.scala 78:19:@43885.4]
  assign regs_446_io_enable = 1'h1; // @[RegFile.scala 74:20:@43879.4]
  assign regs_447_clock = clock; // @[:@43888.4]
  assign regs_447_reset = io_reset; // @[:@43889.4 RegFile.scala 76:16:@43896.4]
  assign regs_447_io_in = 64'h0; // @[RegFile.scala 75:16:@43895.4]
  assign regs_447_io_reset = reset; // @[RegFile.scala 78:19:@43899.4]
  assign regs_447_io_enable = 1'h1; // @[RegFile.scala 74:20:@43893.4]
  assign regs_448_clock = clock; // @[:@43902.4]
  assign regs_448_reset = io_reset; // @[:@43903.4 RegFile.scala 76:16:@43910.4]
  assign regs_448_io_in = 64'h0; // @[RegFile.scala 75:16:@43909.4]
  assign regs_448_io_reset = reset; // @[RegFile.scala 78:19:@43913.4]
  assign regs_448_io_enable = 1'h1; // @[RegFile.scala 74:20:@43907.4]
  assign regs_449_clock = clock; // @[:@43916.4]
  assign regs_449_reset = io_reset; // @[:@43917.4 RegFile.scala 76:16:@43924.4]
  assign regs_449_io_in = 64'h0; // @[RegFile.scala 75:16:@43923.4]
  assign regs_449_io_reset = reset; // @[RegFile.scala 78:19:@43927.4]
  assign regs_449_io_enable = 1'h1; // @[RegFile.scala 74:20:@43921.4]
  assign regs_450_clock = clock; // @[:@43930.4]
  assign regs_450_reset = io_reset; // @[:@43931.4 RegFile.scala 76:16:@43938.4]
  assign regs_450_io_in = 64'h0; // @[RegFile.scala 75:16:@43937.4]
  assign regs_450_io_reset = reset; // @[RegFile.scala 78:19:@43941.4]
  assign regs_450_io_enable = 1'h1; // @[RegFile.scala 74:20:@43935.4]
  assign regs_451_clock = clock; // @[:@43944.4]
  assign regs_451_reset = io_reset; // @[:@43945.4 RegFile.scala 76:16:@43952.4]
  assign regs_451_io_in = 64'h0; // @[RegFile.scala 75:16:@43951.4]
  assign regs_451_io_reset = reset; // @[RegFile.scala 78:19:@43955.4]
  assign regs_451_io_enable = 1'h1; // @[RegFile.scala 74:20:@43949.4]
  assign regs_452_clock = clock; // @[:@43958.4]
  assign regs_452_reset = io_reset; // @[:@43959.4 RegFile.scala 76:16:@43966.4]
  assign regs_452_io_in = 64'h0; // @[RegFile.scala 75:16:@43965.4]
  assign regs_452_io_reset = reset; // @[RegFile.scala 78:19:@43969.4]
  assign regs_452_io_enable = 1'h1; // @[RegFile.scala 74:20:@43963.4]
  assign regs_453_clock = clock; // @[:@43972.4]
  assign regs_453_reset = io_reset; // @[:@43973.4 RegFile.scala 76:16:@43980.4]
  assign regs_453_io_in = 64'h0; // @[RegFile.scala 75:16:@43979.4]
  assign regs_453_io_reset = reset; // @[RegFile.scala 78:19:@43983.4]
  assign regs_453_io_enable = 1'h1; // @[RegFile.scala 74:20:@43977.4]
  assign regs_454_clock = clock; // @[:@43986.4]
  assign regs_454_reset = io_reset; // @[:@43987.4 RegFile.scala 76:16:@43994.4]
  assign regs_454_io_in = 64'h0; // @[RegFile.scala 75:16:@43993.4]
  assign regs_454_io_reset = reset; // @[RegFile.scala 78:19:@43997.4]
  assign regs_454_io_enable = 1'h1; // @[RegFile.scala 74:20:@43991.4]
  assign regs_455_clock = clock; // @[:@44000.4]
  assign regs_455_reset = io_reset; // @[:@44001.4 RegFile.scala 76:16:@44008.4]
  assign regs_455_io_in = 64'h0; // @[RegFile.scala 75:16:@44007.4]
  assign regs_455_io_reset = reset; // @[RegFile.scala 78:19:@44011.4]
  assign regs_455_io_enable = 1'h1; // @[RegFile.scala 74:20:@44005.4]
  assign regs_456_clock = clock; // @[:@44014.4]
  assign regs_456_reset = io_reset; // @[:@44015.4 RegFile.scala 76:16:@44022.4]
  assign regs_456_io_in = 64'h0; // @[RegFile.scala 75:16:@44021.4]
  assign regs_456_io_reset = reset; // @[RegFile.scala 78:19:@44025.4]
  assign regs_456_io_enable = 1'h1; // @[RegFile.scala 74:20:@44019.4]
  assign regs_457_clock = clock; // @[:@44028.4]
  assign regs_457_reset = io_reset; // @[:@44029.4 RegFile.scala 76:16:@44036.4]
  assign regs_457_io_in = 64'h0; // @[RegFile.scala 75:16:@44035.4]
  assign regs_457_io_reset = reset; // @[RegFile.scala 78:19:@44039.4]
  assign regs_457_io_enable = 1'h1; // @[RegFile.scala 74:20:@44033.4]
  assign regs_458_clock = clock; // @[:@44042.4]
  assign regs_458_reset = io_reset; // @[:@44043.4 RegFile.scala 76:16:@44050.4]
  assign regs_458_io_in = 64'h0; // @[RegFile.scala 75:16:@44049.4]
  assign regs_458_io_reset = reset; // @[RegFile.scala 78:19:@44053.4]
  assign regs_458_io_enable = 1'h1; // @[RegFile.scala 74:20:@44047.4]
  assign regs_459_clock = clock; // @[:@44056.4]
  assign regs_459_reset = io_reset; // @[:@44057.4 RegFile.scala 76:16:@44064.4]
  assign regs_459_io_in = 64'h0; // @[RegFile.scala 75:16:@44063.4]
  assign regs_459_io_reset = reset; // @[RegFile.scala 78:19:@44067.4]
  assign regs_459_io_enable = 1'h1; // @[RegFile.scala 74:20:@44061.4]
  assign regs_460_clock = clock; // @[:@44070.4]
  assign regs_460_reset = io_reset; // @[:@44071.4 RegFile.scala 76:16:@44078.4]
  assign regs_460_io_in = 64'h0; // @[RegFile.scala 75:16:@44077.4]
  assign regs_460_io_reset = reset; // @[RegFile.scala 78:19:@44081.4]
  assign regs_460_io_enable = 1'h1; // @[RegFile.scala 74:20:@44075.4]
  assign regs_461_clock = clock; // @[:@44084.4]
  assign regs_461_reset = io_reset; // @[:@44085.4 RegFile.scala 76:16:@44092.4]
  assign regs_461_io_in = 64'h0; // @[RegFile.scala 75:16:@44091.4]
  assign regs_461_io_reset = reset; // @[RegFile.scala 78:19:@44095.4]
  assign regs_461_io_enable = 1'h1; // @[RegFile.scala 74:20:@44089.4]
  assign regs_462_clock = clock; // @[:@44098.4]
  assign regs_462_reset = io_reset; // @[:@44099.4 RegFile.scala 76:16:@44106.4]
  assign regs_462_io_in = 64'h0; // @[RegFile.scala 75:16:@44105.4]
  assign regs_462_io_reset = reset; // @[RegFile.scala 78:19:@44109.4]
  assign regs_462_io_enable = 1'h1; // @[RegFile.scala 74:20:@44103.4]
  assign regs_463_clock = clock; // @[:@44112.4]
  assign regs_463_reset = io_reset; // @[:@44113.4 RegFile.scala 76:16:@44120.4]
  assign regs_463_io_in = 64'h0; // @[RegFile.scala 75:16:@44119.4]
  assign regs_463_io_reset = reset; // @[RegFile.scala 78:19:@44123.4]
  assign regs_463_io_enable = 1'h1; // @[RegFile.scala 74:20:@44117.4]
  assign regs_464_clock = clock; // @[:@44126.4]
  assign regs_464_reset = io_reset; // @[:@44127.4 RegFile.scala 76:16:@44134.4]
  assign regs_464_io_in = 64'h0; // @[RegFile.scala 75:16:@44133.4]
  assign regs_464_io_reset = reset; // @[RegFile.scala 78:19:@44137.4]
  assign regs_464_io_enable = 1'h1; // @[RegFile.scala 74:20:@44131.4]
  assign regs_465_clock = clock; // @[:@44140.4]
  assign regs_465_reset = io_reset; // @[:@44141.4 RegFile.scala 76:16:@44148.4]
  assign regs_465_io_in = 64'h0; // @[RegFile.scala 75:16:@44147.4]
  assign regs_465_io_reset = reset; // @[RegFile.scala 78:19:@44151.4]
  assign regs_465_io_enable = 1'h1; // @[RegFile.scala 74:20:@44145.4]
  assign regs_466_clock = clock; // @[:@44154.4]
  assign regs_466_reset = io_reset; // @[:@44155.4 RegFile.scala 76:16:@44162.4]
  assign regs_466_io_in = 64'h0; // @[RegFile.scala 75:16:@44161.4]
  assign regs_466_io_reset = reset; // @[RegFile.scala 78:19:@44165.4]
  assign regs_466_io_enable = 1'h1; // @[RegFile.scala 74:20:@44159.4]
  assign regs_467_clock = clock; // @[:@44168.4]
  assign regs_467_reset = io_reset; // @[:@44169.4 RegFile.scala 76:16:@44176.4]
  assign regs_467_io_in = 64'h0; // @[RegFile.scala 75:16:@44175.4]
  assign regs_467_io_reset = reset; // @[RegFile.scala 78:19:@44179.4]
  assign regs_467_io_enable = 1'h1; // @[RegFile.scala 74:20:@44173.4]
  assign regs_468_clock = clock; // @[:@44182.4]
  assign regs_468_reset = io_reset; // @[:@44183.4 RegFile.scala 76:16:@44190.4]
  assign regs_468_io_in = 64'h0; // @[RegFile.scala 75:16:@44189.4]
  assign regs_468_io_reset = reset; // @[RegFile.scala 78:19:@44193.4]
  assign regs_468_io_enable = 1'h1; // @[RegFile.scala 74:20:@44187.4]
  assign regs_469_clock = clock; // @[:@44196.4]
  assign regs_469_reset = io_reset; // @[:@44197.4 RegFile.scala 76:16:@44204.4]
  assign regs_469_io_in = 64'h0; // @[RegFile.scala 75:16:@44203.4]
  assign regs_469_io_reset = reset; // @[RegFile.scala 78:19:@44207.4]
  assign regs_469_io_enable = 1'h1; // @[RegFile.scala 74:20:@44201.4]
  assign regs_470_clock = clock; // @[:@44210.4]
  assign regs_470_reset = io_reset; // @[:@44211.4 RegFile.scala 76:16:@44218.4]
  assign regs_470_io_in = 64'h0; // @[RegFile.scala 75:16:@44217.4]
  assign regs_470_io_reset = reset; // @[RegFile.scala 78:19:@44221.4]
  assign regs_470_io_enable = 1'h1; // @[RegFile.scala 74:20:@44215.4]
  assign regs_471_clock = clock; // @[:@44224.4]
  assign regs_471_reset = io_reset; // @[:@44225.4 RegFile.scala 76:16:@44232.4]
  assign regs_471_io_in = 64'h0; // @[RegFile.scala 75:16:@44231.4]
  assign regs_471_io_reset = reset; // @[RegFile.scala 78:19:@44235.4]
  assign regs_471_io_enable = 1'h1; // @[RegFile.scala 74:20:@44229.4]
  assign regs_472_clock = clock; // @[:@44238.4]
  assign regs_472_reset = io_reset; // @[:@44239.4 RegFile.scala 76:16:@44246.4]
  assign regs_472_io_in = 64'h0; // @[RegFile.scala 75:16:@44245.4]
  assign regs_472_io_reset = reset; // @[RegFile.scala 78:19:@44249.4]
  assign regs_472_io_enable = 1'h1; // @[RegFile.scala 74:20:@44243.4]
  assign regs_473_clock = clock; // @[:@44252.4]
  assign regs_473_reset = io_reset; // @[:@44253.4 RegFile.scala 76:16:@44260.4]
  assign regs_473_io_in = 64'h0; // @[RegFile.scala 75:16:@44259.4]
  assign regs_473_io_reset = reset; // @[RegFile.scala 78:19:@44263.4]
  assign regs_473_io_enable = 1'h1; // @[RegFile.scala 74:20:@44257.4]
  assign regs_474_clock = clock; // @[:@44266.4]
  assign regs_474_reset = io_reset; // @[:@44267.4 RegFile.scala 76:16:@44274.4]
  assign regs_474_io_in = 64'h0; // @[RegFile.scala 75:16:@44273.4]
  assign regs_474_io_reset = reset; // @[RegFile.scala 78:19:@44277.4]
  assign regs_474_io_enable = 1'h1; // @[RegFile.scala 74:20:@44271.4]
  assign regs_475_clock = clock; // @[:@44280.4]
  assign regs_475_reset = io_reset; // @[:@44281.4 RegFile.scala 76:16:@44288.4]
  assign regs_475_io_in = 64'h0; // @[RegFile.scala 75:16:@44287.4]
  assign regs_475_io_reset = reset; // @[RegFile.scala 78:19:@44291.4]
  assign regs_475_io_enable = 1'h1; // @[RegFile.scala 74:20:@44285.4]
  assign regs_476_clock = clock; // @[:@44294.4]
  assign regs_476_reset = io_reset; // @[:@44295.4 RegFile.scala 76:16:@44302.4]
  assign regs_476_io_in = 64'h0; // @[RegFile.scala 75:16:@44301.4]
  assign regs_476_io_reset = reset; // @[RegFile.scala 78:19:@44305.4]
  assign regs_476_io_enable = 1'h1; // @[RegFile.scala 74:20:@44299.4]
  assign regs_477_clock = clock; // @[:@44308.4]
  assign regs_477_reset = io_reset; // @[:@44309.4 RegFile.scala 76:16:@44316.4]
  assign regs_477_io_in = 64'h0; // @[RegFile.scala 75:16:@44315.4]
  assign regs_477_io_reset = reset; // @[RegFile.scala 78:19:@44319.4]
  assign regs_477_io_enable = 1'h1; // @[RegFile.scala 74:20:@44313.4]
  assign regs_478_clock = clock; // @[:@44322.4]
  assign regs_478_reset = io_reset; // @[:@44323.4 RegFile.scala 76:16:@44330.4]
  assign regs_478_io_in = 64'h0; // @[RegFile.scala 75:16:@44329.4]
  assign regs_478_io_reset = reset; // @[RegFile.scala 78:19:@44333.4]
  assign regs_478_io_enable = 1'h1; // @[RegFile.scala 74:20:@44327.4]
  assign regs_479_clock = clock; // @[:@44336.4]
  assign regs_479_reset = io_reset; // @[:@44337.4 RegFile.scala 76:16:@44344.4]
  assign regs_479_io_in = 64'h0; // @[RegFile.scala 75:16:@44343.4]
  assign regs_479_io_reset = reset; // @[RegFile.scala 78:19:@44347.4]
  assign regs_479_io_enable = 1'h1; // @[RegFile.scala 74:20:@44341.4]
  assign regs_480_clock = clock; // @[:@44350.4]
  assign regs_480_reset = io_reset; // @[:@44351.4 RegFile.scala 76:16:@44358.4]
  assign regs_480_io_in = 64'h0; // @[RegFile.scala 75:16:@44357.4]
  assign regs_480_io_reset = reset; // @[RegFile.scala 78:19:@44361.4]
  assign regs_480_io_enable = 1'h1; // @[RegFile.scala 74:20:@44355.4]
  assign regs_481_clock = clock; // @[:@44364.4]
  assign regs_481_reset = io_reset; // @[:@44365.4 RegFile.scala 76:16:@44372.4]
  assign regs_481_io_in = 64'h0; // @[RegFile.scala 75:16:@44371.4]
  assign regs_481_io_reset = reset; // @[RegFile.scala 78:19:@44375.4]
  assign regs_481_io_enable = 1'h1; // @[RegFile.scala 74:20:@44369.4]
  assign regs_482_clock = clock; // @[:@44378.4]
  assign regs_482_reset = io_reset; // @[:@44379.4 RegFile.scala 76:16:@44386.4]
  assign regs_482_io_in = 64'h0; // @[RegFile.scala 75:16:@44385.4]
  assign regs_482_io_reset = reset; // @[RegFile.scala 78:19:@44389.4]
  assign regs_482_io_enable = 1'h1; // @[RegFile.scala 74:20:@44383.4]
  assign regs_483_clock = clock; // @[:@44392.4]
  assign regs_483_reset = io_reset; // @[:@44393.4 RegFile.scala 76:16:@44400.4]
  assign regs_483_io_in = 64'h0; // @[RegFile.scala 75:16:@44399.4]
  assign regs_483_io_reset = reset; // @[RegFile.scala 78:19:@44403.4]
  assign regs_483_io_enable = 1'h1; // @[RegFile.scala 74:20:@44397.4]
  assign regs_484_clock = clock; // @[:@44406.4]
  assign regs_484_reset = io_reset; // @[:@44407.4 RegFile.scala 76:16:@44414.4]
  assign regs_484_io_in = 64'h0; // @[RegFile.scala 75:16:@44413.4]
  assign regs_484_io_reset = reset; // @[RegFile.scala 78:19:@44417.4]
  assign regs_484_io_enable = 1'h1; // @[RegFile.scala 74:20:@44411.4]
  assign regs_485_clock = clock; // @[:@44420.4]
  assign regs_485_reset = io_reset; // @[:@44421.4 RegFile.scala 76:16:@44428.4]
  assign regs_485_io_in = 64'h0; // @[RegFile.scala 75:16:@44427.4]
  assign regs_485_io_reset = reset; // @[RegFile.scala 78:19:@44431.4]
  assign regs_485_io_enable = 1'h1; // @[RegFile.scala 74:20:@44425.4]
  assign regs_486_clock = clock; // @[:@44434.4]
  assign regs_486_reset = io_reset; // @[:@44435.4 RegFile.scala 76:16:@44442.4]
  assign regs_486_io_in = 64'h0; // @[RegFile.scala 75:16:@44441.4]
  assign regs_486_io_reset = reset; // @[RegFile.scala 78:19:@44445.4]
  assign regs_486_io_enable = 1'h1; // @[RegFile.scala 74:20:@44439.4]
  assign regs_487_clock = clock; // @[:@44448.4]
  assign regs_487_reset = io_reset; // @[:@44449.4 RegFile.scala 76:16:@44456.4]
  assign regs_487_io_in = 64'h0; // @[RegFile.scala 75:16:@44455.4]
  assign regs_487_io_reset = reset; // @[RegFile.scala 78:19:@44459.4]
  assign regs_487_io_enable = 1'h1; // @[RegFile.scala 74:20:@44453.4]
  assign regs_488_clock = clock; // @[:@44462.4]
  assign regs_488_reset = io_reset; // @[:@44463.4 RegFile.scala 76:16:@44470.4]
  assign regs_488_io_in = 64'h0; // @[RegFile.scala 75:16:@44469.4]
  assign regs_488_io_reset = reset; // @[RegFile.scala 78:19:@44473.4]
  assign regs_488_io_enable = 1'h1; // @[RegFile.scala 74:20:@44467.4]
  assign regs_489_clock = clock; // @[:@44476.4]
  assign regs_489_reset = io_reset; // @[:@44477.4 RegFile.scala 76:16:@44484.4]
  assign regs_489_io_in = 64'h0; // @[RegFile.scala 75:16:@44483.4]
  assign regs_489_io_reset = reset; // @[RegFile.scala 78:19:@44487.4]
  assign regs_489_io_enable = 1'h1; // @[RegFile.scala 74:20:@44481.4]
  assign regs_490_clock = clock; // @[:@44490.4]
  assign regs_490_reset = io_reset; // @[:@44491.4 RegFile.scala 76:16:@44498.4]
  assign regs_490_io_in = 64'h0; // @[RegFile.scala 75:16:@44497.4]
  assign regs_490_io_reset = reset; // @[RegFile.scala 78:19:@44501.4]
  assign regs_490_io_enable = 1'h1; // @[RegFile.scala 74:20:@44495.4]
  assign regs_491_clock = clock; // @[:@44504.4]
  assign regs_491_reset = io_reset; // @[:@44505.4 RegFile.scala 76:16:@44512.4]
  assign regs_491_io_in = 64'h0; // @[RegFile.scala 75:16:@44511.4]
  assign regs_491_io_reset = reset; // @[RegFile.scala 78:19:@44515.4]
  assign regs_491_io_enable = 1'h1; // @[RegFile.scala 74:20:@44509.4]
  assign regs_492_clock = clock; // @[:@44518.4]
  assign regs_492_reset = io_reset; // @[:@44519.4 RegFile.scala 76:16:@44526.4]
  assign regs_492_io_in = 64'h0; // @[RegFile.scala 75:16:@44525.4]
  assign regs_492_io_reset = reset; // @[RegFile.scala 78:19:@44529.4]
  assign regs_492_io_enable = 1'h1; // @[RegFile.scala 74:20:@44523.4]
  assign regs_493_clock = clock; // @[:@44532.4]
  assign regs_493_reset = io_reset; // @[:@44533.4 RegFile.scala 76:16:@44540.4]
  assign regs_493_io_in = 64'h0; // @[RegFile.scala 75:16:@44539.4]
  assign regs_493_io_reset = reset; // @[RegFile.scala 78:19:@44543.4]
  assign regs_493_io_enable = 1'h1; // @[RegFile.scala 74:20:@44537.4]
  assign regs_494_clock = clock; // @[:@44546.4]
  assign regs_494_reset = io_reset; // @[:@44547.4 RegFile.scala 76:16:@44554.4]
  assign regs_494_io_in = 64'h0; // @[RegFile.scala 75:16:@44553.4]
  assign regs_494_io_reset = reset; // @[RegFile.scala 78:19:@44557.4]
  assign regs_494_io_enable = 1'h1; // @[RegFile.scala 74:20:@44551.4]
  assign regs_495_clock = clock; // @[:@44560.4]
  assign regs_495_reset = io_reset; // @[:@44561.4 RegFile.scala 76:16:@44568.4]
  assign regs_495_io_in = 64'h0; // @[RegFile.scala 75:16:@44567.4]
  assign regs_495_io_reset = reset; // @[RegFile.scala 78:19:@44571.4]
  assign regs_495_io_enable = 1'h1; // @[RegFile.scala 74:20:@44565.4]
  assign regs_496_clock = clock; // @[:@44574.4]
  assign regs_496_reset = io_reset; // @[:@44575.4 RegFile.scala 76:16:@44582.4]
  assign regs_496_io_in = 64'h0; // @[RegFile.scala 75:16:@44581.4]
  assign regs_496_io_reset = reset; // @[RegFile.scala 78:19:@44585.4]
  assign regs_496_io_enable = 1'h1; // @[RegFile.scala 74:20:@44579.4]
  assign regs_497_clock = clock; // @[:@44588.4]
  assign regs_497_reset = io_reset; // @[:@44589.4 RegFile.scala 76:16:@44596.4]
  assign regs_497_io_in = 64'h0; // @[RegFile.scala 75:16:@44595.4]
  assign regs_497_io_reset = reset; // @[RegFile.scala 78:19:@44599.4]
  assign regs_497_io_enable = 1'h1; // @[RegFile.scala 74:20:@44593.4]
  assign regs_498_clock = clock; // @[:@44602.4]
  assign regs_498_reset = io_reset; // @[:@44603.4 RegFile.scala 76:16:@44610.4]
  assign regs_498_io_in = 64'h0; // @[RegFile.scala 75:16:@44609.4]
  assign regs_498_io_reset = reset; // @[RegFile.scala 78:19:@44613.4]
  assign regs_498_io_enable = 1'h1; // @[RegFile.scala 74:20:@44607.4]
  assign regs_499_clock = clock; // @[:@44616.4]
  assign regs_499_reset = io_reset; // @[:@44617.4 RegFile.scala 76:16:@44624.4]
  assign regs_499_io_in = 64'h0; // @[RegFile.scala 75:16:@44623.4]
  assign regs_499_io_reset = reset; // @[RegFile.scala 78:19:@44627.4]
  assign regs_499_io_enable = 1'h1; // @[RegFile.scala 74:20:@44621.4]
  assign regs_500_clock = clock; // @[:@44630.4]
  assign regs_500_reset = io_reset; // @[:@44631.4 RegFile.scala 76:16:@44638.4]
  assign regs_500_io_in = 64'h0; // @[RegFile.scala 75:16:@44637.4]
  assign regs_500_io_reset = reset; // @[RegFile.scala 78:19:@44641.4]
  assign regs_500_io_enable = 1'h1; // @[RegFile.scala 74:20:@44635.4]
  assign regs_501_clock = clock; // @[:@44644.4]
  assign regs_501_reset = io_reset; // @[:@44645.4 RegFile.scala 76:16:@44652.4]
  assign regs_501_io_in = 64'h0; // @[RegFile.scala 75:16:@44651.4]
  assign regs_501_io_reset = reset; // @[RegFile.scala 78:19:@44655.4]
  assign regs_501_io_enable = 1'h1; // @[RegFile.scala 74:20:@44649.4]
  assign regs_502_clock = clock; // @[:@44658.4]
  assign regs_502_reset = io_reset; // @[:@44659.4 RegFile.scala 76:16:@44666.4]
  assign regs_502_io_in = 64'h0; // @[RegFile.scala 75:16:@44665.4]
  assign regs_502_io_reset = reset; // @[RegFile.scala 78:19:@44669.4]
  assign regs_502_io_enable = 1'h1; // @[RegFile.scala 74:20:@44663.4]
  assign regs_503_clock = clock; // @[:@44672.4]
  assign regs_503_reset = io_reset; // @[:@44673.4 RegFile.scala 76:16:@44680.4]
  assign regs_503_io_in = 64'h0; // @[RegFile.scala 75:16:@44679.4]
  assign regs_503_io_reset = reset; // @[RegFile.scala 78:19:@44683.4]
  assign regs_503_io_enable = 1'h1; // @[RegFile.scala 74:20:@44677.4]
  assign regs_504_clock = clock; // @[:@44686.4]
  assign regs_504_reset = io_reset; // @[:@44687.4 RegFile.scala 76:16:@44694.4]
  assign regs_504_io_in = 64'h0; // @[RegFile.scala 75:16:@44693.4]
  assign regs_504_io_reset = reset; // @[RegFile.scala 78:19:@44697.4]
  assign regs_504_io_enable = 1'h1; // @[RegFile.scala 74:20:@44691.4]
  assign regs_505_clock = clock; // @[:@44700.4]
  assign regs_505_reset = io_reset; // @[:@44701.4 RegFile.scala 76:16:@44708.4]
  assign regs_505_io_in = 64'h0; // @[RegFile.scala 75:16:@44707.4]
  assign regs_505_io_reset = reset; // @[RegFile.scala 78:19:@44711.4]
  assign regs_505_io_enable = 1'h1; // @[RegFile.scala 74:20:@44705.4]
  assign regs_506_clock = clock; // @[:@44714.4]
  assign regs_506_reset = io_reset; // @[:@44715.4 RegFile.scala 76:16:@44722.4]
  assign regs_506_io_in = 64'h0; // @[RegFile.scala 75:16:@44721.4]
  assign regs_506_io_reset = reset; // @[RegFile.scala 78:19:@44725.4]
  assign regs_506_io_enable = 1'h1; // @[RegFile.scala 74:20:@44719.4]
  assign regs_507_clock = clock; // @[:@44728.4]
  assign regs_507_reset = io_reset; // @[:@44729.4 RegFile.scala 76:16:@44736.4]
  assign regs_507_io_in = 64'h0; // @[RegFile.scala 75:16:@44735.4]
  assign regs_507_io_reset = reset; // @[RegFile.scala 78:19:@44739.4]
  assign regs_507_io_enable = 1'h1; // @[RegFile.scala 74:20:@44733.4]
  assign regs_508_clock = clock; // @[:@44742.4]
  assign regs_508_reset = io_reset; // @[:@44743.4 RegFile.scala 76:16:@44750.4]
  assign regs_508_io_in = 64'h0; // @[RegFile.scala 75:16:@44749.4]
  assign regs_508_io_reset = reset; // @[RegFile.scala 78:19:@44753.4]
  assign regs_508_io_enable = 1'h1; // @[RegFile.scala 74:20:@44747.4]
  assign regs_509_clock = clock; // @[:@44756.4]
  assign regs_509_reset = io_reset; // @[:@44757.4 RegFile.scala 76:16:@44764.4]
  assign regs_509_io_in = 64'h0; // @[RegFile.scala 75:16:@44763.4]
  assign regs_509_io_reset = reset; // @[RegFile.scala 78:19:@44767.4]
  assign regs_509_io_enable = 1'h1; // @[RegFile.scala 74:20:@44761.4]
  assign regs_510_clock = clock; // @[:@44770.4]
  assign regs_510_reset = io_reset; // @[:@44771.4 RegFile.scala 76:16:@44778.4]
  assign regs_510_io_in = 64'h0; // @[RegFile.scala 75:16:@44777.4]
  assign regs_510_io_reset = reset; // @[RegFile.scala 78:19:@44781.4]
  assign regs_510_io_enable = 1'h1; // @[RegFile.scala 74:20:@44775.4]
  assign regs_511_clock = clock; // @[:@44784.4]
  assign regs_511_reset = io_reset; // @[:@44785.4 RegFile.scala 76:16:@44792.4]
  assign regs_511_io_in = 64'h0; // @[RegFile.scala 75:16:@44791.4]
  assign regs_511_io_reset = reset; // @[RegFile.scala 78:19:@44795.4]
  assign regs_511_io_enable = 1'h1; // @[RegFile.scala 74:20:@44789.4]
  assign rport_io_ins_0 = regs_0_io_out; // @[RegFile.scala 97:16:@45313.4]
  assign rport_io_ins_1 = regs_1_io_out; // @[RegFile.scala 97:16:@45314.4]
  assign rport_io_ins_2 = regs_2_io_out; // @[RegFile.scala 97:16:@45315.4]
  assign rport_io_ins_3 = regs_3_io_out; // @[RegFile.scala 97:16:@45316.4]
  assign rport_io_ins_4 = regs_4_io_out; // @[RegFile.scala 97:16:@45317.4]
  assign rport_io_ins_5 = regs_5_io_out; // @[RegFile.scala 97:16:@45318.4]
  assign rport_io_ins_6 = regs_6_io_out; // @[RegFile.scala 97:16:@45319.4]
  assign rport_io_ins_7 = regs_7_io_out; // @[RegFile.scala 97:16:@45320.4]
  assign rport_io_ins_8 = regs_8_io_out; // @[RegFile.scala 97:16:@45321.4]
  assign rport_io_ins_9 = regs_9_io_out; // @[RegFile.scala 97:16:@45322.4]
  assign rport_io_ins_10 = regs_10_io_out; // @[RegFile.scala 97:16:@45323.4]
  assign rport_io_ins_11 = regs_11_io_out; // @[RegFile.scala 97:16:@45324.4]
  assign rport_io_ins_12 = regs_12_io_out; // @[RegFile.scala 97:16:@45325.4]
  assign rport_io_ins_13 = regs_13_io_out; // @[RegFile.scala 97:16:@45326.4]
  assign rport_io_ins_14 = regs_14_io_out; // @[RegFile.scala 97:16:@45327.4]
  assign rport_io_ins_15 = regs_15_io_out; // @[RegFile.scala 97:16:@45328.4]
  assign rport_io_ins_16 = regs_16_io_out; // @[RegFile.scala 97:16:@45329.4]
  assign rport_io_ins_17 = regs_17_io_out; // @[RegFile.scala 97:16:@45330.4]
  assign rport_io_ins_18 = regs_18_io_out; // @[RegFile.scala 97:16:@45331.4]
  assign rport_io_ins_19 = regs_19_io_out; // @[RegFile.scala 97:16:@45332.4]
  assign rport_io_ins_20 = regs_20_io_out; // @[RegFile.scala 97:16:@45333.4]
  assign rport_io_ins_21 = regs_21_io_out; // @[RegFile.scala 97:16:@45334.4]
  assign rport_io_ins_22 = regs_22_io_out; // @[RegFile.scala 97:16:@45335.4]
  assign rport_io_ins_23 = regs_23_io_out; // @[RegFile.scala 97:16:@45336.4]
  assign rport_io_ins_24 = regs_24_io_out; // @[RegFile.scala 97:16:@45337.4]
  assign rport_io_ins_25 = regs_25_io_out; // @[RegFile.scala 97:16:@45338.4]
  assign rport_io_ins_26 = regs_26_io_out; // @[RegFile.scala 97:16:@45339.4]
  assign rport_io_ins_27 = regs_27_io_out; // @[RegFile.scala 97:16:@45340.4]
  assign rport_io_ins_28 = regs_28_io_out; // @[RegFile.scala 97:16:@45341.4]
  assign rport_io_ins_29 = regs_29_io_out; // @[RegFile.scala 97:16:@45342.4]
  assign rport_io_ins_30 = regs_30_io_out; // @[RegFile.scala 97:16:@45343.4]
  assign rport_io_ins_31 = regs_31_io_out; // @[RegFile.scala 97:16:@45344.4]
  assign rport_io_ins_32 = regs_32_io_out; // @[RegFile.scala 97:16:@45345.4]
  assign rport_io_ins_33 = regs_33_io_out; // @[RegFile.scala 97:16:@45346.4]
  assign rport_io_ins_34 = regs_34_io_out; // @[RegFile.scala 97:16:@45347.4]
  assign rport_io_ins_35 = regs_35_io_out; // @[RegFile.scala 97:16:@45348.4]
  assign rport_io_ins_36 = regs_36_io_out; // @[RegFile.scala 97:16:@45349.4]
  assign rport_io_ins_37 = regs_37_io_out; // @[RegFile.scala 97:16:@45350.4]
  assign rport_io_ins_38 = regs_38_io_out; // @[RegFile.scala 97:16:@45351.4]
  assign rport_io_ins_39 = regs_39_io_out; // @[RegFile.scala 97:16:@45352.4]
  assign rport_io_ins_40 = regs_40_io_out; // @[RegFile.scala 97:16:@45353.4]
  assign rport_io_ins_41 = regs_41_io_out; // @[RegFile.scala 97:16:@45354.4]
  assign rport_io_ins_42 = regs_42_io_out; // @[RegFile.scala 97:16:@45355.4]
  assign rport_io_ins_43 = regs_43_io_out; // @[RegFile.scala 97:16:@45356.4]
  assign rport_io_ins_44 = regs_44_io_out; // @[RegFile.scala 97:16:@45357.4]
  assign rport_io_ins_45 = regs_45_io_out; // @[RegFile.scala 97:16:@45358.4]
  assign rport_io_ins_46 = regs_46_io_out; // @[RegFile.scala 97:16:@45359.4]
  assign rport_io_ins_47 = regs_47_io_out; // @[RegFile.scala 97:16:@45360.4]
  assign rport_io_ins_48 = regs_48_io_out; // @[RegFile.scala 97:16:@45361.4]
  assign rport_io_ins_49 = regs_49_io_out; // @[RegFile.scala 97:16:@45362.4]
  assign rport_io_ins_50 = regs_50_io_out; // @[RegFile.scala 97:16:@45363.4]
  assign rport_io_ins_51 = regs_51_io_out; // @[RegFile.scala 97:16:@45364.4]
  assign rport_io_ins_52 = regs_52_io_out; // @[RegFile.scala 97:16:@45365.4]
  assign rport_io_ins_53 = regs_53_io_out; // @[RegFile.scala 97:16:@45366.4]
  assign rport_io_ins_54 = regs_54_io_out; // @[RegFile.scala 97:16:@45367.4]
  assign rport_io_ins_55 = regs_55_io_out; // @[RegFile.scala 97:16:@45368.4]
  assign rport_io_ins_56 = regs_56_io_out; // @[RegFile.scala 97:16:@45369.4]
  assign rport_io_ins_57 = regs_57_io_out; // @[RegFile.scala 97:16:@45370.4]
  assign rport_io_ins_58 = regs_58_io_out; // @[RegFile.scala 97:16:@45371.4]
  assign rport_io_ins_59 = regs_59_io_out; // @[RegFile.scala 97:16:@45372.4]
  assign rport_io_ins_60 = regs_60_io_out; // @[RegFile.scala 97:16:@45373.4]
  assign rport_io_ins_61 = regs_61_io_out; // @[RegFile.scala 97:16:@45374.4]
  assign rport_io_ins_62 = regs_62_io_out; // @[RegFile.scala 97:16:@45375.4]
  assign rport_io_ins_63 = regs_63_io_out; // @[RegFile.scala 97:16:@45376.4]
  assign rport_io_ins_64 = regs_64_io_out; // @[RegFile.scala 97:16:@45377.4]
  assign rport_io_ins_65 = regs_65_io_out; // @[RegFile.scala 97:16:@45378.4]
  assign rport_io_ins_66 = regs_66_io_out; // @[RegFile.scala 97:16:@45379.4]
  assign rport_io_ins_67 = regs_67_io_out; // @[RegFile.scala 97:16:@45380.4]
  assign rport_io_ins_68 = regs_68_io_out; // @[RegFile.scala 97:16:@45381.4]
  assign rport_io_ins_69 = regs_69_io_out; // @[RegFile.scala 97:16:@45382.4]
  assign rport_io_ins_70 = regs_70_io_out; // @[RegFile.scala 97:16:@45383.4]
  assign rport_io_ins_71 = regs_71_io_out; // @[RegFile.scala 97:16:@45384.4]
  assign rport_io_ins_72 = regs_72_io_out; // @[RegFile.scala 97:16:@45385.4]
  assign rport_io_ins_73 = regs_73_io_out; // @[RegFile.scala 97:16:@45386.4]
  assign rport_io_ins_74 = regs_74_io_out; // @[RegFile.scala 97:16:@45387.4]
  assign rport_io_ins_75 = regs_75_io_out; // @[RegFile.scala 97:16:@45388.4]
  assign rport_io_ins_76 = regs_76_io_out; // @[RegFile.scala 97:16:@45389.4]
  assign rport_io_ins_77 = regs_77_io_out; // @[RegFile.scala 97:16:@45390.4]
  assign rport_io_ins_78 = regs_78_io_out; // @[RegFile.scala 97:16:@45391.4]
  assign rport_io_ins_79 = regs_79_io_out; // @[RegFile.scala 97:16:@45392.4]
  assign rport_io_ins_80 = regs_80_io_out; // @[RegFile.scala 97:16:@45393.4]
  assign rport_io_ins_81 = regs_81_io_out; // @[RegFile.scala 97:16:@45394.4]
  assign rport_io_ins_82 = regs_82_io_out; // @[RegFile.scala 97:16:@45395.4]
  assign rport_io_ins_83 = regs_83_io_out; // @[RegFile.scala 97:16:@45396.4]
  assign rport_io_ins_84 = regs_84_io_out; // @[RegFile.scala 97:16:@45397.4]
  assign rport_io_ins_85 = regs_85_io_out; // @[RegFile.scala 97:16:@45398.4]
  assign rport_io_ins_86 = regs_86_io_out; // @[RegFile.scala 97:16:@45399.4]
  assign rport_io_ins_87 = regs_87_io_out; // @[RegFile.scala 97:16:@45400.4]
  assign rport_io_ins_88 = regs_88_io_out; // @[RegFile.scala 97:16:@45401.4]
  assign rport_io_ins_89 = regs_89_io_out; // @[RegFile.scala 97:16:@45402.4]
  assign rport_io_ins_90 = regs_90_io_out; // @[RegFile.scala 97:16:@45403.4]
  assign rport_io_ins_91 = regs_91_io_out; // @[RegFile.scala 97:16:@45404.4]
  assign rport_io_ins_92 = regs_92_io_out; // @[RegFile.scala 97:16:@45405.4]
  assign rport_io_ins_93 = regs_93_io_out; // @[RegFile.scala 97:16:@45406.4]
  assign rport_io_ins_94 = regs_94_io_out; // @[RegFile.scala 97:16:@45407.4]
  assign rport_io_ins_95 = regs_95_io_out; // @[RegFile.scala 97:16:@45408.4]
  assign rport_io_ins_96 = regs_96_io_out; // @[RegFile.scala 97:16:@45409.4]
  assign rport_io_ins_97 = regs_97_io_out; // @[RegFile.scala 97:16:@45410.4]
  assign rport_io_ins_98 = regs_98_io_out; // @[RegFile.scala 97:16:@45411.4]
  assign rport_io_ins_99 = regs_99_io_out; // @[RegFile.scala 97:16:@45412.4]
  assign rport_io_ins_100 = regs_100_io_out; // @[RegFile.scala 97:16:@45413.4]
  assign rport_io_ins_101 = regs_101_io_out; // @[RegFile.scala 97:16:@45414.4]
  assign rport_io_ins_102 = regs_102_io_out; // @[RegFile.scala 97:16:@45415.4]
  assign rport_io_ins_103 = regs_103_io_out; // @[RegFile.scala 97:16:@45416.4]
  assign rport_io_ins_104 = regs_104_io_out; // @[RegFile.scala 97:16:@45417.4]
  assign rport_io_ins_105 = regs_105_io_out; // @[RegFile.scala 97:16:@45418.4]
  assign rport_io_ins_106 = regs_106_io_out; // @[RegFile.scala 97:16:@45419.4]
  assign rport_io_ins_107 = regs_107_io_out; // @[RegFile.scala 97:16:@45420.4]
  assign rport_io_ins_108 = regs_108_io_out; // @[RegFile.scala 97:16:@45421.4]
  assign rport_io_ins_109 = regs_109_io_out; // @[RegFile.scala 97:16:@45422.4]
  assign rport_io_ins_110 = regs_110_io_out; // @[RegFile.scala 97:16:@45423.4]
  assign rport_io_ins_111 = regs_111_io_out; // @[RegFile.scala 97:16:@45424.4]
  assign rport_io_ins_112 = regs_112_io_out; // @[RegFile.scala 97:16:@45425.4]
  assign rport_io_ins_113 = regs_113_io_out; // @[RegFile.scala 97:16:@45426.4]
  assign rport_io_ins_114 = regs_114_io_out; // @[RegFile.scala 97:16:@45427.4]
  assign rport_io_ins_115 = regs_115_io_out; // @[RegFile.scala 97:16:@45428.4]
  assign rport_io_ins_116 = regs_116_io_out; // @[RegFile.scala 97:16:@45429.4]
  assign rport_io_ins_117 = regs_117_io_out; // @[RegFile.scala 97:16:@45430.4]
  assign rport_io_ins_118 = regs_118_io_out; // @[RegFile.scala 97:16:@45431.4]
  assign rport_io_ins_119 = regs_119_io_out; // @[RegFile.scala 97:16:@45432.4]
  assign rport_io_ins_120 = regs_120_io_out; // @[RegFile.scala 97:16:@45433.4]
  assign rport_io_ins_121 = regs_121_io_out; // @[RegFile.scala 97:16:@45434.4]
  assign rport_io_ins_122 = regs_122_io_out; // @[RegFile.scala 97:16:@45435.4]
  assign rport_io_ins_123 = regs_123_io_out; // @[RegFile.scala 97:16:@45436.4]
  assign rport_io_ins_124 = regs_124_io_out; // @[RegFile.scala 97:16:@45437.4]
  assign rport_io_ins_125 = regs_125_io_out; // @[RegFile.scala 97:16:@45438.4]
  assign rport_io_ins_126 = regs_126_io_out; // @[RegFile.scala 97:16:@45439.4]
  assign rport_io_ins_127 = regs_127_io_out; // @[RegFile.scala 97:16:@45440.4]
  assign rport_io_ins_128 = regs_128_io_out; // @[RegFile.scala 97:16:@45441.4]
  assign rport_io_ins_129 = regs_129_io_out; // @[RegFile.scala 97:16:@45442.4]
  assign rport_io_ins_130 = regs_130_io_out; // @[RegFile.scala 97:16:@45443.4]
  assign rport_io_ins_131 = regs_131_io_out; // @[RegFile.scala 97:16:@45444.4]
  assign rport_io_ins_132 = regs_132_io_out; // @[RegFile.scala 97:16:@45445.4]
  assign rport_io_ins_133 = regs_133_io_out; // @[RegFile.scala 97:16:@45446.4]
  assign rport_io_ins_134 = regs_134_io_out; // @[RegFile.scala 97:16:@45447.4]
  assign rport_io_ins_135 = regs_135_io_out; // @[RegFile.scala 97:16:@45448.4]
  assign rport_io_ins_136 = regs_136_io_out; // @[RegFile.scala 97:16:@45449.4]
  assign rport_io_ins_137 = regs_137_io_out; // @[RegFile.scala 97:16:@45450.4]
  assign rport_io_ins_138 = regs_138_io_out; // @[RegFile.scala 97:16:@45451.4]
  assign rport_io_ins_139 = regs_139_io_out; // @[RegFile.scala 97:16:@45452.4]
  assign rport_io_ins_140 = regs_140_io_out; // @[RegFile.scala 97:16:@45453.4]
  assign rport_io_ins_141 = regs_141_io_out; // @[RegFile.scala 97:16:@45454.4]
  assign rport_io_ins_142 = regs_142_io_out; // @[RegFile.scala 97:16:@45455.4]
  assign rport_io_ins_143 = regs_143_io_out; // @[RegFile.scala 97:16:@45456.4]
  assign rport_io_ins_144 = regs_144_io_out; // @[RegFile.scala 97:16:@45457.4]
  assign rport_io_ins_145 = regs_145_io_out; // @[RegFile.scala 97:16:@45458.4]
  assign rport_io_ins_146 = regs_146_io_out; // @[RegFile.scala 97:16:@45459.4]
  assign rport_io_ins_147 = regs_147_io_out; // @[RegFile.scala 97:16:@45460.4]
  assign rport_io_ins_148 = regs_148_io_out; // @[RegFile.scala 97:16:@45461.4]
  assign rport_io_ins_149 = regs_149_io_out; // @[RegFile.scala 97:16:@45462.4]
  assign rport_io_ins_150 = regs_150_io_out; // @[RegFile.scala 97:16:@45463.4]
  assign rport_io_ins_151 = regs_151_io_out; // @[RegFile.scala 97:16:@45464.4]
  assign rport_io_ins_152 = regs_152_io_out; // @[RegFile.scala 97:16:@45465.4]
  assign rport_io_ins_153 = regs_153_io_out; // @[RegFile.scala 97:16:@45466.4]
  assign rport_io_ins_154 = regs_154_io_out; // @[RegFile.scala 97:16:@45467.4]
  assign rport_io_ins_155 = regs_155_io_out; // @[RegFile.scala 97:16:@45468.4]
  assign rport_io_ins_156 = regs_156_io_out; // @[RegFile.scala 97:16:@45469.4]
  assign rport_io_ins_157 = regs_157_io_out; // @[RegFile.scala 97:16:@45470.4]
  assign rport_io_ins_158 = regs_158_io_out; // @[RegFile.scala 97:16:@45471.4]
  assign rport_io_ins_159 = regs_159_io_out; // @[RegFile.scala 97:16:@45472.4]
  assign rport_io_ins_160 = regs_160_io_out; // @[RegFile.scala 97:16:@45473.4]
  assign rport_io_ins_161 = regs_161_io_out; // @[RegFile.scala 97:16:@45474.4]
  assign rport_io_ins_162 = regs_162_io_out; // @[RegFile.scala 97:16:@45475.4]
  assign rport_io_ins_163 = regs_163_io_out; // @[RegFile.scala 97:16:@45476.4]
  assign rport_io_ins_164 = regs_164_io_out; // @[RegFile.scala 97:16:@45477.4]
  assign rport_io_ins_165 = regs_165_io_out; // @[RegFile.scala 97:16:@45478.4]
  assign rport_io_ins_166 = regs_166_io_out; // @[RegFile.scala 97:16:@45479.4]
  assign rport_io_ins_167 = regs_167_io_out; // @[RegFile.scala 97:16:@45480.4]
  assign rport_io_ins_168 = regs_168_io_out; // @[RegFile.scala 97:16:@45481.4]
  assign rport_io_ins_169 = regs_169_io_out; // @[RegFile.scala 97:16:@45482.4]
  assign rport_io_ins_170 = regs_170_io_out; // @[RegFile.scala 97:16:@45483.4]
  assign rport_io_ins_171 = regs_171_io_out; // @[RegFile.scala 97:16:@45484.4]
  assign rport_io_ins_172 = regs_172_io_out; // @[RegFile.scala 97:16:@45485.4]
  assign rport_io_ins_173 = regs_173_io_out; // @[RegFile.scala 97:16:@45486.4]
  assign rport_io_ins_174 = regs_174_io_out; // @[RegFile.scala 97:16:@45487.4]
  assign rport_io_ins_175 = regs_175_io_out; // @[RegFile.scala 97:16:@45488.4]
  assign rport_io_ins_176 = regs_176_io_out; // @[RegFile.scala 97:16:@45489.4]
  assign rport_io_ins_177 = regs_177_io_out; // @[RegFile.scala 97:16:@45490.4]
  assign rport_io_ins_178 = regs_178_io_out; // @[RegFile.scala 97:16:@45491.4]
  assign rport_io_ins_179 = regs_179_io_out; // @[RegFile.scala 97:16:@45492.4]
  assign rport_io_ins_180 = regs_180_io_out; // @[RegFile.scala 97:16:@45493.4]
  assign rport_io_ins_181 = regs_181_io_out; // @[RegFile.scala 97:16:@45494.4]
  assign rport_io_ins_182 = regs_182_io_out; // @[RegFile.scala 97:16:@45495.4]
  assign rport_io_ins_183 = regs_183_io_out; // @[RegFile.scala 97:16:@45496.4]
  assign rport_io_ins_184 = regs_184_io_out; // @[RegFile.scala 97:16:@45497.4]
  assign rport_io_ins_185 = regs_185_io_out; // @[RegFile.scala 97:16:@45498.4]
  assign rport_io_ins_186 = regs_186_io_out; // @[RegFile.scala 97:16:@45499.4]
  assign rport_io_ins_187 = regs_187_io_out; // @[RegFile.scala 97:16:@45500.4]
  assign rport_io_ins_188 = regs_188_io_out; // @[RegFile.scala 97:16:@45501.4]
  assign rport_io_ins_189 = regs_189_io_out; // @[RegFile.scala 97:16:@45502.4]
  assign rport_io_ins_190 = regs_190_io_out; // @[RegFile.scala 97:16:@45503.4]
  assign rport_io_ins_191 = regs_191_io_out; // @[RegFile.scala 97:16:@45504.4]
  assign rport_io_ins_192 = regs_192_io_out; // @[RegFile.scala 97:16:@45505.4]
  assign rport_io_ins_193 = regs_193_io_out; // @[RegFile.scala 97:16:@45506.4]
  assign rport_io_ins_194 = regs_194_io_out; // @[RegFile.scala 97:16:@45507.4]
  assign rport_io_ins_195 = regs_195_io_out; // @[RegFile.scala 97:16:@45508.4]
  assign rport_io_ins_196 = regs_196_io_out; // @[RegFile.scala 97:16:@45509.4]
  assign rport_io_ins_197 = regs_197_io_out; // @[RegFile.scala 97:16:@45510.4]
  assign rport_io_ins_198 = regs_198_io_out; // @[RegFile.scala 97:16:@45511.4]
  assign rport_io_ins_199 = regs_199_io_out; // @[RegFile.scala 97:16:@45512.4]
  assign rport_io_ins_200 = regs_200_io_out; // @[RegFile.scala 97:16:@45513.4]
  assign rport_io_ins_201 = regs_201_io_out; // @[RegFile.scala 97:16:@45514.4]
  assign rport_io_ins_202 = regs_202_io_out; // @[RegFile.scala 97:16:@45515.4]
  assign rport_io_ins_203 = regs_203_io_out; // @[RegFile.scala 97:16:@45516.4]
  assign rport_io_ins_204 = regs_204_io_out; // @[RegFile.scala 97:16:@45517.4]
  assign rport_io_ins_205 = regs_205_io_out; // @[RegFile.scala 97:16:@45518.4]
  assign rport_io_ins_206 = regs_206_io_out; // @[RegFile.scala 97:16:@45519.4]
  assign rport_io_ins_207 = regs_207_io_out; // @[RegFile.scala 97:16:@45520.4]
  assign rport_io_ins_208 = regs_208_io_out; // @[RegFile.scala 97:16:@45521.4]
  assign rport_io_ins_209 = regs_209_io_out; // @[RegFile.scala 97:16:@45522.4]
  assign rport_io_ins_210 = regs_210_io_out; // @[RegFile.scala 97:16:@45523.4]
  assign rport_io_ins_211 = regs_211_io_out; // @[RegFile.scala 97:16:@45524.4]
  assign rport_io_ins_212 = regs_212_io_out; // @[RegFile.scala 97:16:@45525.4]
  assign rport_io_ins_213 = regs_213_io_out; // @[RegFile.scala 97:16:@45526.4]
  assign rport_io_ins_214 = regs_214_io_out; // @[RegFile.scala 97:16:@45527.4]
  assign rport_io_ins_215 = regs_215_io_out; // @[RegFile.scala 97:16:@45528.4]
  assign rport_io_ins_216 = regs_216_io_out; // @[RegFile.scala 97:16:@45529.4]
  assign rport_io_ins_217 = regs_217_io_out; // @[RegFile.scala 97:16:@45530.4]
  assign rport_io_ins_218 = regs_218_io_out; // @[RegFile.scala 97:16:@45531.4]
  assign rport_io_ins_219 = regs_219_io_out; // @[RegFile.scala 97:16:@45532.4]
  assign rport_io_ins_220 = regs_220_io_out; // @[RegFile.scala 97:16:@45533.4]
  assign rport_io_ins_221 = regs_221_io_out; // @[RegFile.scala 97:16:@45534.4]
  assign rport_io_ins_222 = regs_222_io_out; // @[RegFile.scala 97:16:@45535.4]
  assign rport_io_ins_223 = regs_223_io_out; // @[RegFile.scala 97:16:@45536.4]
  assign rport_io_ins_224 = regs_224_io_out; // @[RegFile.scala 97:16:@45537.4]
  assign rport_io_ins_225 = regs_225_io_out; // @[RegFile.scala 97:16:@45538.4]
  assign rport_io_ins_226 = regs_226_io_out; // @[RegFile.scala 97:16:@45539.4]
  assign rport_io_ins_227 = regs_227_io_out; // @[RegFile.scala 97:16:@45540.4]
  assign rport_io_ins_228 = regs_228_io_out; // @[RegFile.scala 97:16:@45541.4]
  assign rport_io_ins_229 = regs_229_io_out; // @[RegFile.scala 97:16:@45542.4]
  assign rport_io_ins_230 = regs_230_io_out; // @[RegFile.scala 97:16:@45543.4]
  assign rport_io_ins_231 = regs_231_io_out; // @[RegFile.scala 97:16:@45544.4]
  assign rport_io_ins_232 = regs_232_io_out; // @[RegFile.scala 97:16:@45545.4]
  assign rport_io_ins_233 = regs_233_io_out; // @[RegFile.scala 97:16:@45546.4]
  assign rport_io_ins_234 = regs_234_io_out; // @[RegFile.scala 97:16:@45547.4]
  assign rport_io_ins_235 = regs_235_io_out; // @[RegFile.scala 97:16:@45548.4]
  assign rport_io_ins_236 = regs_236_io_out; // @[RegFile.scala 97:16:@45549.4]
  assign rport_io_ins_237 = regs_237_io_out; // @[RegFile.scala 97:16:@45550.4]
  assign rport_io_ins_238 = regs_238_io_out; // @[RegFile.scala 97:16:@45551.4]
  assign rport_io_ins_239 = regs_239_io_out; // @[RegFile.scala 97:16:@45552.4]
  assign rport_io_ins_240 = regs_240_io_out; // @[RegFile.scala 97:16:@45553.4]
  assign rport_io_ins_241 = regs_241_io_out; // @[RegFile.scala 97:16:@45554.4]
  assign rport_io_ins_242 = regs_242_io_out; // @[RegFile.scala 97:16:@45555.4]
  assign rport_io_ins_243 = regs_243_io_out; // @[RegFile.scala 97:16:@45556.4]
  assign rport_io_ins_244 = regs_244_io_out; // @[RegFile.scala 97:16:@45557.4]
  assign rport_io_ins_245 = regs_245_io_out; // @[RegFile.scala 97:16:@45558.4]
  assign rport_io_ins_246 = regs_246_io_out; // @[RegFile.scala 97:16:@45559.4]
  assign rport_io_ins_247 = regs_247_io_out; // @[RegFile.scala 97:16:@45560.4]
  assign rport_io_ins_248 = regs_248_io_out; // @[RegFile.scala 97:16:@45561.4]
  assign rport_io_ins_249 = regs_249_io_out; // @[RegFile.scala 97:16:@45562.4]
  assign rport_io_ins_250 = regs_250_io_out; // @[RegFile.scala 97:16:@45563.4]
  assign rport_io_ins_251 = regs_251_io_out; // @[RegFile.scala 97:16:@45564.4]
  assign rport_io_ins_252 = regs_252_io_out; // @[RegFile.scala 97:16:@45565.4]
  assign rport_io_ins_253 = regs_253_io_out; // @[RegFile.scala 97:16:@45566.4]
  assign rport_io_ins_254 = regs_254_io_out; // @[RegFile.scala 97:16:@45567.4]
  assign rport_io_ins_255 = regs_255_io_out; // @[RegFile.scala 97:16:@45568.4]
  assign rport_io_ins_256 = regs_256_io_out; // @[RegFile.scala 97:16:@45569.4]
  assign rport_io_ins_257 = regs_257_io_out; // @[RegFile.scala 97:16:@45570.4]
  assign rport_io_ins_258 = regs_258_io_out; // @[RegFile.scala 97:16:@45571.4]
  assign rport_io_ins_259 = regs_259_io_out; // @[RegFile.scala 97:16:@45572.4]
  assign rport_io_ins_260 = regs_260_io_out; // @[RegFile.scala 97:16:@45573.4]
  assign rport_io_ins_261 = regs_261_io_out; // @[RegFile.scala 97:16:@45574.4]
  assign rport_io_ins_262 = regs_262_io_out; // @[RegFile.scala 97:16:@45575.4]
  assign rport_io_ins_263 = regs_263_io_out; // @[RegFile.scala 97:16:@45576.4]
  assign rport_io_ins_264 = regs_264_io_out; // @[RegFile.scala 97:16:@45577.4]
  assign rport_io_ins_265 = regs_265_io_out; // @[RegFile.scala 97:16:@45578.4]
  assign rport_io_ins_266 = regs_266_io_out; // @[RegFile.scala 97:16:@45579.4]
  assign rport_io_ins_267 = regs_267_io_out; // @[RegFile.scala 97:16:@45580.4]
  assign rport_io_ins_268 = regs_268_io_out; // @[RegFile.scala 97:16:@45581.4]
  assign rport_io_ins_269 = regs_269_io_out; // @[RegFile.scala 97:16:@45582.4]
  assign rport_io_ins_270 = regs_270_io_out; // @[RegFile.scala 97:16:@45583.4]
  assign rport_io_ins_271 = regs_271_io_out; // @[RegFile.scala 97:16:@45584.4]
  assign rport_io_ins_272 = regs_272_io_out; // @[RegFile.scala 97:16:@45585.4]
  assign rport_io_ins_273 = regs_273_io_out; // @[RegFile.scala 97:16:@45586.4]
  assign rport_io_ins_274 = regs_274_io_out; // @[RegFile.scala 97:16:@45587.4]
  assign rport_io_ins_275 = regs_275_io_out; // @[RegFile.scala 97:16:@45588.4]
  assign rport_io_ins_276 = regs_276_io_out; // @[RegFile.scala 97:16:@45589.4]
  assign rport_io_ins_277 = regs_277_io_out; // @[RegFile.scala 97:16:@45590.4]
  assign rport_io_ins_278 = regs_278_io_out; // @[RegFile.scala 97:16:@45591.4]
  assign rport_io_ins_279 = regs_279_io_out; // @[RegFile.scala 97:16:@45592.4]
  assign rport_io_ins_280 = regs_280_io_out; // @[RegFile.scala 97:16:@45593.4]
  assign rport_io_ins_281 = regs_281_io_out; // @[RegFile.scala 97:16:@45594.4]
  assign rport_io_ins_282 = regs_282_io_out; // @[RegFile.scala 97:16:@45595.4]
  assign rport_io_ins_283 = regs_283_io_out; // @[RegFile.scala 97:16:@45596.4]
  assign rport_io_ins_284 = regs_284_io_out; // @[RegFile.scala 97:16:@45597.4]
  assign rport_io_ins_285 = regs_285_io_out; // @[RegFile.scala 97:16:@45598.4]
  assign rport_io_ins_286 = regs_286_io_out; // @[RegFile.scala 97:16:@45599.4]
  assign rport_io_ins_287 = regs_287_io_out; // @[RegFile.scala 97:16:@45600.4]
  assign rport_io_ins_288 = regs_288_io_out; // @[RegFile.scala 97:16:@45601.4]
  assign rport_io_ins_289 = regs_289_io_out; // @[RegFile.scala 97:16:@45602.4]
  assign rport_io_ins_290 = regs_290_io_out; // @[RegFile.scala 97:16:@45603.4]
  assign rport_io_ins_291 = regs_291_io_out; // @[RegFile.scala 97:16:@45604.4]
  assign rport_io_ins_292 = regs_292_io_out; // @[RegFile.scala 97:16:@45605.4]
  assign rport_io_ins_293 = regs_293_io_out; // @[RegFile.scala 97:16:@45606.4]
  assign rport_io_ins_294 = regs_294_io_out; // @[RegFile.scala 97:16:@45607.4]
  assign rport_io_ins_295 = regs_295_io_out; // @[RegFile.scala 97:16:@45608.4]
  assign rport_io_ins_296 = regs_296_io_out; // @[RegFile.scala 97:16:@45609.4]
  assign rport_io_ins_297 = regs_297_io_out; // @[RegFile.scala 97:16:@45610.4]
  assign rport_io_ins_298 = regs_298_io_out; // @[RegFile.scala 97:16:@45611.4]
  assign rport_io_ins_299 = regs_299_io_out; // @[RegFile.scala 97:16:@45612.4]
  assign rport_io_ins_300 = regs_300_io_out; // @[RegFile.scala 97:16:@45613.4]
  assign rport_io_ins_301 = regs_301_io_out; // @[RegFile.scala 97:16:@45614.4]
  assign rport_io_ins_302 = regs_302_io_out; // @[RegFile.scala 97:16:@45615.4]
  assign rport_io_ins_303 = regs_303_io_out; // @[RegFile.scala 97:16:@45616.4]
  assign rport_io_ins_304 = regs_304_io_out; // @[RegFile.scala 97:16:@45617.4]
  assign rport_io_ins_305 = regs_305_io_out; // @[RegFile.scala 97:16:@45618.4]
  assign rport_io_ins_306 = regs_306_io_out; // @[RegFile.scala 97:16:@45619.4]
  assign rport_io_ins_307 = regs_307_io_out; // @[RegFile.scala 97:16:@45620.4]
  assign rport_io_ins_308 = regs_308_io_out; // @[RegFile.scala 97:16:@45621.4]
  assign rport_io_ins_309 = regs_309_io_out; // @[RegFile.scala 97:16:@45622.4]
  assign rport_io_ins_310 = regs_310_io_out; // @[RegFile.scala 97:16:@45623.4]
  assign rport_io_ins_311 = regs_311_io_out; // @[RegFile.scala 97:16:@45624.4]
  assign rport_io_ins_312 = regs_312_io_out; // @[RegFile.scala 97:16:@45625.4]
  assign rport_io_ins_313 = regs_313_io_out; // @[RegFile.scala 97:16:@45626.4]
  assign rport_io_ins_314 = regs_314_io_out; // @[RegFile.scala 97:16:@45627.4]
  assign rport_io_ins_315 = regs_315_io_out; // @[RegFile.scala 97:16:@45628.4]
  assign rport_io_ins_316 = regs_316_io_out; // @[RegFile.scala 97:16:@45629.4]
  assign rport_io_ins_317 = regs_317_io_out; // @[RegFile.scala 97:16:@45630.4]
  assign rport_io_ins_318 = regs_318_io_out; // @[RegFile.scala 97:16:@45631.4]
  assign rport_io_ins_319 = regs_319_io_out; // @[RegFile.scala 97:16:@45632.4]
  assign rport_io_ins_320 = regs_320_io_out; // @[RegFile.scala 97:16:@45633.4]
  assign rport_io_ins_321 = regs_321_io_out; // @[RegFile.scala 97:16:@45634.4]
  assign rport_io_ins_322 = regs_322_io_out; // @[RegFile.scala 97:16:@45635.4]
  assign rport_io_ins_323 = regs_323_io_out; // @[RegFile.scala 97:16:@45636.4]
  assign rport_io_ins_324 = regs_324_io_out; // @[RegFile.scala 97:16:@45637.4]
  assign rport_io_ins_325 = regs_325_io_out; // @[RegFile.scala 97:16:@45638.4]
  assign rport_io_ins_326 = regs_326_io_out; // @[RegFile.scala 97:16:@45639.4]
  assign rport_io_ins_327 = regs_327_io_out; // @[RegFile.scala 97:16:@45640.4]
  assign rport_io_ins_328 = regs_328_io_out; // @[RegFile.scala 97:16:@45641.4]
  assign rport_io_ins_329 = regs_329_io_out; // @[RegFile.scala 97:16:@45642.4]
  assign rport_io_ins_330 = regs_330_io_out; // @[RegFile.scala 97:16:@45643.4]
  assign rport_io_ins_331 = regs_331_io_out; // @[RegFile.scala 97:16:@45644.4]
  assign rport_io_ins_332 = regs_332_io_out; // @[RegFile.scala 97:16:@45645.4]
  assign rport_io_ins_333 = regs_333_io_out; // @[RegFile.scala 97:16:@45646.4]
  assign rport_io_ins_334 = regs_334_io_out; // @[RegFile.scala 97:16:@45647.4]
  assign rport_io_ins_335 = regs_335_io_out; // @[RegFile.scala 97:16:@45648.4]
  assign rport_io_ins_336 = regs_336_io_out; // @[RegFile.scala 97:16:@45649.4]
  assign rport_io_ins_337 = regs_337_io_out; // @[RegFile.scala 97:16:@45650.4]
  assign rport_io_ins_338 = regs_338_io_out; // @[RegFile.scala 97:16:@45651.4]
  assign rport_io_ins_339 = regs_339_io_out; // @[RegFile.scala 97:16:@45652.4]
  assign rport_io_ins_340 = regs_340_io_out; // @[RegFile.scala 97:16:@45653.4]
  assign rport_io_ins_341 = regs_341_io_out; // @[RegFile.scala 97:16:@45654.4]
  assign rport_io_ins_342 = regs_342_io_out; // @[RegFile.scala 97:16:@45655.4]
  assign rport_io_ins_343 = regs_343_io_out; // @[RegFile.scala 97:16:@45656.4]
  assign rport_io_ins_344 = regs_344_io_out; // @[RegFile.scala 97:16:@45657.4]
  assign rport_io_ins_345 = regs_345_io_out; // @[RegFile.scala 97:16:@45658.4]
  assign rport_io_ins_346 = regs_346_io_out; // @[RegFile.scala 97:16:@45659.4]
  assign rport_io_ins_347 = regs_347_io_out; // @[RegFile.scala 97:16:@45660.4]
  assign rport_io_ins_348 = regs_348_io_out; // @[RegFile.scala 97:16:@45661.4]
  assign rport_io_ins_349 = regs_349_io_out; // @[RegFile.scala 97:16:@45662.4]
  assign rport_io_ins_350 = regs_350_io_out; // @[RegFile.scala 97:16:@45663.4]
  assign rport_io_ins_351 = regs_351_io_out; // @[RegFile.scala 97:16:@45664.4]
  assign rport_io_ins_352 = regs_352_io_out; // @[RegFile.scala 97:16:@45665.4]
  assign rport_io_ins_353 = regs_353_io_out; // @[RegFile.scala 97:16:@45666.4]
  assign rport_io_ins_354 = regs_354_io_out; // @[RegFile.scala 97:16:@45667.4]
  assign rport_io_ins_355 = regs_355_io_out; // @[RegFile.scala 97:16:@45668.4]
  assign rport_io_ins_356 = regs_356_io_out; // @[RegFile.scala 97:16:@45669.4]
  assign rport_io_ins_357 = regs_357_io_out; // @[RegFile.scala 97:16:@45670.4]
  assign rport_io_ins_358 = regs_358_io_out; // @[RegFile.scala 97:16:@45671.4]
  assign rport_io_ins_359 = regs_359_io_out; // @[RegFile.scala 97:16:@45672.4]
  assign rport_io_ins_360 = regs_360_io_out; // @[RegFile.scala 97:16:@45673.4]
  assign rport_io_ins_361 = regs_361_io_out; // @[RegFile.scala 97:16:@45674.4]
  assign rport_io_ins_362 = regs_362_io_out; // @[RegFile.scala 97:16:@45675.4]
  assign rport_io_ins_363 = regs_363_io_out; // @[RegFile.scala 97:16:@45676.4]
  assign rport_io_ins_364 = regs_364_io_out; // @[RegFile.scala 97:16:@45677.4]
  assign rport_io_ins_365 = regs_365_io_out; // @[RegFile.scala 97:16:@45678.4]
  assign rport_io_ins_366 = regs_366_io_out; // @[RegFile.scala 97:16:@45679.4]
  assign rport_io_ins_367 = regs_367_io_out; // @[RegFile.scala 97:16:@45680.4]
  assign rport_io_ins_368 = regs_368_io_out; // @[RegFile.scala 97:16:@45681.4]
  assign rport_io_ins_369 = regs_369_io_out; // @[RegFile.scala 97:16:@45682.4]
  assign rport_io_ins_370 = regs_370_io_out; // @[RegFile.scala 97:16:@45683.4]
  assign rport_io_ins_371 = regs_371_io_out; // @[RegFile.scala 97:16:@45684.4]
  assign rport_io_ins_372 = regs_372_io_out; // @[RegFile.scala 97:16:@45685.4]
  assign rport_io_ins_373 = regs_373_io_out; // @[RegFile.scala 97:16:@45686.4]
  assign rport_io_ins_374 = regs_374_io_out; // @[RegFile.scala 97:16:@45687.4]
  assign rport_io_ins_375 = regs_375_io_out; // @[RegFile.scala 97:16:@45688.4]
  assign rport_io_ins_376 = regs_376_io_out; // @[RegFile.scala 97:16:@45689.4]
  assign rport_io_ins_377 = regs_377_io_out; // @[RegFile.scala 97:16:@45690.4]
  assign rport_io_ins_378 = regs_378_io_out; // @[RegFile.scala 97:16:@45691.4]
  assign rport_io_ins_379 = regs_379_io_out; // @[RegFile.scala 97:16:@45692.4]
  assign rport_io_ins_380 = regs_380_io_out; // @[RegFile.scala 97:16:@45693.4]
  assign rport_io_ins_381 = regs_381_io_out; // @[RegFile.scala 97:16:@45694.4]
  assign rport_io_ins_382 = regs_382_io_out; // @[RegFile.scala 97:16:@45695.4]
  assign rport_io_ins_383 = regs_383_io_out; // @[RegFile.scala 97:16:@45696.4]
  assign rport_io_ins_384 = regs_384_io_out; // @[RegFile.scala 97:16:@45697.4]
  assign rport_io_ins_385 = regs_385_io_out; // @[RegFile.scala 97:16:@45698.4]
  assign rport_io_ins_386 = regs_386_io_out; // @[RegFile.scala 97:16:@45699.4]
  assign rport_io_ins_387 = regs_387_io_out; // @[RegFile.scala 97:16:@45700.4]
  assign rport_io_ins_388 = regs_388_io_out; // @[RegFile.scala 97:16:@45701.4]
  assign rport_io_ins_389 = regs_389_io_out; // @[RegFile.scala 97:16:@45702.4]
  assign rport_io_ins_390 = regs_390_io_out; // @[RegFile.scala 97:16:@45703.4]
  assign rport_io_ins_391 = regs_391_io_out; // @[RegFile.scala 97:16:@45704.4]
  assign rport_io_ins_392 = regs_392_io_out; // @[RegFile.scala 97:16:@45705.4]
  assign rport_io_ins_393 = regs_393_io_out; // @[RegFile.scala 97:16:@45706.4]
  assign rport_io_ins_394 = regs_394_io_out; // @[RegFile.scala 97:16:@45707.4]
  assign rport_io_ins_395 = regs_395_io_out; // @[RegFile.scala 97:16:@45708.4]
  assign rport_io_ins_396 = regs_396_io_out; // @[RegFile.scala 97:16:@45709.4]
  assign rport_io_ins_397 = regs_397_io_out; // @[RegFile.scala 97:16:@45710.4]
  assign rport_io_ins_398 = regs_398_io_out; // @[RegFile.scala 97:16:@45711.4]
  assign rport_io_ins_399 = regs_399_io_out; // @[RegFile.scala 97:16:@45712.4]
  assign rport_io_ins_400 = regs_400_io_out; // @[RegFile.scala 97:16:@45713.4]
  assign rport_io_ins_401 = regs_401_io_out; // @[RegFile.scala 97:16:@45714.4]
  assign rport_io_ins_402 = regs_402_io_out; // @[RegFile.scala 97:16:@45715.4]
  assign rport_io_ins_403 = regs_403_io_out; // @[RegFile.scala 97:16:@45716.4]
  assign rport_io_ins_404 = regs_404_io_out; // @[RegFile.scala 97:16:@45717.4]
  assign rport_io_ins_405 = regs_405_io_out; // @[RegFile.scala 97:16:@45718.4]
  assign rport_io_ins_406 = regs_406_io_out; // @[RegFile.scala 97:16:@45719.4]
  assign rport_io_ins_407 = regs_407_io_out; // @[RegFile.scala 97:16:@45720.4]
  assign rport_io_ins_408 = regs_408_io_out; // @[RegFile.scala 97:16:@45721.4]
  assign rport_io_ins_409 = regs_409_io_out; // @[RegFile.scala 97:16:@45722.4]
  assign rport_io_ins_410 = regs_410_io_out; // @[RegFile.scala 97:16:@45723.4]
  assign rport_io_ins_411 = regs_411_io_out; // @[RegFile.scala 97:16:@45724.4]
  assign rport_io_ins_412 = regs_412_io_out; // @[RegFile.scala 97:16:@45725.4]
  assign rport_io_ins_413 = regs_413_io_out; // @[RegFile.scala 97:16:@45726.4]
  assign rport_io_ins_414 = regs_414_io_out; // @[RegFile.scala 97:16:@45727.4]
  assign rport_io_ins_415 = regs_415_io_out; // @[RegFile.scala 97:16:@45728.4]
  assign rport_io_ins_416 = regs_416_io_out; // @[RegFile.scala 97:16:@45729.4]
  assign rport_io_ins_417 = regs_417_io_out; // @[RegFile.scala 97:16:@45730.4]
  assign rport_io_ins_418 = regs_418_io_out; // @[RegFile.scala 97:16:@45731.4]
  assign rport_io_ins_419 = regs_419_io_out; // @[RegFile.scala 97:16:@45732.4]
  assign rport_io_ins_420 = regs_420_io_out; // @[RegFile.scala 97:16:@45733.4]
  assign rport_io_ins_421 = regs_421_io_out; // @[RegFile.scala 97:16:@45734.4]
  assign rport_io_ins_422 = regs_422_io_out; // @[RegFile.scala 97:16:@45735.4]
  assign rport_io_ins_423 = regs_423_io_out; // @[RegFile.scala 97:16:@45736.4]
  assign rport_io_ins_424 = regs_424_io_out; // @[RegFile.scala 97:16:@45737.4]
  assign rport_io_ins_425 = regs_425_io_out; // @[RegFile.scala 97:16:@45738.4]
  assign rport_io_ins_426 = regs_426_io_out; // @[RegFile.scala 97:16:@45739.4]
  assign rport_io_ins_427 = regs_427_io_out; // @[RegFile.scala 97:16:@45740.4]
  assign rport_io_ins_428 = regs_428_io_out; // @[RegFile.scala 97:16:@45741.4]
  assign rport_io_ins_429 = regs_429_io_out; // @[RegFile.scala 97:16:@45742.4]
  assign rport_io_ins_430 = regs_430_io_out; // @[RegFile.scala 97:16:@45743.4]
  assign rport_io_ins_431 = regs_431_io_out; // @[RegFile.scala 97:16:@45744.4]
  assign rport_io_ins_432 = regs_432_io_out; // @[RegFile.scala 97:16:@45745.4]
  assign rport_io_ins_433 = regs_433_io_out; // @[RegFile.scala 97:16:@45746.4]
  assign rport_io_ins_434 = regs_434_io_out; // @[RegFile.scala 97:16:@45747.4]
  assign rport_io_ins_435 = regs_435_io_out; // @[RegFile.scala 97:16:@45748.4]
  assign rport_io_ins_436 = regs_436_io_out; // @[RegFile.scala 97:16:@45749.4]
  assign rport_io_ins_437 = regs_437_io_out; // @[RegFile.scala 97:16:@45750.4]
  assign rport_io_ins_438 = regs_438_io_out; // @[RegFile.scala 97:16:@45751.4]
  assign rport_io_ins_439 = regs_439_io_out; // @[RegFile.scala 97:16:@45752.4]
  assign rport_io_ins_440 = regs_440_io_out; // @[RegFile.scala 97:16:@45753.4]
  assign rport_io_ins_441 = regs_441_io_out; // @[RegFile.scala 97:16:@45754.4]
  assign rport_io_ins_442 = regs_442_io_out; // @[RegFile.scala 97:16:@45755.4]
  assign rport_io_ins_443 = regs_443_io_out; // @[RegFile.scala 97:16:@45756.4]
  assign rport_io_ins_444 = regs_444_io_out; // @[RegFile.scala 97:16:@45757.4]
  assign rport_io_ins_445 = regs_445_io_out; // @[RegFile.scala 97:16:@45758.4]
  assign rport_io_ins_446 = regs_446_io_out; // @[RegFile.scala 97:16:@45759.4]
  assign rport_io_ins_447 = regs_447_io_out; // @[RegFile.scala 97:16:@45760.4]
  assign rport_io_ins_448 = regs_448_io_out; // @[RegFile.scala 97:16:@45761.4]
  assign rport_io_ins_449 = regs_449_io_out; // @[RegFile.scala 97:16:@45762.4]
  assign rport_io_ins_450 = regs_450_io_out; // @[RegFile.scala 97:16:@45763.4]
  assign rport_io_ins_451 = regs_451_io_out; // @[RegFile.scala 97:16:@45764.4]
  assign rport_io_ins_452 = regs_452_io_out; // @[RegFile.scala 97:16:@45765.4]
  assign rport_io_ins_453 = regs_453_io_out; // @[RegFile.scala 97:16:@45766.4]
  assign rport_io_ins_454 = regs_454_io_out; // @[RegFile.scala 97:16:@45767.4]
  assign rport_io_ins_455 = regs_455_io_out; // @[RegFile.scala 97:16:@45768.4]
  assign rport_io_ins_456 = regs_456_io_out; // @[RegFile.scala 97:16:@45769.4]
  assign rport_io_ins_457 = regs_457_io_out; // @[RegFile.scala 97:16:@45770.4]
  assign rport_io_ins_458 = regs_458_io_out; // @[RegFile.scala 97:16:@45771.4]
  assign rport_io_ins_459 = regs_459_io_out; // @[RegFile.scala 97:16:@45772.4]
  assign rport_io_ins_460 = regs_460_io_out; // @[RegFile.scala 97:16:@45773.4]
  assign rport_io_ins_461 = regs_461_io_out; // @[RegFile.scala 97:16:@45774.4]
  assign rport_io_ins_462 = regs_462_io_out; // @[RegFile.scala 97:16:@45775.4]
  assign rport_io_ins_463 = regs_463_io_out; // @[RegFile.scala 97:16:@45776.4]
  assign rport_io_ins_464 = regs_464_io_out; // @[RegFile.scala 97:16:@45777.4]
  assign rport_io_ins_465 = regs_465_io_out; // @[RegFile.scala 97:16:@45778.4]
  assign rport_io_ins_466 = regs_466_io_out; // @[RegFile.scala 97:16:@45779.4]
  assign rport_io_ins_467 = regs_467_io_out; // @[RegFile.scala 97:16:@45780.4]
  assign rport_io_ins_468 = regs_468_io_out; // @[RegFile.scala 97:16:@45781.4]
  assign rport_io_ins_469 = regs_469_io_out; // @[RegFile.scala 97:16:@45782.4]
  assign rport_io_ins_470 = regs_470_io_out; // @[RegFile.scala 97:16:@45783.4]
  assign rport_io_ins_471 = regs_471_io_out; // @[RegFile.scala 97:16:@45784.4]
  assign rport_io_ins_472 = regs_472_io_out; // @[RegFile.scala 97:16:@45785.4]
  assign rport_io_ins_473 = regs_473_io_out; // @[RegFile.scala 97:16:@45786.4]
  assign rport_io_ins_474 = regs_474_io_out; // @[RegFile.scala 97:16:@45787.4]
  assign rport_io_ins_475 = regs_475_io_out; // @[RegFile.scala 97:16:@45788.4]
  assign rport_io_ins_476 = regs_476_io_out; // @[RegFile.scala 97:16:@45789.4]
  assign rport_io_ins_477 = regs_477_io_out; // @[RegFile.scala 97:16:@45790.4]
  assign rport_io_ins_478 = regs_478_io_out; // @[RegFile.scala 97:16:@45791.4]
  assign rport_io_ins_479 = regs_479_io_out; // @[RegFile.scala 97:16:@45792.4]
  assign rport_io_ins_480 = regs_480_io_out; // @[RegFile.scala 97:16:@45793.4]
  assign rport_io_ins_481 = regs_481_io_out; // @[RegFile.scala 97:16:@45794.4]
  assign rport_io_ins_482 = regs_482_io_out; // @[RegFile.scala 97:16:@45795.4]
  assign rport_io_ins_483 = regs_483_io_out; // @[RegFile.scala 97:16:@45796.4]
  assign rport_io_ins_484 = regs_484_io_out; // @[RegFile.scala 97:16:@45797.4]
  assign rport_io_ins_485 = regs_485_io_out; // @[RegFile.scala 97:16:@45798.4]
  assign rport_io_ins_486 = regs_486_io_out; // @[RegFile.scala 97:16:@45799.4]
  assign rport_io_ins_487 = regs_487_io_out; // @[RegFile.scala 97:16:@45800.4]
  assign rport_io_ins_488 = regs_488_io_out; // @[RegFile.scala 97:16:@45801.4]
  assign rport_io_ins_489 = regs_489_io_out; // @[RegFile.scala 97:16:@45802.4]
  assign rport_io_ins_490 = regs_490_io_out; // @[RegFile.scala 97:16:@45803.4]
  assign rport_io_ins_491 = regs_491_io_out; // @[RegFile.scala 97:16:@45804.4]
  assign rport_io_ins_492 = regs_492_io_out; // @[RegFile.scala 97:16:@45805.4]
  assign rport_io_ins_493 = regs_493_io_out; // @[RegFile.scala 97:16:@45806.4]
  assign rport_io_ins_494 = regs_494_io_out; // @[RegFile.scala 97:16:@45807.4]
  assign rport_io_ins_495 = regs_495_io_out; // @[RegFile.scala 97:16:@45808.4]
  assign rport_io_ins_496 = regs_496_io_out; // @[RegFile.scala 97:16:@45809.4]
  assign rport_io_ins_497 = regs_497_io_out; // @[RegFile.scala 97:16:@45810.4]
  assign rport_io_ins_498 = regs_498_io_out; // @[RegFile.scala 97:16:@45811.4]
  assign rport_io_ins_499 = regs_499_io_out; // @[RegFile.scala 97:16:@45812.4]
  assign rport_io_ins_500 = regs_500_io_out; // @[RegFile.scala 97:16:@45813.4]
  assign rport_io_ins_501 = regs_501_io_out; // @[RegFile.scala 97:16:@45814.4]
  assign rport_io_ins_502 = regs_502_io_out; // @[RegFile.scala 97:16:@45815.4]
  assign rport_io_ins_503 = regs_503_io_out; // @[RegFile.scala 97:16:@45816.4]
  assign rport_io_ins_504 = regs_504_io_out; // @[RegFile.scala 97:16:@45817.4]
  assign rport_io_ins_505 = regs_505_io_out; // @[RegFile.scala 97:16:@45818.4]
  assign rport_io_ins_506 = regs_506_io_out; // @[RegFile.scala 97:16:@45819.4]
  assign rport_io_ins_507 = regs_507_io_out; // @[RegFile.scala 97:16:@45820.4]
  assign rport_io_ins_508 = regs_508_io_out; // @[RegFile.scala 97:16:@45821.4]
  assign rport_io_ins_509 = regs_509_io_out; // @[RegFile.scala 97:16:@45822.4]
  assign rport_io_ins_510 = regs_510_io_out; // @[RegFile.scala 97:16:@45823.4]
  assign rport_io_ins_511 = regs_511_io_out; // @[RegFile.scala 97:16:@45824.4]
  assign rport_io_sel = io_raddr[8:0]; // @[RegFile.scala 106:18:@45825.4]
endmodule
module RetimeWrapper_553( // @[:@45847.2]
  input         clock, // @[:@45848.4]
  input         reset, // @[:@45849.4]
  input  [39:0] io_in, // @[:@45850.4]
  output [39:0] io_out // @[:@45850.4]
);
  wire [39:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@45852.4]
  wire [39:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@45852.4]
  wire [39:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@45852.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@45852.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@45852.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@45852.4]
  RetimeShiftRegister #(.WIDTH(40), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@45852.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@45865.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@45864.4]
  assign sr_init = 40'h0; // @[RetimeShiftRegister.scala 19:16:@45863.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@45862.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@45861.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@45859.4]
endmodule
module FringeFF_512( // @[:@45867.2]
  input         clock, // @[:@45868.4]
  input         reset, // @[:@45869.4]
  input  [39:0] io_in, // @[:@45870.4]
  output [39:0] io_out, // @[:@45870.4]
  input         io_enable // @[:@45870.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@45873.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@45873.4]
  wire [39:0] RetimeWrapper_io_in; // @[package.scala 93:22:@45873.4]
  wire [39:0] RetimeWrapper_io_out; // @[package.scala 93:22:@45873.4]
  wire [39:0] _T_18; // @[package.scala 96:25:@45878.4 package.scala 96:25:@45879.4]
  RetimeWrapper_553 RetimeWrapper ( // @[package.scala 93:22:@45873.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@45878.4 package.scala 96:25:@45879.4]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@45890.4]
  assign RetimeWrapper_clock = clock; // @[:@45874.4]
  assign RetimeWrapper_reset = reset; // @[:@45875.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _T_18; // @[package.scala 94:16:@45876.4]
endmodule
module FringeCounter( // @[:@45892.2]
  input   clock, // @[:@45893.4]
  input   reset, // @[:@45894.4]
  input   io_enable, // @[:@45895.4]
  output  io_done // @[:@45895.4]
);
  wire  reg$_clock; // @[FringeCounter.scala 24:19:@45897.4]
  wire  reg$_reset; // @[FringeCounter.scala 24:19:@45897.4]
  wire [39:0] reg$_io_in; // @[FringeCounter.scala 24:19:@45897.4]
  wire [39:0] reg$_io_out; // @[FringeCounter.scala 24:19:@45897.4]
  wire  reg$_io_enable; // @[FringeCounter.scala 24:19:@45897.4]
  wire [40:0] count; // @[Cat.scala 30:58:@45904.4]
  wire [41:0] _T_25; // @[FringeCounter.scala 31:22:@45905.4]
  wire [40:0] newval; // @[FringeCounter.scala 31:22:@45906.4]
  wire  isMax; // @[FringeCounter.scala 32:22:@45907.4]
  wire [40:0] next; // @[FringeCounter.scala 33:17:@45909.4]
  FringeFF_512 reg$ ( // @[FringeCounter.scala 24:19:@45897.4]
    .clock(reg$_clock),
    .reset(reg$_reset),
    .io_in(reg$_io_in),
    .io_out(reg$_io_out),
    .io_enable(reg$_io_enable)
  );
  assign count = {1'h0,reg$_io_out}; // @[Cat.scala 30:58:@45904.4]
  assign _T_25 = count + 41'h1; // @[FringeCounter.scala 31:22:@45905.4]
  assign newval = count + 41'h1; // @[FringeCounter.scala 31:22:@45906.4]
  assign isMax = newval >= 41'h2cb417800; // @[FringeCounter.scala 32:22:@45907.4]
  assign next = isMax ? count : newval; // @[FringeCounter.scala 33:17:@45909.4]
  assign io_done = io_enable & isMax; // @[FringeCounter.scala 43:11:@45920.4]
  assign reg$_clock = clock; // @[:@45898.4]
  assign reg$_reset = reset; // @[:@45899.4]
  assign reg$_io_in = next[39:0]; // @[FringeCounter.scala 35:15:@45911.6 FringeCounter.scala 37:15:@45914.6]
  assign reg$_io_enable = io_enable; // @[FringeCounter.scala 27:17:@45902.4]
endmodule
module FringeFF_513( // @[:@45954.2]
  input   clock, // @[:@45955.4]
  input   reset, // @[:@45956.4]
  input   io_in, // @[:@45957.4]
  input   io_reset, // @[:@45957.4]
  output  io_out, // @[:@45957.4]
  input   io_enable // @[:@45957.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@45960.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@45960.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@45960.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@45960.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@45960.4]
  wire  _T_18; // @[package.scala 96:25:@45965.4 package.scala 96:25:@45966.4]
  wire  _GEN_0; // @[FringeFF.scala 21:27:@45971.6]
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@45960.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@45965.4 package.scala 96:25:@45966.4]
  assign _GEN_0 = io_reset ? 1'h0 : _T_18; // @[FringeFF.scala 21:27:@45971.6]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@45977.4]
  assign RetimeWrapper_clock = clock; // @[:@45961.4]
  assign RetimeWrapper_reset = reset; // @[:@45962.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@45964.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _GEN_0; // @[package.scala 94:16:@45963.4]
endmodule
module Depulser( // @[:@45979.2]
  input   clock, // @[:@45980.4]
  input   reset, // @[:@45981.4]
  input   io_in, // @[:@45982.4]
  input   io_rst, // @[:@45982.4]
  output  io_out // @[:@45982.4]
);
  wire  r_clock; // @[Depulser.scala 14:17:@45984.4]
  wire  r_reset; // @[Depulser.scala 14:17:@45984.4]
  wire  r_io_in; // @[Depulser.scala 14:17:@45984.4]
  wire  r_io_reset; // @[Depulser.scala 14:17:@45984.4]
  wire  r_io_out; // @[Depulser.scala 14:17:@45984.4]
  wire  r_io_enable; // @[Depulser.scala 14:17:@45984.4]
  FringeFF_513 r ( // @[Depulser.scala 14:17:@45984.4]
    .clock(r_clock),
    .reset(r_reset),
    .io_in(r_io_in),
    .io_reset(r_io_reset),
    .io_out(r_io_out),
    .io_enable(r_io_enable)
  );
  assign io_out = r_io_out; // @[Depulser.scala 19:10:@45993.4]
  assign r_clock = clock; // @[:@45985.4]
  assign r_reset = reset; // @[:@45986.4]
  assign r_io_in = io_rst ? 1'h0 : io_in; // @[Depulser.scala 15:11:@45988.4]
  assign r_io_reset = io_rst; // @[Depulser.scala 18:14:@45992.4]
  assign r_io_enable = io_in | io_rst; // @[Depulser.scala 17:15:@45991.4]
endmodule
module Fringe( // @[:@45995.2]
  input         clock, // @[:@45996.4]
  input         reset, // @[:@45997.4]
  input  [31:0] io_raddr, // @[:@45998.4]
  input         io_wen, // @[:@45998.4]
  input  [31:0] io_waddr, // @[:@45998.4]
  input  [63:0] io_wdata, // @[:@45998.4]
  output [63:0] io_rdata, // @[:@45998.4]
  output        io_enable, // @[:@45998.4]
  input         io_done, // @[:@45998.4]
  output        io_reset, // @[:@45998.4]
  output [63:0] io_argIns_0, // @[:@45998.4]
  input         io_argOuts_0_valid, // @[:@45998.4]
  input  [63:0] io_argOuts_0_bits, // @[:@45998.4]
  input         io_argOuts_1_valid, // @[:@45998.4]
  input  [63:0] io_argOuts_1_bits, // @[:@45998.4]
  input         io_argOuts_2_valid, // @[:@45998.4]
  input  [63:0] io_argOuts_2_bits, // @[:@45998.4]
  input         io_argOuts_3_valid, // @[:@45998.4]
  input  [63:0] io_argOuts_3_bits, // @[:@45998.4]
  input         io_argOuts_4_valid, // @[:@45998.4]
  input  [63:0] io_argOuts_4_bits, // @[:@45998.4]
  input         io_argOuts_5_valid, // @[:@45998.4]
  input  [63:0] io_argOuts_5_bits, // @[:@45998.4]
  input         io_argOuts_6_valid, // @[:@45998.4]
  input  [63:0] io_argOuts_6_bits, // @[:@45998.4]
  input         io_argOuts_7_valid, // @[:@45998.4]
  input  [63:0] io_argOuts_7_bits, // @[:@45998.4]
  input         io_argOuts_8_valid, // @[:@45998.4]
  input  [63:0] io_argOuts_8_bits, // @[:@45998.4]
  input         io_argOuts_9_valid, // @[:@45998.4]
  input  [63:0] io_argOuts_9_bits, // @[:@45998.4]
  input         io_heap_0_req_valid, // @[:@45998.4]
  input         io_heap_0_req_bits_allocDealloc, // @[:@45998.4]
  input  [63:0] io_heap_0_req_bits_sizeAddr, // @[:@45998.4]
  output        io_heap_0_resp_valid, // @[:@45998.4]
  output        io_heap_0_resp_bits_allocDealloc, // @[:@45998.4]
  output [63:0] io_heap_0_resp_bits_sizeAddr // @[:@45998.4]
);
  wire  heap_io_accel_0_req_valid; // @[Fringe.scala 107:20:@47063.4]
  wire  heap_io_accel_0_req_bits_allocDealloc; // @[Fringe.scala 107:20:@47063.4]
  wire [63:0] heap_io_accel_0_req_bits_sizeAddr; // @[Fringe.scala 107:20:@47063.4]
  wire  heap_io_accel_0_resp_valid; // @[Fringe.scala 107:20:@47063.4]
  wire  heap_io_accel_0_resp_bits_allocDealloc; // @[Fringe.scala 107:20:@47063.4]
  wire [63:0] heap_io_accel_0_resp_bits_sizeAddr; // @[Fringe.scala 107:20:@47063.4]
  wire  heap_io_host_0_req_valid; // @[Fringe.scala 107:20:@47063.4]
  wire  heap_io_host_0_req_bits_allocDealloc; // @[Fringe.scala 107:20:@47063.4]
  wire [63:0] heap_io_host_0_req_bits_sizeAddr; // @[Fringe.scala 107:20:@47063.4]
  wire  heap_io_host_0_resp_valid; // @[Fringe.scala 107:20:@47063.4]
  wire  heap_io_host_0_resp_bits_allocDealloc; // @[Fringe.scala 107:20:@47063.4]
  wire [63:0] heap_io_host_0_resp_bits_sizeAddr; // @[Fringe.scala 107:20:@47063.4]
  wire  regs_clock; // @[Fringe.scala 116:20:@47072.4]
  wire  regs_reset; // @[Fringe.scala 116:20:@47072.4]
  wire [31:0] regs_io_raddr; // @[Fringe.scala 116:20:@47072.4]
  wire  regs_io_wen; // @[Fringe.scala 116:20:@47072.4]
  wire [31:0] regs_io_waddr; // @[Fringe.scala 116:20:@47072.4]
  wire [63:0] regs_io_wdata; // @[Fringe.scala 116:20:@47072.4]
  wire [63:0] regs_io_rdata; // @[Fringe.scala 116:20:@47072.4]
  wire  regs_io_reset; // @[Fringe.scala 116:20:@47072.4]
  wire [63:0] regs_io_argIns_0; // @[Fringe.scala 116:20:@47072.4]
  wire [63:0] regs_io_argIns_1; // @[Fringe.scala 116:20:@47072.4]
  wire [63:0] regs_io_argIns_2; // @[Fringe.scala 116:20:@47072.4]
  wire  regs_io_argOuts_0_valid; // @[Fringe.scala 116:20:@47072.4]
  wire [63:0] regs_io_argOuts_0_bits; // @[Fringe.scala 116:20:@47072.4]
  wire  regs_io_argOuts_1_valid; // @[Fringe.scala 116:20:@47072.4]
  wire [63:0] regs_io_argOuts_1_bits; // @[Fringe.scala 116:20:@47072.4]
  wire  regs_io_argOuts_2_valid; // @[Fringe.scala 116:20:@47072.4]
  wire [63:0] regs_io_argOuts_2_bits; // @[Fringe.scala 116:20:@47072.4]
  wire  regs_io_argOuts_3_valid; // @[Fringe.scala 116:20:@47072.4]
  wire [63:0] regs_io_argOuts_3_bits; // @[Fringe.scala 116:20:@47072.4]
  wire  regs_io_argOuts_4_valid; // @[Fringe.scala 116:20:@47072.4]
  wire [63:0] regs_io_argOuts_4_bits; // @[Fringe.scala 116:20:@47072.4]
  wire  regs_io_argOuts_5_valid; // @[Fringe.scala 116:20:@47072.4]
  wire [63:0] regs_io_argOuts_5_bits; // @[Fringe.scala 116:20:@47072.4]
  wire  regs_io_argOuts_6_valid; // @[Fringe.scala 116:20:@47072.4]
  wire [63:0] regs_io_argOuts_6_bits; // @[Fringe.scala 116:20:@47072.4]
  wire  regs_io_argOuts_7_valid; // @[Fringe.scala 116:20:@47072.4]
  wire [63:0] regs_io_argOuts_7_bits; // @[Fringe.scala 116:20:@47072.4]
  wire  regs_io_argOuts_8_valid; // @[Fringe.scala 116:20:@47072.4]
  wire [63:0] regs_io_argOuts_8_bits; // @[Fringe.scala 116:20:@47072.4]
  wire  regs_io_argOuts_9_valid; // @[Fringe.scala 116:20:@47072.4]
  wire [63:0] regs_io_argOuts_9_bits; // @[Fringe.scala 116:20:@47072.4]
  wire  regs_io_argOuts_10_valid; // @[Fringe.scala 116:20:@47072.4]
  wire [63:0] regs_io_argOuts_10_bits; // @[Fringe.scala 116:20:@47072.4]
  wire  timeoutCtr_clock; // @[Fringe.scala 143:26:@49157.4]
  wire  timeoutCtr_reset; // @[Fringe.scala 143:26:@49157.4]
  wire  timeoutCtr_io_enable; // @[Fringe.scala 143:26:@49157.4]
  wire  timeoutCtr_io_done; // @[Fringe.scala 143:26:@49157.4]
  wire  depulser_clock; // @[Fringe.scala 153:24:@49175.4]
  wire  depulser_reset; // @[Fringe.scala 153:24:@49175.4]
  wire  depulser_io_in; // @[Fringe.scala 153:24:@49175.4]
  wire  depulser_io_rst; // @[Fringe.scala 153:24:@49175.4]
  wire  depulser_io_out; // @[Fringe.scala 153:24:@49175.4]
  wire [63:0] _T_880; // @[:@49134.4 :@49135.4]
  wire  curStatus_done; // @[Fringe.scala 133:45:@49136.4]
  wire  curStatus_timeout; // @[Fringe.scala 133:45:@49138.4]
  wire [2:0] curStatus_allocDealloc; // @[Fringe.scala 133:45:@49140.4]
  wire [58:0] curStatus_sizeAddr; // @[Fringe.scala 133:45:@49142.4]
  wire  _T_885; // @[Fringe.scala 134:28:@49144.4]
  wire  _T_889; // @[Fringe.scala 134:42:@49146.4]
  wire  _T_890; // @[Fringe.scala 135:27:@49148.4]
  wire [63:0] _T_900; // @[Fringe.scala 156:22:@49183.4]
  reg  _T_907; // @[package.scala 152:20:@49186.4]
  reg [31:0] _RAND_0;
  wire  _T_908; // @[package.scala 153:13:@49188.4]
  wire  _T_909; // @[package.scala 153:8:@49189.4]
  wire  _T_912; // @[Fringe.scala 160:55:@49193.4]
  wire  status_bits_done; // @[Fringe.scala 160:26:@49194.4]
  wire  _T_915; // @[Fringe.scala 161:58:@49197.4]
  wire  status_bits_timeout; // @[Fringe.scala 161:29:@49198.4]
  wire [1:0] _T_919; // @[Fringe.scala 162:57:@49200.4]
  wire [1:0] _T_921; // @[Fringe.scala 162:34:@49201.4]
  wire [63:0] _T_923; // @[Fringe.scala 163:30:@49203.4]
  wire [1:0] _T_924; // @[Fringe.scala 171:37:@49206.4]
  wire [58:0] status_bits_sizeAddr; // @[Fringe.scala 158:20:@49185.4 Fringe.scala 163:24:@49204.4]
  wire [2:0] status_bits_allocDealloc; // @[Fringe.scala 158:20:@49185.4 Fringe.scala 162:28:@49202.4]
  wire [61:0] _T_925; // @[Fringe.scala 171:37:@49207.4]
  wire  alloc; // @[Fringe.scala 202:38:@50519.4]
  wire  dealloc; // @[Fringe.scala 203:40:@50520.4]
  wire  _T_1429; // @[Fringe.scala 204:37:@50521.4]
  reg  _T_1432; // @[package.scala 152:20:@50522.4]
  reg [31:0] _RAND_1;
  wire  _T_1433; // @[package.scala 153:13:@50524.4]
  DRAMHeap heap ( // @[Fringe.scala 107:20:@47063.4]
    .io_accel_0_req_valid(heap_io_accel_0_req_valid),
    .io_accel_0_req_bits_allocDealloc(heap_io_accel_0_req_bits_allocDealloc),
    .io_accel_0_req_bits_sizeAddr(heap_io_accel_0_req_bits_sizeAddr),
    .io_accel_0_resp_valid(heap_io_accel_0_resp_valid),
    .io_accel_0_resp_bits_allocDealloc(heap_io_accel_0_resp_bits_allocDealloc),
    .io_accel_0_resp_bits_sizeAddr(heap_io_accel_0_resp_bits_sizeAddr),
    .io_host_0_req_valid(heap_io_host_0_req_valid),
    .io_host_0_req_bits_allocDealloc(heap_io_host_0_req_bits_allocDealloc),
    .io_host_0_req_bits_sizeAddr(heap_io_host_0_req_bits_sizeAddr),
    .io_host_0_resp_valid(heap_io_host_0_resp_valid),
    .io_host_0_resp_bits_allocDealloc(heap_io_host_0_resp_bits_allocDealloc),
    .io_host_0_resp_bits_sizeAddr(heap_io_host_0_resp_bits_sizeAddr)
  );
  RegFile regs ( // @[Fringe.scala 116:20:@47072.4]
    .clock(regs_clock),
    .reset(regs_reset),
    .io_raddr(regs_io_raddr),
    .io_wen(regs_io_wen),
    .io_waddr(regs_io_waddr),
    .io_wdata(regs_io_wdata),
    .io_rdata(regs_io_rdata),
    .io_reset(regs_io_reset),
    .io_argIns_0(regs_io_argIns_0),
    .io_argIns_1(regs_io_argIns_1),
    .io_argIns_2(regs_io_argIns_2),
    .io_argOuts_0_valid(regs_io_argOuts_0_valid),
    .io_argOuts_0_bits(regs_io_argOuts_0_bits),
    .io_argOuts_1_valid(regs_io_argOuts_1_valid),
    .io_argOuts_1_bits(regs_io_argOuts_1_bits),
    .io_argOuts_2_valid(regs_io_argOuts_2_valid),
    .io_argOuts_2_bits(regs_io_argOuts_2_bits),
    .io_argOuts_3_valid(regs_io_argOuts_3_valid),
    .io_argOuts_3_bits(regs_io_argOuts_3_bits),
    .io_argOuts_4_valid(regs_io_argOuts_4_valid),
    .io_argOuts_4_bits(regs_io_argOuts_4_bits),
    .io_argOuts_5_valid(regs_io_argOuts_5_valid),
    .io_argOuts_5_bits(regs_io_argOuts_5_bits),
    .io_argOuts_6_valid(regs_io_argOuts_6_valid),
    .io_argOuts_6_bits(regs_io_argOuts_6_bits),
    .io_argOuts_7_valid(regs_io_argOuts_7_valid),
    .io_argOuts_7_bits(regs_io_argOuts_7_bits),
    .io_argOuts_8_valid(regs_io_argOuts_8_valid),
    .io_argOuts_8_bits(regs_io_argOuts_8_bits),
    .io_argOuts_9_valid(regs_io_argOuts_9_valid),
    .io_argOuts_9_bits(regs_io_argOuts_9_bits),
    .io_argOuts_10_valid(regs_io_argOuts_10_valid),
    .io_argOuts_10_bits(regs_io_argOuts_10_bits)
  );
  FringeCounter timeoutCtr ( // @[Fringe.scala 143:26:@49157.4]
    .clock(timeoutCtr_clock),
    .reset(timeoutCtr_reset),
    .io_enable(timeoutCtr_io_enable),
    .io_done(timeoutCtr_io_done)
  );
  Depulser depulser ( // @[Fringe.scala 153:24:@49175.4]
    .clock(depulser_clock),
    .reset(depulser_reset),
    .io_in(depulser_io_in),
    .io_rst(depulser_io_rst),
    .io_out(depulser_io_out)
  );
  assign _T_880 = regs_io_argIns_1; // @[:@49134.4 :@49135.4]
  assign curStatus_done = _T_880[0]; // @[Fringe.scala 133:45:@49136.4]
  assign curStatus_timeout = _T_880[1]; // @[Fringe.scala 133:45:@49138.4]
  assign curStatus_allocDealloc = _T_880[4:2]; // @[Fringe.scala 133:45:@49140.4]
  assign curStatus_sizeAddr = _T_880[63:5]; // @[Fringe.scala 133:45:@49142.4]
  assign _T_885 = regs_io_argIns_0[0]; // @[Fringe.scala 134:28:@49144.4]
  assign _T_889 = curStatus_done == 1'h0; // @[Fringe.scala 134:42:@49146.4]
  assign _T_890 = regs_io_argIns_0[1]; // @[Fringe.scala 135:27:@49148.4]
  assign _T_900 = ~ regs_io_argIns_0; // @[Fringe.scala 156:22:@49183.4]
  assign _T_908 = _T_907 ^ heap_io_host_0_req_valid; // @[package.scala 153:13:@49188.4]
  assign _T_909 = heap_io_host_0_req_valid & _T_908; // @[package.scala 153:8:@49189.4]
  assign _T_912 = _T_885 & depulser_io_out; // @[Fringe.scala 160:55:@49193.4]
  assign status_bits_done = depulser_io_out ? _T_912 : curStatus_done; // @[Fringe.scala 160:26:@49194.4]
  assign _T_915 = _T_885 & timeoutCtr_io_done; // @[Fringe.scala 161:58:@49197.4]
  assign status_bits_timeout = depulser_io_out ? _T_915 : curStatus_timeout; // @[Fringe.scala 161:29:@49198.4]
  assign _T_919 = heap_io_host_0_req_bits_allocDealloc ? 2'h1 : 2'h2; // @[Fringe.scala 162:57:@49200.4]
  assign _T_921 = heap_io_host_0_req_valid ? _T_919 : 2'h0; // @[Fringe.scala 162:34:@49201.4]
  assign _T_923 = heap_io_host_0_req_valid ? heap_io_host_0_req_bits_sizeAddr : 64'h0; // @[Fringe.scala 163:30:@49203.4]
  assign _T_924 = {status_bits_timeout,status_bits_done}; // @[Fringe.scala 171:37:@49206.4]
  assign status_bits_sizeAddr = _T_923[58:0]; // @[Fringe.scala 158:20:@49185.4 Fringe.scala 163:24:@49204.4]
  assign status_bits_allocDealloc = {{1'd0}, _T_921}; // @[Fringe.scala 158:20:@49185.4 Fringe.scala 162:28:@49202.4]
  assign _T_925 = {status_bits_sizeAddr,status_bits_allocDealloc}; // @[Fringe.scala 171:37:@49207.4]
  assign alloc = curStatus_allocDealloc == 3'h3; // @[Fringe.scala 202:38:@50519.4]
  assign dealloc = curStatus_allocDealloc == 3'h4; // @[Fringe.scala 203:40:@50520.4]
  assign _T_1429 = alloc | dealloc; // @[Fringe.scala 204:37:@50521.4]
  assign _T_1433 = _T_1432 ^ _T_1429; // @[package.scala 153:13:@50524.4]
  assign io_rdata = regs_io_rdata; // @[Fringe.scala 125:14:@49132.4]
  assign io_enable = _T_885 & _T_889; // @[Fringe.scala 136:13:@49152.4]
  assign io_reset = _T_890 | reset; // @[Fringe.scala 137:12:@49153.4]
  assign io_argIns_0 = regs_io_argIns_2; // @[Fringe.scala 151:51:@49174.4]
  assign io_heap_0_resp_valid = heap_io_accel_0_resp_valid; // @[Fringe.scala 108:17:@47068.4]
  assign io_heap_0_resp_bits_allocDealloc = heap_io_accel_0_resp_bits_allocDealloc; // @[Fringe.scala 108:17:@47067.4]
  assign io_heap_0_resp_bits_sizeAddr = heap_io_accel_0_resp_bits_sizeAddr; // @[Fringe.scala 108:17:@47066.4]
  assign heap_io_accel_0_req_valid = io_heap_0_req_valid; // @[Fringe.scala 108:17:@47071.4]
  assign heap_io_accel_0_req_bits_allocDealloc = io_heap_0_req_bits_allocDealloc; // @[Fringe.scala 108:17:@47070.4]
  assign heap_io_accel_0_req_bits_sizeAddr = io_heap_0_req_bits_sizeAddr; // @[Fringe.scala 108:17:@47069.4]
  assign heap_io_host_0_resp_valid = _T_1429 & _T_1433; // @[Fringe.scala 204:22:@50526.4]
  assign heap_io_host_0_resp_bits_allocDealloc = curStatus_allocDealloc == 3'h3; // @[Fringe.scala 205:34:@50527.4]
  assign heap_io_host_0_resp_bits_sizeAddr = {{5'd0}, curStatus_sizeAddr}; // @[Fringe.scala 206:30:@50528.4]
  assign regs_clock = clock; // @[:@47073.4]
  assign regs_reset = reset; // @[:@47074.4 Fringe.scala 139:14:@49156.4]
  assign regs_io_raddr = io_raddr; // @[Fringe.scala 118:17:@49128.4]
  assign regs_io_wen = io_wen; // @[Fringe.scala 120:15:@49130.4]
  assign regs_io_waddr = io_waddr; // @[Fringe.scala 119:17:@49129.4]
  assign regs_io_wdata = io_wdata; // @[Fringe.scala 121:17:@49131.4]
  assign regs_io_reset = _T_890 | reset; // @[Fringe.scala 138:17:@49154.4]
  assign regs_io_argOuts_0_valid = depulser_io_out | _T_909; // @[Fringe.scala 170:23:@49205.4]
  assign regs_io_argOuts_0_bits = {_T_925,_T_924}; // @[Fringe.scala 171:22:@49209.4]
  assign regs_io_argOuts_1_valid = io_argOuts_0_valid; // @[Fringe.scala 176:23:@49212.4]
  assign regs_io_argOuts_1_bits = io_argOuts_0_bits; // @[Fringe.scala 175:22:@49211.4]
  assign regs_io_argOuts_2_valid = io_argOuts_1_valid; // @[Fringe.scala 176:23:@49215.4]
  assign regs_io_argOuts_2_bits = io_argOuts_1_bits; // @[Fringe.scala 175:22:@49214.4]
  assign regs_io_argOuts_3_valid = io_argOuts_2_valid; // @[Fringe.scala 176:23:@49218.4]
  assign regs_io_argOuts_3_bits = io_argOuts_2_bits; // @[Fringe.scala 175:22:@49217.4]
  assign regs_io_argOuts_4_valid = io_argOuts_3_valid; // @[Fringe.scala 176:23:@49221.4]
  assign regs_io_argOuts_4_bits = io_argOuts_3_bits; // @[Fringe.scala 175:22:@49220.4]
  assign regs_io_argOuts_5_valid = io_argOuts_4_valid; // @[Fringe.scala 176:23:@49224.4]
  assign regs_io_argOuts_5_bits = io_argOuts_4_bits; // @[Fringe.scala 175:22:@49223.4]
  assign regs_io_argOuts_6_valid = io_argOuts_5_valid; // @[Fringe.scala 176:23:@49227.4]
  assign regs_io_argOuts_6_bits = io_argOuts_5_bits; // @[Fringe.scala 175:22:@49226.4]
  assign regs_io_argOuts_7_valid = io_argOuts_6_valid; // @[Fringe.scala 176:23:@49230.4]
  assign regs_io_argOuts_7_bits = io_argOuts_6_bits; // @[Fringe.scala 175:22:@49229.4]
  assign regs_io_argOuts_8_valid = io_argOuts_7_valid; // @[Fringe.scala 176:23:@49233.4]
  assign regs_io_argOuts_8_bits = io_argOuts_7_bits; // @[Fringe.scala 175:22:@49232.4]
  assign regs_io_argOuts_9_valid = io_argOuts_8_valid; // @[Fringe.scala 176:23:@49236.4]
  assign regs_io_argOuts_9_bits = io_argOuts_8_bits; // @[Fringe.scala 175:22:@49235.4]
  assign regs_io_argOuts_10_valid = io_argOuts_9_valid; // @[Fringe.scala 176:23:@49239.4]
  assign regs_io_argOuts_10_bits = io_argOuts_9_bits; // @[Fringe.scala 175:22:@49238.4]
  assign timeoutCtr_clock = clock; // @[:@49158.4]
  assign timeoutCtr_reset = reset; // @[:@49159.4]
  assign timeoutCtr_io_enable = _T_885 & _T_889; // @[Fringe.scala 149:24:@49173.4]
  assign depulser_clock = clock; // @[:@49176.4]
  assign depulser_reset = reset; // @[:@49177.4]
  assign depulser_io_in = io_done | timeoutCtr_io_done; // @[Fringe.scala 155:18:@49182.4]
  assign depulser_io_rst = _T_900[0]; // @[Fringe.scala 156:19:@49184.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_907 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1432 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_907 <= 1'h0;
    end else begin
      _T_907 <= heap_io_host_0_req_valid;
    end
    if (reset) begin
      _T_1432 <= 1'h0;
    end else begin
      _T_1432 <= _T_1429;
    end
  end
endmodule
module AXI4LiteToRFBridgeKCU1500( // @[:@50543.2]
  input         clock, // @[:@50544.4]
  input         reset, // @[:@50545.4]
  input  [31:0] io_S_AXI_AWADDR, // @[:@50546.4]
  input  [2:0]  io_S_AXI_AWPROT, // @[:@50546.4]
  input         io_S_AXI_AWVALID, // @[:@50546.4]
  output        io_S_AXI_AWREADY, // @[:@50546.4]
  input  [31:0] io_S_AXI_ARADDR, // @[:@50546.4]
  input  [2:0]  io_S_AXI_ARPROT, // @[:@50546.4]
  input         io_S_AXI_ARVALID, // @[:@50546.4]
  output        io_S_AXI_ARREADY, // @[:@50546.4]
  input  [31:0] io_S_AXI_WDATA, // @[:@50546.4]
  input  [3:0]  io_S_AXI_WSTRB, // @[:@50546.4]
  input         io_S_AXI_WVALID, // @[:@50546.4]
  output        io_S_AXI_WREADY, // @[:@50546.4]
  output [31:0] io_S_AXI_RDATA, // @[:@50546.4]
  output [1:0]  io_S_AXI_RRESP, // @[:@50546.4]
  output        io_S_AXI_RVALID, // @[:@50546.4]
  input         io_S_AXI_RREADY, // @[:@50546.4]
  output [1:0]  io_S_AXI_BRESP, // @[:@50546.4]
  output        io_S_AXI_BVALID, // @[:@50546.4]
  input         io_S_AXI_BREADY, // @[:@50546.4]
  output [31:0] io_raddr, // @[:@50546.4]
  output        io_wen, // @[:@50546.4]
  output [31:0] io_waddr, // @[:@50546.4]
  output [31:0] io_wdata, // @[:@50546.4]
  input  [31:0] io_rdata // @[:@50546.4]
);
  wire [31:0] d_rf_rdata; // @[AXI4LiteToRFBridge.scala 109:17:@50548.4]
  wire [31:0] d_rf_wdata; // @[AXI4LiteToRFBridge.scala 109:17:@50548.4]
  wire [31:0] d_rf_waddr; // @[AXI4LiteToRFBridge.scala 109:17:@50548.4]
  wire  d_rf_wen; // @[AXI4LiteToRFBridge.scala 109:17:@50548.4]
  wire [31:0] d_rf_raddr; // @[AXI4LiteToRFBridge.scala 109:17:@50548.4]
  wire  d_S_AXI_ARESETN; // @[AXI4LiteToRFBridge.scala 109:17:@50548.4]
  wire  d_S_AXI_ACLK; // @[AXI4LiteToRFBridge.scala 109:17:@50548.4]
  wire [31:0] d_S_AXI_AWADDR; // @[AXI4LiteToRFBridge.scala 109:17:@50548.4]
  wire [2:0] d_S_AXI_AWPROT; // @[AXI4LiteToRFBridge.scala 109:17:@50548.4]
  wire  d_S_AXI_AWVALID; // @[AXI4LiteToRFBridge.scala 109:17:@50548.4]
  wire  d_S_AXI_AWREADY; // @[AXI4LiteToRFBridge.scala 109:17:@50548.4]
  wire [31:0] d_S_AXI_ARADDR; // @[AXI4LiteToRFBridge.scala 109:17:@50548.4]
  wire [2:0] d_S_AXI_ARPROT; // @[AXI4LiteToRFBridge.scala 109:17:@50548.4]
  wire  d_S_AXI_ARVALID; // @[AXI4LiteToRFBridge.scala 109:17:@50548.4]
  wire  d_S_AXI_ARREADY; // @[AXI4LiteToRFBridge.scala 109:17:@50548.4]
  wire [31:0] d_S_AXI_WDATA; // @[AXI4LiteToRFBridge.scala 109:17:@50548.4]
  wire [3:0] d_S_AXI_WSTRB; // @[AXI4LiteToRFBridge.scala 109:17:@50548.4]
  wire  d_S_AXI_WVALID; // @[AXI4LiteToRFBridge.scala 109:17:@50548.4]
  wire  d_S_AXI_WREADY; // @[AXI4LiteToRFBridge.scala 109:17:@50548.4]
  wire [31:0] d_S_AXI_RDATA; // @[AXI4LiteToRFBridge.scala 109:17:@50548.4]
  wire [1:0] d_S_AXI_RRESP; // @[AXI4LiteToRFBridge.scala 109:17:@50548.4]
  wire  d_S_AXI_RVALID; // @[AXI4LiteToRFBridge.scala 109:17:@50548.4]
  wire  d_S_AXI_RREADY; // @[AXI4LiteToRFBridge.scala 109:17:@50548.4]
  wire [1:0] d_S_AXI_BRESP; // @[AXI4LiteToRFBridge.scala 109:17:@50548.4]
  wire  d_S_AXI_BVALID; // @[AXI4LiteToRFBridge.scala 109:17:@50548.4]
  wire  d_S_AXI_BREADY; // @[AXI4LiteToRFBridge.scala 109:17:@50548.4]
  AXI4LiteToRFBridgeVerilog d ( // @[AXI4LiteToRFBridge.scala 109:17:@50548.4]
    .rf_rdata(d_rf_rdata),
    .rf_wdata(d_rf_wdata),
    .rf_waddr(d_rf_waddr),
    .rf_wen(d_rf_wen),
    .rf_raddr(d_rf_raddr),
    .S_AXI_ARESETN(d_S_AXI_ARESETN),
    .S_AXI_ACLK(d_S_AXI_ACLK),
    .S_AXI_AWADDR(d_S_AXI_AWADDR),
    .S_AXI_AWPROT(d_S_AXI_AWPROT),
    .S_AXI_AWVALID(d_S_AXI_AWVALID),
    .S_AXI_AWREADY(d_S_AXI_AWREADY),
    .S_AXI_ARADDR(d_S_AXI_ARADDR),
    .S_AXI_ARPROT(d_S_AXI_ARPROT),
    .S_AXI_ARVALID(d_S_AXI_ARVALID),
    .S_AXI_ARREADY(d_S_AXI_ARREADY),
    .S_AXI_WDATA(d_S_AXI_WDATA),
    .S_AXI_WSTRB(d_S_AXI_WSTRB),
    .S_AXI_WVALID(d_S_AXI_WVALID),
    .S_AXI_WREADY(d_S_AXI_WREADY),
    .S_AXI_RDATA(d_S_AXI_RDATA),
    .S_AXI_RRESP(d_S_AXI_RRESP),
    .S_AXI_RVALID(d_S_AXI_RVALID),
    .S_AXI_RREADY(d_S_AXI_RREADY),
    .S_AXI_BRESP(d_S_AXI_BRESP),
    .S_AXI_BVALID(d_S_AXI_BVALID),
    .S_AXI_BREADY(d_S_AXI_BREADY)
  );
  assign io_S_AXI_AWREADY = d_S_AXI_AWREADY; // @[AXI4LiteToRFBridge.scala 111:14:@50572.4]
  assign io_S_AXI_ARREADY = d_S_AXI_ARREADY; // @[AXI4LiteToRFBridge.scala 111:14:@50568.4]
  assign io_S_AXI_WREADY = d_S_AXI_WREADY; // @[AXI4LiteToRFBridge.scala 111:14:@50564.4]
  assign io_S_AXI_RDATA = d_S_AXI_RDATA; // @[AXI4LiteToRFBridge.scala 111:14:@50563.4]
  assign io_S_AXI_RRESP = d_S_AXI_RRESP; // @[AXI4LiteToRFBridge.scala 111:14:@50562.4]
  assign io_S_AXI_RVALID = d_S_AXI_RVALID; // @[AXI4LiteToRFBridge.scala 111:14:@50561.4]
  assign io_S_AXI_BRESP = d_S_AXI_BRESP; // @[AXI4LiteToRFBridge.scala 111:14:@50559.4]
  assign io_S_AXI_BVALID = d_S_AXI_BVALID; // @[AXI4LiteToRFBridge.scala 111:14:@50558.4]
  assign io_raddr = d_rf_raddr; // @[AXI4LiteToRFBridge.scala 115:12:@50580.4]
  assign io_wen = d_rf_wen; // @[AXI4LiteToRFBridge.scala 118:12:@50583.4]
  assign io_waddr = d_rf_waddr; // @[AXI4LiteToRFBridge.scala 116:12:@50581.4]
  assign io_wdata = d_rf_wdata; // @[AXI4LiteToRFBridge.scala 117:12:@50582.4]
  assign d_rf_rdata = io_rdata; // @[AXI4LiteToRFBridge.scala 119:17:@50584.4]
  assign d_S_AXI_ARESETN = ~ reset; // @[AXI4LiteToRFBridge.scala 113:22:@50579.4]
  assign d_S_AXI_ACLK = clock; // @[AXI4LiteToRFBridge.scala 112:19:@50576.4]
  assign d_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[AXI4LiteToRFBridge.scala 111:14:@50575.4]
  assign d_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[AXI4LiteToRFBridge.scala 111:14:@50574.4]
  assign d_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[AXI4LiteToRFBridge.scala 111:14:@50573.4]
  assign d_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[AXI4LiteToRFBridge.scala 111:14:@50571.4]
  assign d_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[AXI4LiteToRFBridge.scala 111:14:@50570.4]
  assign d_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[AXI4LiteToRFBridge.scala 111:14:@50569.4]
  assign d_S_AXI_WDATA = io_S_AXI_WDATA; // @[AXI4LiteToRFBridge.scala 111:14:@50567.4]
  assign d_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[AXI4LiteToRFBridge.scala 111:14:@50566.4]
  assign d_S_AXI_WVALID = io_S_AXI_WVALID; // @[AXI4LiteToRFBridge.scala 111:14:@50565.4]
  assign d_S_AXI_RREADY = io_S_AXI_RREADY; // @[AXI4LiteToRFBridge.scala 111:14:@50560.4]
  assign d_S_AXI_BREADY = io_S_AXI_BREADY; // @[AXI4LiteToRFBridge.scala 111:14:@50557.4]
endmodule
module MAGToAXI4Bridge( // @[:@50586.2]
  output [7:0] io_M_AXI_AWLEN, // @[:@50589.4]
  output [7:0] io_M_AXI_ARLEN // @[:@50589.4]
);
  wire [32:0] _T_218; // @[MAGToAXI4Bridge.scala 27:29:@50746.4]
  wire [32:0] _T_219; // @[MAGToAXI4Bridge.scala 27:29:@50747.4]
  wire [31:0] _T_220; // @[MAGToAXI4Bridge.scala 27:29:@50748.4]
  assign _T_218 = 32'h0 - 32'h1; // @[MAGToAXI4Bridge.scala 27:29:@50746.4]
  assign _T_219 = $unsigned(_T_218); // @[MAGToAXI4Bridge.scala 27:29:@50747.4]
  assign _T_220 = _T_219[31:0]; // @[MAGToAXI4Bridge.scala 27:29:@50748.4]
  assign io_M_AXI_AWLEN = _T_220[7:0]; // @[MAGToAXI4Bridge.scala 41:21:@50766.4]
  assign io_M_AXI_ARLEN = _T_220[7:0]; // @[MAGToAXI4Bridge.scala 27:21:@50749.4]
endmodule
module FringeZynq( // @[:@50914.2]
  input         clock, // @[:@50915.4]
  input         reset, // @[:@50916.4]
  input  [31:0] io_S_AXI_AWADDR, // @[:@50917.4]
  input  [2:0]  io_S_AXI_AWPROT, // @[:@50917.4]
  input         io_S_AXI_AWVALID, // @[:@50917.4]
  output        io_S_AXI_AWREADY, // @[:@50917.4]
  input  [31:0] io_S_AXI_ARADDR, // @[:@50917.4]
  input  [2:0]  io_S_AXI_ARPROT, // @[:@50917.4]
  input         io_S_AXI_ARVALID, // @[:@50917.4]
  output        io_S_AXI_ARREADY, // @[:@50917.4]
  input  [31:0] io_S_AXI_WDATA, // @[:@50917.4]
  input  [3:0]  io_S_AXI_WSTRB, // @[:@50917.4]
  input         io_S_AXI_WVALID, // @[:@50917.4]
  output        io_S_AXI_WREADY, // @[:@50917.4]
  output [31:0] io_S_AXI_RDATA, // @[:@50917.4]
  output [1:0]  io_S_AXI_RRESP, // @[:@50917.4]
  output        io_S_AXI_RVALID, // @[:@50917.4]
  input         io_S_AXI_RREADY, // @[:@50917.4]
  output [1:0]  io_S_AXI_BRESP, // @[:@50917.4]
  output        io_S_AXI_BVALID, // @[:@50917.4]
  input         io_S_AXI_BREADY, // @[:@50917.4]
  output [7:0]  io_M_AXI_0_AWLEN, // @[:@50917.4]
  output [7:0]  io_M_AXI_0_ARLEN, // @[:@50917.4]
  output        io_enable, // @[:@50917.4]
  input         io_done, // @[:@50917.4]
  output        io_reset, // @[:@50917.4]
  output [63:0] io_argIns_0, // @[:@50917.4]
  input         io_argOuts_0_valid, // @[:@50917.4]
  input  [63:0] io_argOuts_0_bits, // @[:@50917.4]
  input         io_argOuts_1_valid, // @[:@50917.4]
  input  [63:0] io_argOuts_1_bits, // @[:@50917.4]
  input         io_argOuts_2_valid, // @[:@50917.4]
  input  [63:0] io_argOuts_2_bits, // @[:@50917.4]
  input         io_argOuts_3_valid, // @[:@50917.4]
  input  [63:0] io_argOuts_3_bits, // @[:@50917.4]
  input         io_argOuts_4_valid, // @[:@50917.4]
  input  [63:0] io_argOuts_4_bits, // @[:@50917.4]
  input         io_argOuts_5_valid, // @[:@50917.4]
  input  [63:0] io_argOuts_5_bits, // @[:@50917.4]
  input         io_argOuts_6_valid, // @[:@50917.4]
  input  [63:0] io_argOuts_6_bits, // @[:@50917.4]
  input         io_argOuts_7_valid, // @[:@50917.4]
  input  [63:0] io_argOuts_7_bits, // @[:@50917.4]
  input         io_argOuts_8_valid, // @[:@50917.4]
  input  [63:0] io_argOuts_8_bits, // @[:@50917.4]
  input         io_argOuts_9_valid, // @[:@50917.4]
  input  [63:0] io_argOuts_9_bits, // @[:@50917.4]
  input         io_heap_0_req_valid, // @[:@50917.4]
  input         io_heap_0_req_bits_allocDealloc, // @[:@50917.4]
  input  [63:0] io_heap_0_req_bits_sizeAddr, // @[:@50917.4]
  output        io_heap_0_resp_valid, // @[:@50917.4]
  output        io_heap_0_resp_bits_allocDealloc, // @[:@50917.4]
  output [63:0] io_heap_0_resp_bits_sizeAddr // @[:@50917.4]
);
  wire  fringeCommon_clock; // @[FringeZynq.scala 68:28:@51315.4]
  wire  fringeCommon_reset; // @[FringeZynq.scala 68:28:@51315.4]
  wire [31:0] fringeCommon_io_raddr; // @[FringeZynq.scala 68:28:@51315.4]
  wire  fringeCommon_io_wen; // @[FringeZynq.scala 68:28:@51315.4]
  wire [31:0] fringeCommon_io_waddr; // @[FringeZynq.scala 68:28:@51315.4]
  wire [63:0] fringeCommon_io_wdata; // @[FringeZynq.scala 68:28:@51315.4]
  wire [63:0] fringeCommon_io_rdata; // @[FringeZynq.scala 68:28:@51315.4]
  wire  fringeCommon_io_enable; // @[FringeZynq.scala 68:28:@51315.4]
  wire  fringeCommon_io_done; // @[FringeZynq.scala 68:28:@51315.4]
  wire  fringeCommon_io_reset; // @[FringeZynq.scala 68:28:@51315.4]
  wire [63:0] fringeCommon_io_argIns_0; // @[FringeZynq.scala 68:28:@51315.4]
  wire  fringeCommon_io_argOuts_0_valid; // @[FringeZynq.scala 68:28:@51315.4]
  wire [63:0] fringeCommon_io_argOuts_0_bits; // @[FringeZynq.scala 68:28:@51315.4]
  wire  fringeCommon_io_argOuts_1_valid; // @[FringeZynq.scala 68:28:@51315.4]
  wire [63:0] fringeCommon_io_argOuts_1_bits; // @[FringeZynq.scala 68:28:@51315.4]
  wire  fringeCommon_io_argOuts_2_valid; // @[FringeZynq.scala 68:28:@51315.4]
  wire [63:0] fringeCommon_io_argOuts_2_bits; // @[FringeZynq.scala 68:28:@51315.4]
  wire  fringeCommon_io_argOuts_3_valid; // @[FringeZynq.scala 68:28:@51315.4]
  wire [63:0] fringeCommon_io_argOuts_3_bits; // @[FringeZynq.scala 68:28:@51315.4]
  wire  fringeCommon_io_argOuts_4_valid; // @[FringeZynq.scala 68:28:@51315.4]
  wire [63:0] fringeCommon_io_argOuts_4_bits; // @[FringeZynq.scala 68:28:@51315.4]
  wire  fringeCommon_io_argOuts_5_valid; // @[FringeZynq.scala 68:28:@51315.4]
  wire [63:0] fringeCommon_io_argOuts_5_bits; // @[FringeZynq.scala 68:28:@51315.4]
  wire  fringeCommon_io_argOuts_6_valid; // @[FringeZynq.scala 68:28:@51315.4]
  wire [63:0] fringeCommon_io_argOuts_6_bits; // @[FringeZynq.scala 68:28:@51315.4]
  wire  fringeCommon_io_argOuts_7_valid; // @[FringeZynq.scala 68:28:@51315.4]
  wire [63:0] fringeCommon_io_argOuts_7_bits; // @[FringeZynq.scala 68:28:@51315.4]
  wire  fringeCommon_io_argOuts_8_valid; // @[FringeZynq.scala 68:28:@51315.4]
  wire [63:0] fringeCommon_io_argOuts_8_bits; // @[FringeZynq.scala 68:28:@51315.4]
  wire  fringeCommon_io_argOuts_9_valid; // @[FringeZynq.scala 68:28:@51315.4]
  wire [63:0] fringeCommon_io_argOuts_9_bits; // @[FringeZynq.scala 68:28:@51315.4]
  wire  fringeCommon_io_heap_0_req_valid; // @[FringeZynq.scala 68:28:@51315.4]
  wire  fringeCommon_io_heap_0_req_bits_allocDealloc; // @[FringeZynq.scala 68:28:@51315.4]
  wire [63:0] fringeCommon_io_heap_0_req_bits_sizeAddr; // @[FringeZynq.scala 68:28:@51315.4]
  wire  fringeCommon_io_heap_0_resp_valid; // @[FringeZynq.scala 68:28:@51315.4]
  wire  fringeCommon_io_heap_0_resp_bits_allocDealloc; // @[FringeZynq.scala 68:28:@51315.4]
  wire [63:0] fringeCommon_io_heap_0_resp_bits_sizeAddr; // @[FringeZynq.scala 68:28:@51315.4]
  wire  AXI4LiteToRFBridgeKCU1500_clock; // @[FringeZynq.scala 78:31:@51935.4]
  wire  AXI4LiteToRFBridgeKCU1500_reset; // @[FringeZynq.scala 78:31:@51935.4]
  wire [31:0] AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWADDR; // @[FringeZynq.scala 78:31:@51935.4]
  wire [2:0] AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWPROT; // @[FringeZynq.scala 78:31:@51935.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWVALID; // @[FringeZynq.scala 78:31:@51935.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWREADY; // @[FringeZynq.scala 78:31:@51935.4]
  wire [31:0] AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARADDR; // @[FringeZynq.scala 78:31:@51935.4]
  wire [2:0] AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARPROT; // @[FringeZynq.scala 78:31:@51935.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARVALID; // @[FringeZynq.scala 78:31:@51935.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARREADY; // @[FringeZynq.scala 78:31:@51935.4]
  wire [31:0] AXI4LiteToRFBridgeKCU1500_io_S_AXI_WDATA; // @[FringeZynq.scala 78:31:@51935.4]
  wire [3:0] AXI4LiteToRFBridgeKCU1500_io_S_AXI_WSTRB; // @[FringeZynq.scala 78:31:@51935.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_WVALID; // @[FringeZynq.scala 78:31:@51935.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_WREADY; // @[FringeZynq.scala 78:31:@51935.4]
  wire [31:0] AXI4LiteToRFBridgeKCU1500_io_S_AXI_RDATA; // @[FringeZynq.scala 78:31:@51935.4]
  wire [1:0] AXI4LiteToRFBridgeKCU1500_io_S_AXI_RRESP; // @[FringeZynq.scala 78:31:@51935.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_RVALID; // @[FringeZynq.scala 78:31:@51935.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_RREADY; // @[FringeZynq.scala 78:31:@51935.4]
  wire [1:0] AXI4LiteToRFBridgeKCU1500_io_S_AXI_BRESP; // @[FringeZynq.scala 78:31:@51935.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_BVALID; // @[FringeZynq.scala 78:31:@51935.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_S_AXI_BREADY; // @[FringeZynq.scala 78:31:@51935.4]
  wire [31:0] AXI4LiteToRFBridgeKCU1500_io_raddr; // @[FringeZynq.scala 78:31:@51935.4]
  wire  AXI4LiteToRFBridgeKCU1500_io_wen; // @[FringeZynq.scala 78:31:@51935.4]
  wire [31:0] AXI4LiteToRFBridgeKCU1500_io_waddr; // @[FringeZynq.scala 78:31:@51935.4]
  wire [31:0] AXI4LiteToRFBridgeKCU1500_io_wdata; // @[FringeZynq.scala 78:31:@51935.4]
  wire [31:0] AXI4LiteToRFBridgeKCU1500_io_rdata; // @[FringeZynq.scala 78:31:@51935.4]
  wire [7:0] MAGToAXI4Bridge_io_M_AXI_AWLEN; // @[FringeZynq.scala 130:27:@52128.4]
  wire [7:0] MAGToAXI4Bridge_io_M_AXI_ARLEN; // @[FringeZynq.scala 130:27:@52128.4]
  Fringe fringeCommon ( // @[FringeZynq.scala 68:28:@51315.4]
    .clock(fringeCommon_clock),
    .reset(fringeCommon_reset),
    .io_raddr(fringeCommon_io_raddr),
    .io_wen(fringeCommon_io_wen),
    .io_waddr(fringeCommon_io_waddr),
    .io_wdata(fringeCommon_io_wdata),
    .io_rdata(fringeCommon_io_rdata),
    .io_enable(fringeCommon_io_enable),
    .io_done(fringeCommon_io_done),
    .io_reset(fringeCommon_io_reset),
    .io_argIns_0(fringeCommon_io_argIns_0),
    .io_argOuts_0_valid(fringeCommon_io_argOuts_0_valid),
    .io_argOuts_0_bits(fringeCommon_io_argOuts_0_bits),
    .io_argOuts_1_valid(fringeCommon_io_argOuts_1_valid),
    .io_argOuts_1_bits(fringeCommon_io_argOuts_1_bits),
    .io_argOuts_2_valid(fringeCommon_io_argOuts_2_valid),
    .io_argOuts_2_bits(fringeCommon_io_argOuts_2_bits),
    .io_argOuts_3_valid(fringeCommon_io_argOuts_3_valid),
    .io_argOuts_3_bits(fringeCommon_io_argOuts_3_bits),
    .io_argOuts_4_valid(fringeCommon_io_argOuts_4_valid),
    .io_argOuts_4_bits(fringeCommon_io_argOuts_4_bits),
    .io_argOuts_5_valid(fringeCommon_io_argOuts_5_valid),
    .io_argOuts_5_bits(fringeCommon_io_argOuts_5_bits),
    .io_argOuts_6_valid(fringeCommon_io_argOuts_6_valid),
    .io_argOuts_6_bits(fringeCommon_io_argOuts_6_bits),
    .io_argOuts_7_valid(fringeCommon_io_argOuts_7_valid),
    .io_argOuts_7_bits(fringeCommon_io_argOuts_7_bits),
    .io_argOuts_8_valid(fringeCommon_io_argOuts_8_valid),
    .io_argOuts_8_bits(fringeCommon_io_argOuts_8_bits),
    .io_argOuts_9_valid(fringeCommon_io_argOuts_9_valid),
    .io_argOuts_9_bits(fringeCommon_io_argOuts_9_bits),
    .io_heap_0_req_valid(fringeCommon_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(fringeCommon_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(fringeCommon_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(fringeCommon_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(fringeCommon_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(fringeCommon_io_heap_0_resp_bits_sizeAddr)
  );
  AXI4LiteToRFBridgeKCU1500 AXI4LiteToRFBridgeKCU1500 ( // @[FringeZynq.scala 78:31:@51935.4]
    .clock(AXI4LiteToRFBridgeKCU1500_clock),
    .reset(AXI4LiteToRFBridgeKCU1500_reset),
    .io_S_AXI_AWADDR(AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWADDR),
    .io_S_AXI_AWPROT(AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWPROT),
    .io_S_AXI_AWVALID(AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWVALID),
    .io_S_AXI_AWREADY(AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWREADY),
    .io_S_AXI_ARADDR(AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARADDR),
    .io_S_AXI_ARPROT(AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARPROT),
    .io_S_AXI_ARVALID(AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARVALID),
    .io_S_AXI_ARREADY(AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARREADY),
    .io_S_AXI_WDATA(AXI4LiteToRFBridgeKCU1500_io_S_AXI_WDATA),
    .io_S_AXI_WSTRB(AXI4LiteToRFBridgeKCU1500_io_S_AXI_WSTRB),
    .io_S_AXI_WVALID(AXI4LiteToRFBridgeKCU1500_io_S_AXI_WVALID),
    .io_S_AXI_WREADY(AXI4LiteToRFBridgeKCU1500_io_S_AXI_WREADY),
    .io_S_AXI_RDATA(AXI4LiteToRFBridgeKCU1500_io_S_AXI_RDATA),
    .io_S_AXI_RRESP(AXI4LiteToRFBridgeKCU1500_io_S_AXI_RRESP),
    .io_S_AXI_RVALID(AXI4LiteToRFBridgeKCU1500_io_S_AXI_RVALID),
    .io_S_AXI_RREADY(AXI4LiteToRFBridgeKCU1500_io_S_AXI_RREADY),
    .io_S_AXI_BRESP(AXI4LiteToRFBridgeKCU1500_io_S_AXI_BRESP),
    .io_S_AXI_BVALID(AXI4LiteToRFBridgeKCU1500_io_S_AXI_BVALID),
    .io_S_AXI_BREADY(AXI4LiteToRFBridgeKCU1500_io_S_AXI_BREADY),
    .io_raddr(AXI4LiteToRFBridgeKCU1500_io_raddr),
    .io_wen(AXI4LiteToRFBridgeKCU1500_io_wen),
    .io_waddr(AXI4LiteToRFBridgeKCU1500_io_waddr),
    .io_wdata(AXI4LiteToRFBridgeKCU1500_io_wdata),
    .io_rdata(AXI4LiteToRFBridgeKCU1500_io_rdata)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge ( // @[FringeZynq.scala 130:27:@52128.4]
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_io_M_AXI_AWLEN),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_io_M_AXI_ARLEN)
  );
  assign io_S_AXI_AWREADY = AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWREADY; // @[FringeZynq.scala 79:28:@51953.4]
  assign io_S_AXI_ARREADY = AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARREADY; // @[FringeZynq.scala 79:28:@51949.4]
  assign io_S_AXI_WREADY = AXI4LiteToRFBridgeKCU1500_io_S_AXI_WREADY; // @[FringeZynq.scala 79:28:@51945.4]
  assign io_S_AXI_RDATA = AXI4LiteToRFBridgeKCU1500_io_S_AXI_RDATA; // @[FringeZynq.scala 79:28:@51944.4]
  assign io_S_AXI_RRESP = AXI4LiteToRFBridgeKCU1500_io_S_AXI_RRESP; // @[FringeZynq.scala 79:28:@51943.4]
  assign io_S_AXI_RVALID = AXI4LiteToRFBridgeKCU1500_io_S_AXI_RVALID; // @[FringeZynq.scala 79:28:@51942.4]
  assign io_S_AXI_BRESP = AXI4LiteToRFBridgeKCU1500_io_S_AXI_BRESP; // @[FringeZynq.scala 79:28:@51940.4]
  assign io_S_AXI_BVALID = AXI4LiteToRFBridgeKCU1500_io_S_AXI_BVALID; // @[FringeZynq.scala 79:28:@51939.4]
  assign io_M_AXI_0_AWLEN = MAGToAXI4Bridge_io_M_AXI_AWLEN; // @[FringeZynq.scala 132:10:@52280.4]
  assign io_M_AXI_0_ARLEN = MAGToAXI4Bridge_io_M_AXI_ARLEN; // @[FringeZynq.scala 132:10:@52268.4]
  assign io_enable = fringeCommon_io_enable; // @[FringeZynq.scala 114:13:@51965.4]
  assign io_reset = fringeCommon_io_reset; // @[FringeZynq.scala 118:12:@51969.4]
  assign io_argIns_0 = fringeCommon_io_argIns_0; // @[FringeZynq.scala 120:13:@51970.4]
  assign io_heap_0_resp_valid = fringeCommon_io_heap_0_resp_valid; // @[FringeZynq.scala 126:11:@52124.4]
  assign io_heap_0_resp_bits_allocDealloc = fringeCommon_io_heap_0_resp_bits_allocDealloc; // @[FringeZynq.scala 126:11:@52123.4]
  assign io_heap_0_resp_bits_sizeAddr = fringeCommon_io_heap_0_resp_bits_sizeAddr; // @[FringeZynq.scala 126:11:@52122.4]
  assign fringeCommon_clock = clock; // @[:@51316.4]
  assign fringeCommon_reset = reset; // @[:@51317.4 FringeZynq.scala 81:24:@51958.4 FringeZynq.scala 116:22:@51968.4]
  assign fringeCommon_io_raddr = AXI4LiteToRFBridgeKCU1500_io_raddr; // @[FringeZynq.scala 82:27:@51959.4]
  assign fringeCommon_io_wen = AXI4LiteToRFBridgeKCU1500_io_wen; // @[FringeZynq.scala 83:27:@51960.4]
  assign fringeCommon_io_waddr = AXI4LiteToRFBridgeKCU1500_io_waddr; // @[FringeZynq.scala 84:27:@51961.4]
  assign fringeCommon_io_wdata = {{32'd0}, AXI4LiteToRFBridgeKCU1500_io_wdata}; // @[FringeZynq.scala 85:27:@51962.4]
  assign fringeCommon_io_done = io_done; // @[FringeZynq.scala 115:24:@51966.4]
  assign fringeCommon_io_argOuts_0_valid = io_argOuts_0_valid; // @[FringeZynq.scala 121:27:@51972.4]
  assign fringeCommon_io_argOuts_0_bits = io_argOuts_0_bits; // @[FringeZynq.scala 121:27:@51971.4]
  assign fringeCommon_io_argOuts_1_valid = io_argOuts_1_valid; // @[FringeZynq.scala 121:27:@51975.4]
  assign fringeCommon_io_argOuts_1_bits = io_argOuts_1_bits; // @[FringeZynq.scala 121:27:@51974.4]
  assign fringeCommon_io_argOuts_2_valid = io_argOuts_2_valid; // @[FringeZynq.scala 121:27:@51978.4]
  assign fringeCommon_io_argOuts_2_bits = io_argOuts_2_bits; // @[FringeZynq.scala 121:27:@51977.4]
  assign fringeCommon_io_argOuts_3_valid = io_argOuts_3_valid; // @[FringeZynq.scala 121:27:@51981.4]
  assign fringeCommon_io_argOuts_3_bits = io_argOuts_3_bits; // @[FringeZynq.scala 121:27:@51980.4]
  assign fringeCommon_io_argOuts_4_valid = io_argOuts_4_valid; // @[FringeZynq.scala 121:27:@51984.4]
  assign fringeCommon_io_argOuts_4_bits = io_argOuts_4_bits; // @[FringeZynq.scala 121:27:@51983.4]
  assign fringeCommon_io_argOuts_5_valid = io_argOuts_5_valid; // @[FringeZynq.scala 121:27:@51987.4]
  assign fringeCommon_io_argOuts_5_bits = io_argOuts_5_bits; // @[FringeZynq.scala 121:27:@51986.4]
  assign fringeCommon_io_argOuts_6_valid = io_argOuts_6_valid; // @[FringeZynq.scala 121:27:@51990.4]
  assign fringeCommon_io_argOuts_6_bits = io_argOuts_6_bits; // @[FringeZynq.scala 121:27:@51989.4]
  assign fringeCommon_io_argOuts_7_valid = io_argOuts_7_valid; // @[FringeZynq.scala 121:27:@51993.4]
  assign fringeCommon_io_argOuts_7_bits = io_argOuts_7_bits; // @[FringeZynq.scala 121:27:@51992.4]
  assign fringeCommon_io_argOuts_8_valid = io_argOuts_8_valid; // @[FringeZynq.scala 121:27:@51996.4]
  assign fringeCommon_io_argOuts_8_bits = io_argOuts_8_bits; // @[FringeZynq.scala 121:27:@51995.4]
  assign fringeCommon_io_argOuts_9_valid = io_argOuts_9_valid; // @[FringeZynq.scala 121:27:@51999.4]
  assign fringeCommon_io_argOuts_9_bits = io_argOuts_9_bits; // @[FringeZynq.scala 121:27:@51998.4]
  assign fringeCommon_io_heap_0_req_valid = io_heap_0_req_valid; // @[FringeZynq.scala 126:11:@52127.4]
  assign fringeCommon_io_heap_0_req_bits_allocDealloc = io_heap_0_req_bits_allocDealloc; // @[FringeZynq.scala 126:11:@52126.4]
  assign fringeCommon_io_heap_0_req_bits_sizeAddr = io_heap_0_req_bits_sizeAddr; // @[FringeZynq.scala 126:11:@52125.4]
  assign AXI4LiteToRFBridgeKCU1500_clock = clock; // @[:@51936.4]
  assign AXI4LiteToRFBridgeKCU1500_reset = reset; // @[:@51937.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[FringeZynq.scala 79:28:@51956.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[FringeZynq.scala 79:28:@51955.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[FringeZynq.scala 79:28:@51954.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[FringeZynq.scala 79:28:@51952.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[FringeZynq.scala 79:28:@51951.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[FringeZynq.scala 79:28:@51950.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_WDATA = io_S_AXI_WDATA; // @[FringeZynq.scala 79:28:@51948.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[FringeZynq.scala 79:28:@51947.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_WVALID = io_S_AXI_WVALID; // @[FringeZynq.scala 79:28:@51946.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_RREADY = io_S_AXI_RREADY; // @[FringeZynq.scala 79:28:@51941.4]
  assign AXI4LiteToRFBridgeKCU1500_io_S_AXI_BREADY = io_S_AXI_BREADY; // @[FringeZynq.scala 79:28:@51938.4]
  assign AXI4LiteToRFBridgeKCU1500_io_rdata = fringeCommon_io_rdata[31:0]; // @[FringeZynq.scala 86:28:@51963.4]
endmodule
module SpatialIP( // @[:@52285.2]
  input          clock, // @[:@52286.4]
  input          reset, // @[:@52287.4]
  input          io_raddr, // @[:@52288.4]
  input          io_wen, // @[:@52288.4]
  input          io_waddr, // @[:@52288.4]
  input          io_wdata, // @[:@52288.4]
  output         io_rdata, // @[:@52288.4]
  input  [31:0]  io_S_AXI_AWADDR, // @[:@52288.4]
  input  [2:0]   io_S_AXI_AWPROT, // @[:@52288.4]
  input          io_S_AXI_AWVALID, // @[:@52288.4]
  output         io_S_AXI_AWREADY, // @[:@52288.4]
  input  [31:0]  io_S_AXI_ARADDR, // @[:@52288.4]
  input  [2:0]   io_S_AXI_ARPROT, // @[:@52288.4]
  input          io_S_AXI_ARVALID, // @[:@52288.4]
  output         io_S_AXI_ARREADY, // @[:@52288.4]
  input  [31:0]  io_S_AXI_WDATA, // @[:@52288.4]
  input  [3:0]   io_S_AXI_WSTRB, // @[:@52288.4]
  input          io_S_AXI_WVALID, // @[:@52288.4]
  output         io_S_AXI_WREADY, // @[:@52288.4]
  output [31:0]  io_S_AXI_RDATA, // @[:@52288.4]
  output [1:0]   io_S_AXI_RRESP, // @[:@52288.4]
  output         io_S_AXI_RVALID, // @[:@52288.4]
  input          io_S_AXI_RREADY, // @[:@52288.4]
  output [1:0]   io_S_AXI_BRESP, // @[:@52288.4]
  output         io_S_AXI_BVALID, // @[:@52288.4]
  input          io_S_AXI_BREADY, // @[:@52288.4]
  output [3:0]   io_M_AXI_0_AWID, // @[:@52288.4]
  output [3:0]   io_M_AXI_0_AWUSER, // @[:@52288.4]
  output [31:0]  io_M_AXI_0_AWADDR, // @[:@52288.4]
  output [7:0]   io_M_AXI_0_AWLEN, // @[:@52288.4]
  output [2:0]   io_M_AXI_0_AWSIZE, // @[:@52288.4]
  output [1:0]   io_M_AXI_0_AWBURST, // @[:@52288.4]
  output         io_M_AXI_0_AWLOCK, // @[:@52288.4]
  output [3:0]   io_M_AXI_0_AWCACHE, // @[:@52288.4]
  output [2:0]   io_M_AXI_0_AWPROT, // @[:@52288.4]
  output [3:0]   io_M_AXI_0_AWQOS, // @[:@52288.4]
  output         io_M_AXI_0_AWVALID, // @[:@52288.4]
  input          io_M_AXI_0_AWREADY, // @[:@52288.4]
  output [3:0]   io_M_AXI_0_ARID, // @[:@52288.4]
  output [3:0]   io_M_AXI_0_ARUSER, // @[:@52288.4]
  output [31:0]  io_M_AXI_0_ARADDR, // @[:@52288.4]
  output [7:0]   io_M_AXI_0_ARLEN, // @[:@52288.4]
  output [2:0]   io_M_AXI_0_ARSIZE, // @[:@52288.4]
  output [1:0]   io_M_AXI_0_ARBURST, // @[:@52288.4]
  output         io_M_AXI_0_ARLOCK, // @[:@52288.4]
  output [3:0]   io_M_AXI_0_ARCACHE, // @[:@52288.4]
  output [2:0]   io_M_AXI_0_ARPROT, // @[:@52288.4]
  output [3:0]   io_M_AXI_0_ARQOS, // @[:@52288.4]
  output         io_M_AXI_0_ARVALID, // @[:@52288.4]
  input          io_M_AXI_0_ARREADY, // @[:@52288.4]
  output [511:0] io_M_AXI_0_WDATA, // @[:@52288.4]
  output [63:0]  io_M_AXI_0_WSTRB, // @[:@52288.4]
  output         io_M_AXI_0_WLAST, // @[:@52288.4]
  output         io_M_AXI_0_WVALID, // @[:@52288.4]
  input          io_M_AXI_0_WREADY, // @[:@52288.4]
  input  [3:0]   io_M_AXI_0_RID, // @[:@52288.4]
  input  [31:0]  io_M_AXI_0_RUSER, // @[:@52288.4]
  input  [511:0] io_M_AXI_0_RDATA, // @[:@52288.4]
  input  [1:0]   io_M_AXI_0_RRESP, // @[:@52288.4]
  input          io_M_AXI_0_RLAST, // @[:@52288.4]
  input          io_M_AXI_0_RVALID, // @[:@52288.4]
  output         io_M_AXI_0_RREADY, // @[:@52288.4]
  input  [3:0]   io_M_AXI_0_BID, // @[:@52288.4]
  input  [3:0]   io_M_AXI_0_BUSER, // @[:@52288.4]
  input  [1:0]   io_M_AXI_0_BRESP, // @[:@52288.4]
  input          io_M_AXI_0_BVALID, // @[:@52288.4]
  output         io_M_AXI_0_BREADY, // @[:@52288.4]
  input          io_AXIS_IN_TVALID, // @[:@52288.4]
  output         io_AXIS_IN_TREADY, // @[:@52288.4]
  input  [511:0] io_AXIS_IN_TDATA, // @[:@52288.4]
  input  [63:0]  io_AXIS_IN_TSTRB, // @[:@52288.4]
  input  [63:0]  io_AXIS_IN_TKEEP, // @[:@52288.4]
  input          io_AXIS_IN_TLAST, // @[:@52288.4]
  input  [7:0]   io_AXIS_IN_TID, // @[:@52288.4]
  input  [7:0]   io_AXIS_IN_TDEST, // @[:@52288.4]
  input  [511:0] io_AXIS_IN_TUSER, // @[:@52288.4]
  output         io_AXIS_OUT_TVALID, // @[:@52288.4]
  input          io_AXIS_OUT_TREADY, // @[:@52288.4]
  output [511:0] io_AXIS_OUT_TDATA, // @[:@52288.4]
  output [63:0]  io_AXIS_OUT_TSTRB, // @[:@52288.4]
  output [63:0]  io_AXIS_OUT_TKEEP, // @[:@52288.4]
  output         io_AXIS_OUT_TLAST, // @[:@52288.4]
  output [7:0]   io_AXIS_OUT_TID, // @[:@52288.4]
  output [7:0]   io_AXIS_OUT_TDEST, // @[:@52288.4]
  output [511:0] io_AXIS_OUT_TUSER // @[:@52288.4]
);
  wire  accel_clock; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_reset; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_enable; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_done; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_reset; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_memStreams_loads_0_cmd_ready; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_memStreams_loads_0_cmd_valid; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_memStreams_loads_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_loads_0_cmd_bits_size; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_memStreams_loads_0_data_ready; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_memStreams_loads_0_data_valid; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_0; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_1; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_2; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_3; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_4; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_5; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_6; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_7; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_8; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_9; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_10; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_11; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_12; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_13; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_14; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_15; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_memStreams_stores_0_cmd_ready; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_memStreams_stores_0_cmd_valid; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_memStreams_stores_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_stores_0_cmd_bits_size; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_memStreams_stores_0_data_ready; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_memStreams_stores_0_data_valid; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_0; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_1; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_2; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_3; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_4; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_5; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_6; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_7; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_8; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_9; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_10; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_11; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_12; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_13; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_14; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_15; // @[Instantiator.scala 53:44:@52290.4]
  wire [15:0] accel_io_memStreams_stores_0_data_bits_wstrb; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_memStreams_stores_0_wresp_ready; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_memStreams_stores_0_wresp_valid; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_memStreams_stores_0_wresp_bits; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_memStreams_gathers_0_cmd_ready; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_memStreams_gathers_0_cmd_valid; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_0; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_1; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_2; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_3; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_4; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_5; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_6; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_7; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_8; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_9; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_10; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_11; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_12; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_13; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_14; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_15; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_memStreams_gathers_0_data_ready; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_memStreams_gathers_0_data_valid; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_0; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_1; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_2; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_3; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_4; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_5; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_6; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_7; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_8; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_9; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_10; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_11; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_12; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_13; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_14; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_15; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_memStreams_scatters_0_cmd_ready; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_memStreams_scatters_0_cmd_valid; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_0; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_1; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_2; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_3; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_4; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_5; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_6; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_7; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_8; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_9; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_10; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_11; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_12; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_13; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_14; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_15; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_memStreams_scatters_0_wresp_ready; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_memStreams_scatters_0_wresp_valid; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_memStreams_scatters_0_wresp_bits; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_axiStreamsIn_0_TVALID; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_axiStreamsIn_0_TREADY; // @[Instantiator.scala 53:44:@52290.4]
  wire [255:0] accel_io_axiStreamsIn_0_TDATA; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_axiStreamsIn_0_TSTRB; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_axiStreamsIn_0_TKEEP; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_axiStreamsIn_0_TLAST; // @[Instantiator.scala 53:44:@52290.4]
  wire [7:0] accel_io_axiStreamsIn_0_TID; // @[Instantiator.scala 53:44:@52290.4]
  wire [7:0] accel_io_axiStreamsIn_0_TDEST; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_axiStreamsIn_0_TUSER; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_axiStreamsOut_0_TVALID; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_axiStreamsOut_0_TREADY; // @[Instantiator.scala 53:44:@52290.4]
  wire [511:0] accel_io_axiStreamsOut_0_TDATA; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_axiStreamsOut_0_TSTRB; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_axiStreamsOut_0_TKEEP; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_axiStreamsOut_0_TLAST; // @[Instantiator.scala 53:44:@52290.4]
  wire [7:0] accel_io_axiStreamsOut_0_TID; // @[Instantiator.scala 53:44:@52290.4]
  wire [7:0] accel_io_axiStreamsOut_0_TDEST; // @[Instantiator.scala 53:44:@52290.4]
  wire [31:0] accel_io_axiStreamsOut_0_TUSER; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_heap_0_req_valid; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_heap_0_req_bits_allocDealloc; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_heap_0_req_bits_sizeAddr; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_heap_0_resp_valid; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_heap_0_resp_bits_allocDealloc; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_heap_0_resp_bits_sizeAddr; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_argIns_0; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_argOuts_0_port_ready; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_argOuts_0_port_valid; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_argOuts_0_port_bits; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_argOuts_0_echo; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_argOuts_1_port_ready; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_argOuts_1_port_valid; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_argOuts_1_port_bits; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_argOuts_1_echo; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_argOuts_2_port_ready; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_argOuts_2_port_valid; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_argOuts_2_port_bits; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_argOuts_2_echo; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_argOuts_3_port_ready; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_argOuts_3_port_valid; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_argOuts_3_port_bits; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_argOuts_3_echo; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_argOuts_4_port_ready; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_argOuts_4_port_valid; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_argOuts_4_port_bits; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_argOuts_4_echo; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_argOuts_5_port_ready; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_argOuts_5_port_valid; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_argOuts_5_port_bits; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_argOuts_5_echo; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_argOuts_6_port_ready; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_argOuts_6_port_valid; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_argOuts_6_port_bits; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_argOuts_6_echo; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_argOuts_7_port_ready; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_argOuts_7_port_valid; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_argOuts_7_port_bits; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_argOuts_7_echo; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_argOuts_8_port_ready; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_argOuts_8_port_valid; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_argOuts_8_port_bits; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_argOuts_8_echo; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_argOuts_9_port_ready; // @[Instantiator.scala 53:44:@52290.4]
  wire  accel_io_argOuts_9_port_valid; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_argOuts_9_port_bits; // @[Instantiator.scala 53:44:@52290.4]
  wire [63:0] accel_io_argOuts_9_echo; // @[Instantiator.scala 53:44:@52290.4]
  wire  FringeZynq_clock; // @[KCU1500.scala 21:24:@52482.4]
  wire  FringeZynq_reset; // @[KCU1500.scala 21:24:@52482.4]
  wire [31:0] FringeZynq_io_S_AXI_AWADDR; // @[KCU1500.scala 21:24:@52482.4]
  wire [2:0] FringeZynq_io_S_AXI_AWPROT; // @[KCU1500.scala 21:24:@52482.4]
  wire  FringeZynq_io_S_AXI_AWVALID; // @[KCU1500.scala 21:24:@52482.4]
  wire  FringeZynq_io_S_AXI_AWREADY; // @[KCU1500.scala 21:24:@52482.4]
  wire [31:0] FringeZynq_io_S_AXI_ARADDR; // @[KCU1500.scala 21:24:@52482.4]
  wire [2:0] FringeZynq_io_S_AXI_ARPROT; // @[KCU1500.scala 21:24:@52482.4]
  wire  FringeZynq_io_S_AXI_ARVALID; // @[KCU1500.scala 21:24:@52482.4]
  wire  FringeZynq_io_S_AXI_ARREADY; // @[KCU1500.scala 21:24:@52482.4]
  wire [31:0] FringeZynq_io_S_AXI_WDATA; // @[KCU1500.scala 21:24:@52482.4]
  wire [3:0] FringeZynq_io_S_AXI_WSTRB; // @[KCU1500.scala 21:24:@52482.4]
  wire  FringeZynq_io_S_AXI_WVALID; // @[KCU1500.scala 21:24:@52482.4]
  wire  FringeZynq_io_S_AXI_WREADY; // @[KCU1500.scala 21:24:@52482.4]
  wire [31:0] FringeZynq_io_S_AXI_RDATA; // @[KCU1500.scala 21:24:@52482.4]
  wire [1:0] FringeZynq_io_S_AXI_RRESP; // @[KCU1500.scala 21:24:@52482.4]
  wire  FringeZynq_io_S_AXI_RVALID; // @[KCU1500.scala 21:24:@52482.4]
  wire  FringeZynq_io_S_AXI_RREADY; // @[KCU1500.scala 21:24:@52482.4]
  wire [1:0] FringeZynq_io_S_AXI_BRESP; // @[KCU1500.scala 21:24:@52482.4]
  wire  FringeZynq_io_S_AXI_BVALID; // @[KCU1500.scala 21:24:@52482.4]
  wire  FringeZynq_io_S_AXI_BREADY; // @[KCU1500.scala 21:24:@52482.4]
  wire [7:0] FringeZynq_io_M_AXI_0_AWLEN; // @[KCU1500.scala 21:24:@52482.4]
  wire [7:0] FringeZynq_io_M_AXI_0_ARLEN; // @[KCU1500.scala 21:24:@52482.4]
  wire  FringeZynq_io_enable; // @[KCU1500.scala 21:24:@52482.4]
  wire  FringeZynq_io_done; // @[KCU1500.scala 21:24:@52482.4]
  wire  FringeZynq_io_reset; // @[KCU1500.scala 21:24:@52482.4]
  wire [63:0] FringeZynq_io_argIns_0; // @[KCU1500.scala 21:24:@52482.4]
  wire  FringeZynq_io_argOuts_0_valid; // @[KCU1500.scala 21:24:@52482.4]
  wire [63:0] FringeZynq_io_argOuts_0_bits; // @[KCU1500.scala 21:24:@52482.4]
  wire  FringeZynq_io_argOuts_1_valid; // @[KCU1500.scala 21:24:@52482.4]
  wire [63:0] FringeZynq_io_argOuts_1_bits; // @[KCU1500.scala 21:24:@52482.4]
  wire  FringeZynq_io_argOuts_2_valid; // @[KCU1500.scala 21:24:@52482.4]
  wire [63:0] FringeZynq_io_argOuts_2_bits; // @[KCU1500.scala 21:24:@52482.4]
  wire  FringeZynq_io_argOuts_3_valid; // @[KCU1500.scala 21:24:@52482.4]
  wire [63:0] FringeZynq_io_argOuts_3_bits; // @[KCU1500.scala 21:24:@52482.4]
  wire  FringeZynq_io_argOuts_4_valid; // @[KCU1500.scala 21:24:@52482.4]
  wire [63:0] FringeZynq_io_argOuts_4_bits; // @[KCU1500.scala 21:24:@52482.4]
  wire  FringeZynq_io_argOuts_5_valid; // @[KCU1500.scala 21:24:@52482.4]
  wire [63:0] FringeZynq_io_argOuts_5_bits; // @[KCU1500.scala 21:24:@52482.4]
  wire  FringeZynq_io_argOuts_6_valid; // @[KCU1500.scala 21:24:@52482.4]
  wire [63:0] FringeZynq_io_argOuts_6_bits; // @[KCU1500.scala 21:24:@52482.4]
  wire  FringeZynq_io_argOuts_7_valid; // @[KCU1500.scala 21:24:@52482.4]
  wire [63:0] FringeZynq_io_argOuts_7_bits; // @[KCU1500.scala 21:24:@52482.4]
  wire  FringeZynq_io_argOuts_8_valid; // @[KCU1500.scala 21:24:@52482.4]
  wire [63:0] FringeZynq_io_argOuts_8_bits; // @[KCU1500.scala 21:24:@52482.4]
  wire  FringeZynq_io_argOuts_9_valid; // @[KCU1500.scala 21:24:@52482.4]
  wire [63:0] FringeZynq_io_argOuts_9_bits; // @[KCU1500.scala 21:24:@52482.4]
  wire  FringeZynq_io_heap_0_req_valid; // @[KCU1500.scala 21:24:@52482.4]
  wire  FringeZynq_io_heap_0_req_bits_allocDealloc; // @[KCU1500.scala 21:24:@52482.4]
  wire [63:0] FringeZynq_io_heap_0_req_bits_sizeAddr; // @[KCU1500.scala 21:24:@52482.4]
  wire  FringeZynq_io_heap_0_resp_valid; // @[KCU1500.scala 21:24:@52482.4]
  wire  FringeZynq_io_heap_0_resp_bits_allocDealloc; // @[KCU1500.scala 21:24:@52482.4]
  wire [63:0] FringeZynq_io_heap_0_resp_bits_sizeAddr; // @[KCU1500.scala 21:24:@52482.4]
  AccelUnit accel ( // @[Instantiator.scala 53:44:@52290.4]
    .clock(accel_clock),
    .reset(accel_reset),
    .io_enable(accel_io_enable),
    .io_done(accel_io_done),
    .io_reset(accel_io_reset),
    .io_memStreams_loads_0_cmd_ready(accel_io_memStreams_loads_0_cmd_ready),
    .io_memStreams_loads_0_cmd_valid(accel_io_memStreams_loads_0_cmd_valid),
    .io_memStreams_loads_0_cmd_bits_addr(accel_io_memStreams_loads_0_cmd_bits_addr),
    .io_memStreams_loads_0_cmd_bits_size(accel_io_memStreams_loads_0_cmd_bits_size),
    .io_memStreams_loads_0_data_ready(accel_io_memStreams_loads_0_data_ready),
    .io_memStreams_loads_0_data_valid(accel_io_memStreams_loads_0_data_valid),
    .io_memStreams_loads_0_data_bits_rdata_0(accel_io_memStreams_loads_0_data_bits_rdata_0),
    .io_memStreams_loads_0_data_bits_rdata_1(accel_io_memStreams_loads_0_data_bits_rdata_1),
    .io_memStreams_loads_0_data_bits_rdata_2(accel_io_memStreams_loads_0_data_bits_rdata_2),
    .io_memStreams_loads_0_data_bits_rdata_3(accel_io_memStreams_loads_0_data_bits_rdata_3),
    .io_memStreams_loads_0_data_bits_rdata_4(accel_io_memStreams_loads_0_data_bits_rdata_4),
    .io_memStreams_loads_0_data_bits_rdata_5(accel_io_memStreams_loads_0_data_bits_rdata_5),
    .io_memStreams_loads_0_data_bits_rdata_6(accel_io_memStreams_loads_0_data_bits_rdata_6),
    .io_memStreams_loads_0_data_bits_rdata_7(accel_io_memStreams_loads_0_data_bits_rdata_7),
    .io_memStreams_loads_0_data_bits_rdata_8(accel_io_memStreams_loads_0_data_bits_rdata_8),
    .io_memStreams_loads_0_data_bits_rdata_9(accel_io_memStreams_loads_0_data_bits_rdata_9),
    .io_memStreams_loads_0_data_bits_rdata_10(accel_io_memStreams_loads_0_data_bits_rdata_10),
    .io_memStreams_loads_0_data_bits_rdata_11(accel_io_memStreams_loads_0_data_bits_rdata_11),
    .io_memStreams_loads_0_data_bits_rdata_12(accel_io_memStreams_loads_0_data_bits_rdata_12),
    .io_memStreams_loads_0_data_bits_rdata_13(accel_io_memStreams_loads_0_data_bits_rdata_13),
    .io_memStreams_loads_0_data_bits_rdata_14(accel_io_memStreams_loads_0_data_bits_rdata_14),
    .io_memStreams_loads_0_data_bits_rdata_15(accel_io_memStreams_loads_0_data_bits_rdata_15),
    .io_memStreams_stores_0_cmd_ready(accel_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(accel_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(accel_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(accel_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(accel_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(accel_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(accel_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wdata_1(accel_io_memStreams_stores_0_data_bits_wdata_1),
    .io_memStreams_stores_0_data_bits_wdata_2(accel_io_memStreams_stores_0_data_bits_wdata_2),
    .io_memStreams_stores_0_data_bits_wdata_3(accel_io_memStreams_stores_0_data_bits_wdata_3),
    .io_memStreams_stores_0_data_bits_wdata_4(accel_io_memStreams_stores_0_data_bits_wdata_4),
    .io_memStreams_stores_0_data_bits_wdata_5(accel_io_memStreams_stores_0_data_bits_wdata_5),
    .io_memStreams_stores_0_data_bits_wdata_6(accel_io_memStreams_stores_0_data_bits_wdata_6),
    .io_memStreams_stores_0_data_bits_wdata_7(accel_io_memStreams_stores_0_data_bits_wdata_7),
    .io_memStreams_stores_0_data_bits_wdata_8(accel_io_memStreams_stores_0_data_bits_wdata_8),
    .io_memStreams_stores_0_data_bits_wdata_9(accel_io_memStreams_stores_0_data_bits_wdata_9),
    .io_memStreams_stores_0_data_bits_wdata_10(accel_io_memStreams_stores_0_data_bits_wdata_10),
    .io_memStreams_stores_0_data_bits_wdata_11(accel_io_memStreams_stores_0_data_bits_wdata_11),
    .io_memStreams_stores_0_data_bits_wdata_12(accel_io_memStreams_stores_0_data_bits_wdata_12),
    .io_memStreams_stores_0_data_bits_wdata_13(accel_io_memStreams_stores_0_data_bits_wdata_13),
    .io_memStreams_stores_0_data_bits_wdata_14(accel_io_memStreams_stores_0_data_bits_wdata_14),
    .io_memStreams_stores_0_data_bits_wdata_15(accel_io_memStreams_stores_0_data_bits_wdata_15),
    .io_memStreams_stores_0_data_bits_wstrb(accel_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(accel_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(accel_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(accel_io_memStreams_stores_0_wresp_bits),
    .io_memStreams_gathers_0_cmd_ready(accel_io_memStreams_gathers_0_cmd_ready),
    .io_memStreams_gathers_0_cmd_valid(accel_io_memStreams_gathers_0_cmd_valid),
    .io_memStreams_gathers_0_cmd_bits_addr_0(accel_io_memStreams_gathers_0_cmd_bits_addr_0),
    .io_memStreams_gathers_0_cmd_bits_addr_1(accel_io_memStreams_gathers_0_cmd_bits_addr_1),
    .io_memStreams_gathers_0_cmd_bits_addr_2(accel_io_memStreams_gathers_0_cmd_bits_addr_2),
    .io_memStreams_gathers_0_cmd_bits_addr_3(accel_io_memStreams_gathers_0_cmd_bits_addr_3),
    .io_memStreams_gathers_0_cmd_bits_addr_4(accel_io_memStreams_gathers_0_cmd_bits_addr_4),
    .io_memStreams_gathers_0_cmd_bits_addr_5(accel_io_memStreams_gathers_0_cmd_bits_addr_5),
    .io_memStreams_gathers_0_cmd_bits_addr_6(accel_io_memStreams_gathers_0_cmd_bits_addr_6),
    .io_memStreams_gathers_0_cmd_bits_addr_7(accel_io_memStreams_gathers_0_cmd_bits_addr_7),
    .io_memStreams_gathers_0_cmd_bits_addr_8(accel_io_memStreams_gathers_0_cmd_bits_addr_8),
    .io_memStreams_gathers_0_cmd_bits_addr_9(accel_io_memStreams_gathers_0_cmd_bits_addr_9),
    .io_memStreams_gathers_0_cmd_bits_addr_10(accel_io_memStreams_gathers_0_cmd_bits_addr_10),
    .io_memStreams_gathers_0_cmd_bits_addr_11(accel_io_memStreams_gathers_0_cmd_bits_addr_11),
    .io_memStreams_gathers_0_cmd_bits_addr_12(accel_io_memStreams_gathers_0_cmd_bits_addr_12),
    .io_memStreams_gathers_0_cmd_bits_addr_13(accel_io_memStreams_gathers_0_cmd_bits_addr_13),
    .io_memStreams_gathers_0_cmd_bits_addr_14(accel_io_memStreams_gathers_0_cmd_bits_addr_14),
    .io_memStreams_gathers_0_cmd_bits_addr_15(accel_io_memStreams_gathers_0_cmd_bits_addr_15),
    .io_memStreams_gathers_0_data_ready(accel_io_memStreams_gathers_0_data_ready),
    .io_memStreams_gathers_0_data_valid(accel_io_memStreams_gathers_0_data_valid),
    .io_memStreams_gathers_0_data_bits_0(accel_io_memStreams_gathers_0_data_bits_0),
    .io_memStreams_gathers_0_data_bits_1(accel_io_memStreams_gathers_0_data_bits_1),
    .io_memStreams_gathers_0_data_bits_2(accel_io_memStreams_gathers_0_data_bits_2),
    .io_memStreams_gathers_0_data_bits_3(accel_io_memStreams_gathers_0_data_bits_3),
    .io_memStreams_gathers_0_data_bits_4(accel_io_memStreams_gathers_0_data_bits_4),
    .io_memStreams_gathers_0_data_bits_5(accel_io_memStreams_gathers_0_data_bits_5),
    .io_memStreams_gathers_0_data_bits_6(accel_io_memStreams_gathers_0_data_bits_6),
    .io_memStreams_gathers_0_data_bits_7(accel_io_memStreams_gathers_0_data_bits_7),
    .io_memStreams_gathers_0_data_bits_8(accel_io_memStreams_gathers_0_data_bits_8),
    .io_memStreams_gathers_0_data_bits_9(accel_io_memStreams_gathers_0_data_bits_9),
    .io_memStreams_gathers_0_data_bits_10(accel_io_memStreams_gathers_0_data_bits_10),
    .io_memStreams_gathers_0_data_bits_11(accel_io_memStreams_gathers_0_data_bits_11),
    .io_memStreams_gathers_0_data_bits_12(accel_io_memStreams_gathers_0_data_bits_12),
    .io_memStreams_gathers_0_data_bits_13(accel_io_memStreams_gathers_0_data_bits_13),
    .io_memStreams_gathers_0_data_bits_14(accel_io_memStreams_gathers_0_data_bits_14),
    .io_memStreams_gathers_0_data_bits_15(accel_io_memStreams_gathers_0_data_bits_15),
    .io_memStreams_scatters_0_cmd_ready(accel_io_memStreams_scatters_0_cmd_ready),
    .io_memStreams_scatters_0_cmd_valid(accel_io_memStreams_scatters_0_cmd_valid),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_0(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_1(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_2(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_3(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_4(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_5(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_6(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_7(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_8(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_9(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_10(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_11(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_12(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_13(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_14(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_15(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15),
    .io_memStreams_scatters_0_cmd_bits_wdata_0(accel_io_memStreams_scatters_0_cmd_bits_wdata_0),
    .io_memStreams_scatters_0_cmd_bits_wdata_1(accel_io_memStreams_scatters_0_cmd_bits_wdata_1),
    .io_memStreams_scatters_0_cmd_bits_wdata_2(accel_io_memStreams_scatters_0_cmd_bits_wdata_2),
    .io_memStreams_scatters_0_cmd_bits_wdata_3(accel_io_memStreams_scatters_0_cmd_bits_wdata_3),
    .io_memStreams_scatters_0_cmd_bits_wdata_4(accel_io_memStreams_scatters_0_cmd_bits_wdata_4),
    .io_memStreams_scatters_0_cmd_bits_wdata_5(accel_io_memStreams_scatters_0_cmd_bits_wdata_5),
    .io_memStreams_scatters_0_cmd_bits_wdata_6(accel_io_memStreams_scatters_0_cmd_bits_wdata_6),
    .io_memStreams_scatters_0_cmd_bits_wdata_7(accel_io_memStreams_scatters_0_cmd_bits_wdata_7),
    .io_memStreams_scatters_0_cmd_bits_wdata_8(accel_io_memStreams_scatters_0_cmd_bits_wdata_8),
    .io_memStreams_scatters_0_cmd_bits_wdata_9(accel_io_memStreams_scatters_0_cmd_bits_wdata_9),
    .io_memStreams_scatters_0_cmd_bits_wdata_10(accel_io_memStreams_scatters_0_cmd_bits_wdata_10),
    .io_memStreams_scatters_0_cmd_bits_wdata_11(accel_io_memStreams_scatters_0_cmd_bits_wdata_11),
    .io_memStreams_scatters_0_cmd_bits_wdata_12(accel_io_memStreams_scatters_0_cmd_bits_wdata_12),
    .io_memStreams_scatters_0_cmd_bits_wdata_13(accel_io_memStreams_scatters_0_cmd_bits_wdata_13),
    .io_memStreams_scatters_0_cmd_bits_wdata_14(accel_io_memStreams_scatters_0_cmd_bits_wdata_14),
    .io_memStreams_scatters_0_cmd_bits_wdata_15(accel_io_memStreams_scatters_0_cmd_bits_wdata_15),
    .io_memStreams_scatters_0_wresp_ready(accel_io_memStreams_scatters_0_wresp_ready),
    .io_memStreams_scatters_0_wresp_valid(accel_io_memStreams_scatters_0_wresp_valid),
    .io_memStreams_scatters_0_wresp_bits(accel_io_memStreams_scatters_0_wresp_bits),
    .io_axiStreamsIn_0_TVALID(accel_io_axiStreamsIn_0_TVALID),
    .io_axiStreamsIn_0_TREADY(accel_io_axiStreamsIn_0_TREADY),
    .io_axiStreamsIn_0_TDATA(accel_io_axiStreamsIn_0_TDATA),
    .io_axiStreamsIn_0_TSTRB(accel_io_axiStreamsIn_0_TSTRB),
    .io_axiStreamsIn_0_TKEEP(accel_io_axiStreamsIn_0_TKEEP),
    .io_axiStreamsIn_0_TLAST(accel_io_axiStreamsIn_0_TLAST),
    .io_axiStreamsIn_0_TID(accel_io_axiStreamsIn_0_TID),
    .io_axiStreamsIn_0_TDEST(accel_io_axiStreamsIn_0_TDEST),
    .io_axiStreamsIn_0_TUSER(accel_io_axiStreamsIn_0_TUSER),
    .io_axiStreamsOut_0_TVALID(accel_io_axiStreamsOut_0_TVALID),
    .io_axiStreamsOut_0_TREADY(accel_io_axiStreamsOut_0_TREADY),
    .io_axiStreamsOut_0_TDATA(accel_io_axiStreamsOut_0_TDATA),
    .io_axiStreamsOut_0_TSTRB(accel_io_axiStreamsOut_0_TSTRB),
    .io_axiStreamsOut_0_TKEEP(accel_io_axiStreamsOut_0_TKEEP),
    .io_axiStreamsOut_0_TLAST(accel_io_axiStreamsOut_0_TLAST),
    .io_axiStreamsOut_0_TID(accel_io_axiStreamsOut_0_TID),
    .io_axiStreamsOut_0_TDEST(accel_io_axiStreamsOut_0_TDEST),
    .io_axiStreamsOut_0_TUSER(accel_io_axiStreamsOut_0_TUSER),
    .io_heap_0_req_valid(accel_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(accel_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(accel_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(accel_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(accel_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(accel_io_heap_0_resp_bits_sizeAddr),
    .io_argIns_0(accel_io_argIns_0),
    .io_argOuts_0_port_ready(accel_io_argOuts_0_port_ready),
    .io_argOuts_0_port_valid(accel_io_argOuts_0_port_valid),
    .io_argOuts_0_port_bits(accel_io_argOuts_0_port_bits),
    .io_argOuts_0_echo(accel_io_argOuts_0_echo),
    .io_argOuts_1_port_ready(accel_io_argOuts_1_port_ready),
    .io_argOuts_1_port_valid(accel_io_argOuts_1_port_valid),
    .io_argOuts_1_port_bits(accel_io_argOuts_1_port_bits),
    .io_argOuts_1_echo(accel_io_argOuts_1_echo),
    .io_argOuts_2_port_ready(accel_io_argOuts_2_port_ready),
    .io_argOuts_2_port_valid(accel_io_argOuts_2_port_valid),
    .io_argOuts_2_port_bits(accel_io_argOuts_2_port_bits),
    .io_argOuts_2_echo(accel_io_argOuts_2_echo),
    .io_argOuts_3_port_ready(accel_io_argOuts_3_port_ready),
    .io_argOuts_3_port_valid(accel_io_argOuts_3_port_valid),
    .io_argOuts_3_port_bits(accel_io_argOuts_3_port_bits),
    .io_argOuts_3_echo(accel_io_argOuts_3_echo),
    .io_argOuts_4_port_ready(accel_io_argOuts_4_port_ready),
    .io_argOuts_4_port_valid(accel_io_argOuts_4_port_valid),
    .io_argOuts_4_port_bits(accel_io_argOuts_4_port_bits),
    .io_argOuts_4_echo(accel_io_argOuts_4_echo),
    .io_argOuts_5_port_ready(accel_io_argOuts_5_port_ready),
    .io_argOuts_5_port_valid(accel_io_argOuts_5_port_valid),
    .io_argOuts_5_port_bits(accel_io_argOuts_5_port_bits),
    .io_argOuts_5_echo(accel_io_argOuts_5_echo),
    .io_argOuts_6_port_ready(accel_io_argOuts_6_port_ready),
    .io_argOuts_6_port_valid(accel_io_argOuts_6_port_valid),
    .io_argOuts_6_port_bits(accel_io_argOuts_6_port_bits),
    .io_argOuts_6_echo(accel_io_argOuts_6_echo),
    .io_argOuts_7_port_ready(accel_io_argOuts_7_port_ready),
    .io_argOuts_7_port_valid(accel_io_argOuts_7_port_valid),
    .io_argOuts_7_port_bits(accel_io_argOuts_7_port_bits),
    .io_argOuts_7_echo(accel_io_argOuts_7_echo),
    .io_argOuts_8_port_ready(accel_io_argOuts_8_port_ready),
    .io_argOuts_8_port_valid(accel_io_argOuts_8_port_valid),
    .io_argOuts_8_port_bits(accel_io_argOuts_8_port_bits),
    .io_argOuts_8_echo(accel_io_argOuts_8_echo),
    .io_argOuts_9_port_ready(accel_io_argOuts_9_port_ready),
    .io_argOuts_9_port_valid(accel_io_argOuts_9_port_valid),
    .io_argOuts_9_port_bits(accel_io_argOuts_9_port_bits),
    .io_argOuts_9_echo(accel_io_argOuts_9_echo)
  );
  FringeZynq FringeZynq ( // @[KCU1500.scala 21:24:@52482.4]
    .clock(FringeZynq_clock),
    .reset(FringeZynq_reset),
    .io_S_AXI_AWADDR(FringeZynq_io_S_AXI_AWADDR),
    .io_S_AXI_AWPROT(FringeZynq_io_S_AXI_AWPROT),
    .io_S_AXI_AWVALID(FringeZynq_io_S_AXI_AWVALID),
    .io_S_AXI_AWREADY(FringeZynq_io_S_AXI_AWREADY),
    .io_S_AXI_ARADDR(FringeZynq_io_S_AXI_ARADDR),
    .io_S_AXI_ARPROT(FringeZynq_io_S_AXI_ARPROT),
    .io_S_AXI_ARVALID(FringeZynq_io_S_AXI_ARVALID),
    .io_S_AXI_ARREADY(FringeZynq_io_S_AXI_ARREADY),
    .io_S_AXI_WDATA(FringeZynq_io_S_AXI_WDATA),
    .io_S_AXI_WSTRB(FringeZynq_io_S_AXI_WSTRB),
    .io_S_AXI_WVALID(FringeZynq_io_S_AXI_WVALID),
    .io_S_AXI_WREADY(FringeZynq_io_S_AXI_WREADY),
    .io_S_AXI_RDATA(FringeZynq_io_S_AXI_RDATA),
    .io_S_AXI_RRESP(FringeZynq_io_S_AXI_RRESP),
    .io_S_AXI_RVALID(FringeZynq_io_S_AXI_RVALID),
    .io_S_AXI_RREADY(FringeZynq_io_S_AXI_RREADY),
    .io_S_AXI_BRESP(FringeZynq_io_S_AXI_BRESP),
    .io_S_AXI_BVALID(FringeZynq_io_S_AXI_BVALID),
    .io_S_AXI_BREADY(FringeZynq_io_S_AXI_BREADY),
    .io_M_AXI_0_AWLEN(FringeZynq_io_M_AXI_0_AWLEN),
    .io_M_AXI_0_ARLEN(FringeZynq_io_M_AXI_0_ARLEN),
    .io_enable(FringeZynq_io_enable),
    .io_done(FringeZynq_io_done),
    .io_reset(FringeZynq_io_reset),
    .io_argIns_0(FringeZynq_io_argIns_0),
    .io_argOuts_0_valid(FringeZynq_io_argOuts_0_valid),
    .io_argOuts_0_bits(FringeZynq_io_argOuts_0_bits),
    .io_argOuts_1_valid(FringeZynq_io_argOuts_1_valid),
    .io_argOuts_1_bits(FringeZynq_io_argOuts_1_bits),
    .io_argOuts_2_valid(FringeZynq_io_argOuts_2_valid),
    .io_argOuts_2_bits(FringeZynq_io_argOuts_2_bits),
    .io_argOuts_3_valid(FringeZynq_io_argOuts_3_valid),
    .io_argOuts_3_bits(FringeZynq_io_argOuts_3_bits),
    .io_argOuts_4_valid(FringeZynq_io_argOuts_4_valid),
    .io_argOuts_4_bits(FringeZynq_io_argOuts_4_bits),
    .io_argOuts_5_valid(FringeZynq_io_argOuts_5_valid),
    .io_argOuts_5_bits(FringeZynq_io_argOuts_5_bits),
    .io_argOuts_6_valid(FringeZynq_io_argOuts_6_valid),
    .io_argOuts_6_bits(FringeZynq_io_argOuts_6_bits),
    .io_argOuts_7_valid(FringeZynq_io_argOuts_7_valid),
    .io_argOuts_7_bits(FringeZynq_io_argOuts_7_bits),
    .io_argOuts_8_valid(FringeZynq_io_argOuts_8_valid),
    .io_argOuts_8_bits(FringeZynq_io_argOuts_8_bits),
    .io_argOuts_9_valid(FringeZynq_io_argOuts_9_valid),
    .io_argOuts_9_bits(FringeZynq_io_argOuts_9_bits),
    .io_heap_0_req_valid(FringeZynq_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(FringeZynq_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(FringeZynq_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(FringeZynq_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(FringeZynq_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(FringeZynq_io_heap_0_resp_bits_sizeAddr)
  );
  assign io_rdata = 1'h0;
  assign io_S_AXI_AWREADY = FringeZynq_io_S_AXI_AWREADY; // @[KCU1500.scala 24:21:@52500.4]
  assign io_S_AXI_ARREADY = FringeZynq_io_S_AXI_ARREADY; // @[KCU1500.scala 24:21:@52496.4]
  assign io_S_AXI_WREADY = FringeZynq_io_S_AXI_WREADY; // @[KCU1500.scala 24:21:@52492.4]
  assign io_S_AXI_RDATA = FringeZynq_io_S_AXI_RDATA; // @[KCU1500.scala 24:21:@52491.4]
  assign io_S_AXI_RRESP = FringeZynq_io_S_AXI_RRESP; // @[KCU1500.scala 24:21:@52490.4]
  assign io_S_AXI_RVALID = FringeZynq_io_S_AXI_RVALID; // @[KCU1500.scala 24:21:@52489.4]
  assign io_S_AXI_BRESP = FringeZynq_io_S_AXI_BRESP; // @[KCU1500.scala 24:21:@52487.4]
  assign io_S_AXI_BVALID = FringeZynq_io_S_AXI_BVALID; // @[KCU1500.scala 24:21:@52486.4]
  assign io_M_AXI_0_AWID = 4'h0; // @[KCU1500.scala 31:14:@52562.4]
  assign io_M_AXI_0_AWUSER = 4'h0; // @[KCU1500.scala 31:14:@52561.4]
  assign io_M_AXI_0_AWADDR = 32'h0; // @[KCU1500.scala 31:14:@52560.4]
  assign io_M_AXI_0_AWLEN = FringeZynq_io_M_AXI_0_AWLEN; // @[KCU1500.scala 31:14:@52559.4]
  assign io_M_AXI_0_AWSIZE = 3'h6; // @[KCU1500.scala 31:14:@52558.4]
  assign io_M_AXI_0_AWBURST = 2'h1; // @[KCU1500.scala 31:14:@52557.4]
  assign io_M_AXI_0_AWLOCK = 1'h0; // @[KCU1500.scala 31:14:@52556.4]
  assign io_M_AXI_0_AWCACHE = 4'h3; // @[KCU1500.scala 31:14:@52555.4]
  assign io_M_AXI_0_AWPROT = 3'h0; // @[KCU1500.scala 31:14:@52554.4]
  assign io_M_AXI_0_AWQOS = 4'h0; // @[KCU1500.scala 31:14:@52553.4]
  assign io_M_AXI_0_AWVALID = 1'h0; // @[KCU1500.scala 31:14:@52552.4]
  assign io_M_AXI_0_ARID = 4'h0; // @[KCU1500.scala 31:14:@52550.4]
  assign io_M_AXI_0_ARUSER = 4'h0; // @[KCU1500.scala 31:14:@52549.4]
  assign io_M_AXI_0_ARADDR = 32'h0; // @[KCU1500.scala 31:14:@52548.4]
  assign io_M_AXI_0_ARLEN = FringeZynq_io_M_AXI_0_ARLEN; // @[KCU1500.scala 31:14:@52547.4]
  assign io_M_AXI_0_ARSIZE = 3'h6; // @[KCU1500.scala 31:14:@52546.4]
  assign io_M_AXI_0_ARBURST = 2'h1; // @[KCU1500.scala 31:14:@52545.4]
  assign io_M_AXI_0_ARLOCK = 1'h0; // @[KCU1500.scala 31:14:@52544.4]
  assign io_M_AXI_0_ARCACHE = 4'h3; // @[KCU1500.scala 31:14:@52543.4]
  assign io_M_AXI_0_ARPROT = 3'h0; // @[KCU1500.scala 31:14:@52542.4]
  assign io_M_AXI_0_ARQOS = 4'h0; // @[KCU1500.scala 31:14:@52541.4]
  assign io_M_AXI_0_ARVALID = 1'h0; // @[KCU1500.scala 31:14:@52540.4]
  assign io_M_AXI_0_WDATA = 512'h0; // @[KCU1500.scala 31:14:@52538.4]
  assign io_M_AXI_0_WSTRB = 64'h0; // @[KCU1500.scala 31:14:@52537.4]
  assign io_M_AXI_0_WLAST = 1'h0; // @[KCU1500.scala 31:14:@52536.4]
  assign io_M_AXI_0_WVALID = 1'h0; // @[KCU1500.scala 31:14:@52535.4]
  assign io_M_AXI_0_RREADY = 1'h0; // @[KCU1500.scala 31:14:@52527.4]
  assign io_M_AXI_0_BREADY = 1'h0; // @[KCU1500.scala 31:14:@52522.4]
  assign io_AXIS_IN_TREADY = accel_io_axiStreamsIn_0_TREADY; // @[KCU1500.scala 27:16:@52511.4]
  assign io_AXIS_OUT_TVALID = accel_io_axiStreamsOut_0_TVALID; // @[KCU1500.scala 28:17:@52521.4]
  assign io_AXIS_OUT_TDATA = accel_io_axiStreamsOut_0_TDATA; // @[KCU1500.scala 28:17:@52519.4]
  assign io_AXIS_OUT_TSTRB = accel_io_axiStreamsOut_0_TSTRB; // @[KCU1500.scala 28:17:@52518.4]
  assign io_AXIS_OUT_TKEEP = accel_io_axiStreamsOut_0_TKEEP; // @[KCU1500.scala 28:17:@52517.4]
  assign io_AXIS_OUT_TLAST = accel_io_axiStreamsOut_0_TLAST; // @[KCU1500.scala 28:17:@52516.4]
  assign io_AXIS_OUT_TID = accel_io_axiStreamsOut_0_TID; // @[KCU1500.scala 28:17:@52515.4]
  assign io_AXIS_OUT_TDEST = accel_io_axiStreamsOut_0_TDEST; // @[KCU1500.scala 28:17:@52514.4]
  assign io_AXIS_OUT_TUSER = {{480'd0}, accel_io_axiStreamsOut_0_TUSER}; // @[KCU1500.scala 28:17:@52513.4]
  assign accel_clock = clock; // @[:@52291.4]
  assign accel_reset = FringeZynq_io_reset; // @[:@52292.4 KCU1500.scala 61:17:@52891.4]
  assign accel_io_enable = FringeZynq_io_enable; // @[KCU1500.scala 58:21:@52887.4]
  assign accel_io_reset = 1'h0;
  assign accel_io_memStreams_loads_0_cmd_ready = 1'h0; // @[KCU1500.scala 56:26:@52880.4]
  assign accel_io_memStreams_loads_0_data_valid = 1'h0; // @[KCU1500.scala 56:26:@52875.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_0 = 32'h0; // @[KCU1500.scala 56:26:@52859.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_1 = 32'h0; // @[KCU1500.scala 56:26:@52860.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_2 = 32'h0; // @[KCU1500.scala 56:26:@52861.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_3 = 32'h0; // @[KCU1500.scala 56:26:@52862.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_4 = 32'h0; // @[KCU1500.scala 56:26:@52863.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_5 = 32'h0; // @[KCU1500.scala 56:26:@52864.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_6 = 32'h0; // @[KCU1500.scala 56:26:@52865.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_7 = 32'h0; // @[KCU1500.scala 56:26:@52866.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_8 = 32'h0; // @[KCU1500.scala 56:26:@52867.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_9 = 32'h0; // @[KCU1500.scala 56:26:@52868.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_10 = 32'h0; // @[KCU1500.scala 56:26:@52869.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_11 = 32'h0; // @[KCU1500.scala 56:26:@52870.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_12 = 32'h0; // @[KCU1500.scala 56:26:@52871.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_13 = 32'h0; // @[KCU1500.scala 56:26:@52872.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_14 = 32'h0; // @[KCU1500.scala 56:26:@52873.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_15 = 32'h0; // @[KCU1500.scala 56:26:@52874.4]
  assign accel_io_memStreams_stores_0_cmd_ready = 1'h0; // @[KCU1500.scala 56:26:@52858.4]
  assign accel_io_memStreams_stores_0_data_ready = 1'h0; // @[KCU1500.scala 56:26:@52854.4]
  assign accel_io_memStreams_stores_0_wresp_valid = 1'h0; // @[KCU1500.scala 56:26:@52834.4]
  assign accel_io_memStreams_stores_0_wresp_bits = 1'h0; // @[KCU1500.scala 56:26:@52833.4]
  assign accel_io_memStreams_gathers_0_cmd_ready = 1'h0; // @[KCU1500.scala 56:26:@52832.4]
  assign accel_io_memStreams_gathers_0_data_valid = 1'h0; // @[KCU1500.scala 56:26:@52813.4]
  assign accel_io_memStreams_gathers_0_data_bits_0 = 32'h0; // @[KCU1500.scala 56:26:@52797.4]
  assign accel_io_memStreams_gathers_0_data_bits_1 = 32'h0; // @[KCU1500.scala 56:26:@52798.4]
  assign accel_io_memStreams_gathers_0_data_bits_2 = 32'h0; // @[KCU1500.scala 56:26:@52799.4]
  assign accel_io_memStreams_gathers_0_data_bits_3 = 32'h0; // @[KCU1500.scala 56:26:@52800.4]
  assign accel_io_memStreams_gathers_0_data_bits_4 = 32'h0; // @[KCU1500.scala 56:26:@52801.4]
  assign accel_io_memStreams_gathers_0_data_bits_5 = 32'h0; // @[KCU1500.scala 56:26:@52802.4]
  assign accel_io_memStreams_gathers_0_data_bits_6 = 32'h0; // @[KCU1500.scala 56:26:@52803.4]
  assign accel_io_memStreams_gathers_0_data_bits_7 = 32'h0; // @[KCU1500.scala 56:26:@52804.4]
  assign accel_io_memStreams_gathers_0_data_bits_8 = 32'h0; // @[KCU1500.scala 56:26:@52805.4]
  assign accel_io_memStreams_gathers_0_data_bits_9 = 32'h0; // @[KCU1500.scala 56:26:@52806.4]
  assign accel_io_memStreams_gathers_0_data_bits_10 = 32'h0; // @[KCU1500.scala 56:26:@52807.4]
  assign accel_io_memStreams_gathers_0_data_bits_11 = 32'h0; // @[KCU1500.scala 56:26:@52808.4]
  assign accel_io_memStreams_gathers_0_data_bits_12 = 32'h0; // @[KCU1500.scala 56:26:@52809.4]
  assign accel_io_memStreams_gathers_0_data_bits_13 = 32'h0; // @[KCU1500.scala 56:26:@52810.4]
  assign accel_io_memStreams_gathers_0_data_bits_14 = 32'h0; // @[KCU1500.scala 56:26:@52811.4]
  assign accel_io_memStreams_gathers_0_data_bits_15 = 32'h0; // @[KCU1500.scala 56:26:@52812.4]
  assign accel_io_memStreams_scatters_0_cmd_ready = 1'h0; // @[KCU1500.scala 56:26:@52796.4]
  assign accel_io_memStreams_scatters_0_wresp_valid = 1'h0; // @[KCU1500.scala 56:26:@52761.4]
  assign accel_io_memStreams_scatters_0_wresp_bits = 1'h0; // @[KCU1500.scala 56:26:@52760.4]
  assign accel_io_axiStreamsIn_0_TVALID = io_AXIS_IN_TVALID; // @[KCU1500.scala 27:16:@52512.4]
  assign accel_io_axiStreamsIn_0_TDATA = io_AXIS_IN_TDATA[255:0]; // @[KCU1500.scala 27:16:@52510.4]
  assign accel_io_axiStreamsIn_0_TSTRB = io_AXIS_IN_TSTRB[31:0]; // @[KCU1500.scala 27:16:@52509.4]
  assign accel_io_axiStreamsIn_0_TKEEP = io_AXIS_IN_TKEEP[31:0]; // @[KCU1500.scala 27:16:@52508.4]
  assign accel_io_axiStreamsIn_0_TLAST = io_AXIS_IN_TLAST; // @[KCU1500.scala 27:16:@52507.4]
  assign accel_io_axiStreamsIn_0_TID = io_AXIS_IN_TID; // @[KCU1500.scala 27:16:@52506.4]
  assign accel_io_axiStreamsIn_0_TDEST = io_AXIS_IN_TDEST; // @[KCU1500.scala 27:16:@52505.4]
  assign accel_io_axiStreamsIn_0_TUSER = io_AXIS_IN_TUSER[31:0]; // @[KCU1500.scala 27:16:@52504.4]
  assign accel_io_axiStreamsOut_0_TREADY = io_AXIS_OUT_TREADY; // @[KCU1500.scala 28:17:@52520.4]
  assign accel_io_heap_0_resp_valid = FringeZynq_io_heap_0_resp_valid; // @[KCU1500.scala 57:20:@52883.4]
  assign accel_io_heap_0_resp_bits_allocDealloc = FringeZynq_io_heap_0_resp_bits_allocDealloc; // @[KCU1500.scala 57:20:@52882.4]
  assign accel_io_heap_0_resp_bits_sizeAddr = FringeZynq_io_heap_0_resp_bits_sizeAddr; // @[KCU1500.scala 57:20:@52881.4]
  assign accel_io_argIns_0 = FringeZynq_io_argIns_0; // @[KCU1500.scala 41:21:@52728.4]
  assign accel_io_argOuts_0_port_ready = 1'h0;
  assign accel_io_argOuts_0_echo = 64'h0; // @[KCU1500.scala 47:24:@52749.4]
  assign accel_io_argOuts_1_port_ready = 1'h0;
  assign accel_io_argOuts_1_echo = 64'h0; // @[KCU1500.scala 47:24:@52750.4]
  assign accel_io_argOuts_2_port_ready = 1'h0;
  assign accel_io_argOuts_2_echo = 64'h0; // @[KCU1500.scala 47:24:@52751.4]
  assign accel_io_argOuts_3_port_ready = 1'h0;
  assign accel_io_argOuts_3_echo = 64'h0; // @[KCU1500.scala 47:24:@52752.4]
  assign accel_io_argOuts_4_port_ready = 1'h0;
  assign accel_io_argOuts_4_echo = 64'h0; // @[KCU1500.scala 47:24:@52753.4]
  assign accel_io_argOuts_5_port_ready = 1'h0;
  assign accel_io_argOuts_5_echo = 64'h0; // @[KCU1500.scala 47:24:@52754.4]
  assign accel_io_argOuts_6_port_ready = 1'h0;
  assign accel_io_argOuts_6_echo = 64'h0; // @[KCU1500.scala 47:24:@52755.4]
  assign accel_io_argOuts_7_port_ready = 1'h0;
  assign accel_io_argOuts_7_echo = 64'h0; // @[KCU1500.scala 47:24:@52756.4]
  assign accel_io_argOuts_8_port_ready = 1'h0;
  assign accel_io_argOuts_8_echo = 64'h0; // @[KCU1500.scala 47:24:@52757.4]
  assign accel_io_argOuts_9_port_ready = 1'h0;
  assign accel_io_argOuts_9_echo = 64'h0; // @[KCU1500.scala 47:24:@52758.4]
  assign FringeZynq_clock = clock; // @[:@52483.4]
  assign FringeZynq_reset = reset; // @[:@52484.4 KCU1500.scala 60:18:@52890.4]
  assign FringeZynq_io_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[KCU1500.scala 24:21:@52503.4]
  assign FringeZynq_io_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[KCU1500.scala 24:21:@52502.4]
  assign FringeZynq_io_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[KCU1500.scala 24:21:@52501.4]
  assign FringeZynq_io_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[KCU1500.scala 24:21:@52499.4]
  assign FringeZynq_io_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[KCU1500.scala 24:21:@52498.4]
  assign FringeZynq_io_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[KCU1500.scala 24:21:@52497.4]
  assign FringeZynq_io_S_AXI_WDATA = io_S_AXI_WDATA; // @[KCU1500.scala 24:21:@52495.4]
  assign FringeZynq_io_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[KCU1500.scala 24:21:@52494.4]
  assign FringeZynq_io_S_AXI_WVALID = io_S_AXI_WVALID; // @[KCU1500.scala 24:21:@52493.4]
  assign FringeZynq_io_S_AXI_RREADY = io_S_AXI_RREADY; // @[KCU1500.scala 24:21:@52488.4]
  assign FringeZynq_io_S_AXI_BREADY = io_S_AXI_BREADY; // @[KCU1500.scala 24:21:@52485.4]
  assign FringeZynq_io_done = accel_io_done; // @[KCU1500.scala 59:20:@52888.4]
  assign FringeZynq_io_argOuts_0_valid = accel_io_argOuts_0_port_valid; // @[KCU1500.scala 44:26:@52730.4]
  assign FringeZynq_io_argOuts_0_bits = accel_io_argOuts_0_port_bits; // @[KCU1500.scala 43:25:@52729.4]
  assign FringeZynq_io_argOuts_1_valid = accel_io_argOuts_1_port_valid; // @[KCU1500.scala 44:26:@52732.4]
  assign FringeZynq_io_argOuts_1_bits = accel_io_argOuts_1_port_bits; // @[KCU1500.scala 43:25:@52731.4]
  assign FringeZynq_io_argOuts_2_valid = accel_io_argOuts_2_port_valid; // @[KCU1500.scala 44:26:@52734.4]
  assign FringeZynq_io_argOuts_2_bits = accel_io_argOuts_2_port_bits; // @[KCU1500.scala 43:25:@52733.4]
  assign FringeZynq_io_argOuts_3_valid = accel_io_argOuts_3_port_valid; // @[KCU1500.scala 44:26:@52736.4]
  assign FringeZynq_io_argOuts_3_bits = accel_io_argOuts_3_port_bits; // @[KCU1500.scala 43:25:@52735.4]
  assign FringeZynq_io_argOuts_4_valid = accel_io_argOuts_4_port_valid; // @[KCU1500.scala 44:26:@52738.4]
  assign FringeZynq_io_argOuts_4_bits = accel_io_argOuts_4_port_bits; // @[KCU1500.scala 43:25:@52737.4]
  assign FringeZynq_io_argOuts_5_valid = accel_io_argOuts_5_port_valid; // @[KCU1500.scala 44:26:@52740.4]
  assign FringeZynq_io_argOuts_5_bits = accel_io_argOuts_5_port_bits; // @[KCU1500.scala 43:25:@52739.4]
  assign FringeZynq_io_argOuts_6_valid = accel_io_argOuts_6_port_valid; // @[KCU1500.scala 44:26:@52742.4]
  assign FringeZynq_io_argOuts_6_bits = accel_io_argOuts_6_port_bits; // @[KCU1500.scala 43:25:@52741.4]
  assign FringeZynq_io_argOuts_7_valid = accel_io_argOuts_7_port_valid; // @[KCU1500.scala 44:26:@52744.4]
  assign FringeZynq_io_argOuts_7_bits = accel_io_argOuts_7_port_bits; // @[KCU1500.scala 43:25:@52743.4]
  assign FringeZynq_io_argOuts_8_valid = accel_io_argOuts_8_port_valid; // @[KCU1500.scala 44:26:@52746.4]
  assign FringeZynq_io_argOuts_8_bits = accel_io_argOuts_8_port_bits; // @[KCU1500.scala 43:25:@52745.4]
  assign FringeZynq_io_argOuts_9_valid = accel_io_argOuts_9_port_valid; // @[KCU1500.scala 44:26:@52748.4]
  assign FringeZynq_io_argOuts_9_bits = accel_io_argOuts_9_port_bits; // @[KCU1500.scala 43:25:@52747.4]
  assign FringeZynq_io_heap_0_req_valid = accel_io_heap_0_req_valid; // @[KCU1500.scala 57:20:@52886.4]
  assign FringeZynq_io_heap_0_req_bits_allocDealloc = accel_io_heap_0_req_bits_allocDealloc; // @[KCU1500.scala 57:20:@52885.4]
  assign FringeZynq_io_heap_0_req_bits_sizeAddr = accel_io_heap_0_req_bits_sizeAddr; // @[KCU1500.scala 57:20:@52884.4]
endmodule
module SRAMVerilogAWS
#(
    parameter WORDS = 1024,
    parameter AWIDTH = 10,
    parameter DWIDTH = 32)
(
    input clk,
    input [AWIDTH-1:0] raddr,
    input [AWIDTH-1:0] waddr,
    input raddrEn,
    input waddrEn,
    input wen,
    input [DWIDTH-1:0] wdata,
    input backpressure,
    output reg [DWIDTH-1:0] rdata
);

    reg [DWIDTH-1:0] mem [0:WORDS-1];

    always @(posedge clk) begin
      if (wen) mem[waddr] <= wdata;
      if (backpressure) rdata <= mem[raddr];
    end

endmodule
